PK   W�X�Ή�0  Jt    cirkitFile.json�}K�$7��_Y���	���:f}�=�=H��?[�[]Y�J��W�_�gd)�a�atm���A���F{�����K����c���?��������0�w?�/�/��_���/O�_���R���ï��������_�<�?�>j��Jk[�U���_u���7�i�۶k�����ﯞ.����UטN��(�
]ʾh�4E��֭��<�;f��l8���V�4�wE�;_辩����B�ږNԃiţd}�f�VԆd����襁t9NW�h��Ei���Z�A6�]O�#(�PS<���8�)&�P{j�����ǥ����!� ̖�ނ���CB�O(x�tA+/l�`Η���9_3�3e����s>����$��$��$��$s�$s�$��`��ڮ0Z���R�4R��JuVhc"�+4�^}h:���t��C��M�O>4�fh:�7�����N�;f����M���N�;4��wh:s��v���aVb�J9N��U5Ⱥ��U�N[u�:�׹:�*5�8A�)gCM9NjނS����e�r� Ԕ߄��'5�#c�)�I��������U;um��mݘ��Ck��ܔ���}7m�`�i��cL5�^��LE*��
F�8���
�9��\R���pPS���qPS��䠦l0��15)� rPS�K����1�H��n��M_��A�x]8[��M�e���~C�#-2=��"ә��
�;NȘs��9���k�a(��eT�^m������Z:7X��4�u�*��Van �p���r��2�j�^�������T1vInυL[���0���Sf)$�h��N� P�1mJOC�n�Ov�M�>>�H
֚��eс>>5�fA���2�@�����A����pH��Gs�y�i��N�E�t:�M��Eh:��^P�d�&b;�.�5�y���]��hk��A7�Q-�k�v��b��)��hJ&b�)���d"��R�jނS
B͒�d�BM� jJB�)���r��y���t��OǊ1�T��X16���#�b��bɈH�@��D�X16���A<Xު�3jުQf���0Ԕ� �f)p2V�f)p2V�f��H��O[��2��*h�2n/��j�X�ܛR�49�)� �����Ej�|��"5�@c���4�1A�@M,�ꋃ�441�AM,�:���,X M�W����#Z�)N�z�&v��C����7
:�7
�q���s�	fB�#�Lh~ġ��G���H@��d��Iw&���xh>��"�|��E
 o>Vl8j�.<P�M����|8]�
��%�l�K}4��ӱ�M�����������r���k��#ʃ"�Т�h��&�C�j��zg��g@1�/B��/�MIdˠ��#-fP����=�upP�=�}Y:bu�Z� Ŕ��Y9f	�EK�ú���DvZ-��_\(>�0p9p0I� ���#e��&�<L,�p����2�<\,�l�̳�2��h�q(�}B��3@I��&9���A+�3@I�Z��J�_���P����2g�����9�<���Rh�r���G0^U����$��0�zѕm�s���怙��Nږ���u�[b��S�X`&�*���&�m+��5�L28��*?��Y���05�Gٔ�ך�#p�h<,׀�#p=g<��f��p�eS"m{�U���mr��2�<�SV Z��--� %�Gh�Y
X4�J���:�����t��4�:+n���Vq+���ih�S�FC+��;�4e��<hyS(IO-v� %�	��O�$�h�")��ꢻ���T��d}��U?�z�y5�oӵv8`&���8�
���ԝ�=A��%�	µ+9�^��+Yr��$��ay��n����KU�k�k=�0�=A��$�5��W�0��=Տ�
�T�k�3q�u�� ,#�Zc��w0�`�h��H{�p1EZS�J�|�eq��V<�5&Z�W�hB\_�%qu�V$�%��8�`�~Bʀ��	� f�'����`~{��s�r
L;O�)0�<��5�&�� ��f���`�>%�l�LښAS�s���ÀM��g ��hvz0y�8����� ��p4�=�r3Д��$e�����\��ؔ�E�ǿ��{*�����禂�~}�?Qā��|(2���Ť����|(�=�S��P�{�����#�J������L̛�{E�y�W�a`���EyxX�ab���e.��dp.�y6\��p��p8�%�Op*8JR����|(II���$�N�CI��
·��8�%�/p*8J~IJ)8<�eb�<ܛ���T�`�0pڶ�S�3����i�
O� ��pqڶ�S�3����2�<\�6�T�`�p����*�<\�2�i�M�CI��h*8J�uI��h*x
�
·��#8<M�CI�
·��:8�%�uh*8JR����|(I~�S��P�����$�N�C��/I�N��u��7��=A<<�<���T�`��p��S�3H�<\���T�`�pq��S�3����iOO� &�=A<<�L�D���Tp>������|(y�%y��Tp>��цS��l����O�
·��h*8JZ���|(y�%��T�\��y�p/`�é���a`�&�S�3���ÀM��g�zy����T�`�l8`�©�Q0p*8
����� ��`*8JR����|(�l��}�Ͽ���|��~�A���_�^���_>�m�=>}~|~����?lwm���TE���Т��(��ʲur(��zw]�^�Bv�*t�tQ��/�ol٨F�J��������ui�v���G_��֕,��4�w�З�#�6����k����B�R�.�КJ7u/]3=����M "Fb�,����j
����vE���/�F۲U6���G}f� �T����U��hM!î� �jы�-���fob.��z3被��pTN՚��j��y?Tӳsٿ� ̜o����3�q�kk���a�{z胶l|UT�J�\]
���&����E�.������ F��
��6��{���D	D5�af�j���L��D0Kf��Ln3���,X��:w���6GO�>�h&�6B�u>��U��J^�_m/ʶ����L̂0K ��z��`{�1.�`�6;�T�Lp0Se���`��h`R��������6�N�.����mP\�ڞ���a��[V
�
3�38,��f�����,����0b��o&�'5X�s���f�z�,'��*��w�J�� ;X%`#������v�9�ٚ!V�"xQ�j!l��M[X%E[J]�c�O�ߴo�n�E5Fuӹ`?�����J���N��*hךb�}�k[�ި���Y�}'���+����У��%����z�x��}��(��y��>��gf؀�@��	"X�4���%�V3Q�
�k���U�+�	jt�+WԲ�S�f��`ii�f�u$�7��V�F���2�G�!��-۶��2L��B-HGzԤ=�?jҫ����[2m~B�k��R�E���`��ht�e[��.��M+�~(u�᫛Vښ�������]]��2S%�&fh�xG�(�s]?Rm�@��UP�U�5�n\��ZHZ��0�f����l��^R^�M!|]��Vu�w�,_4&Lk�0CQ�}�U���U��%3�a$f�n�ߤ�3�� e�湴��/����Nٲ�|W�)���ҫ.XY����*��j�Cd���`f�.|���h��iҖ��ں��q�4!�!̴����i����l�)�7M'zz�AeG��m崯mѶU3f~[2X�R��4�y�e�V]S�e��]D�Y8SWEk+�Mi۾��H2Tm�il�X��@�h]_˰;m����	S��nuo�33�Q�l�z����N뀺iDQ��g
���egˈ7�J�mM]
;�>��*h���e�~]����Rw���N&�P�p()O �D�:�$f#E�j�)G�S���eg;�e?��%�HW¼��bj��=؛'O�ٜ��s�a��LFm Y��L��a���b�����ˏ?�D�A�f1Zs�2Ci/�l���"B���"��!݉֫�H�L��;���ʶ�}عH�����|��S��F�M��骐�sd[v���KKd6�
��f3���38�yr�L�9<1a&��M%ذ|;�.�'^�3�8�y&+F�2�8�AWa̠��f�U��y���b�A��W�ו�5�������Ҩ��j��BM����yY�T�3��G:}�$t�Y��=� n���I�Ēqw��P�
K��)[g�PS��٭*f8��������/X�u*�%��������L�c����ͼ}�|3�Xq0�D	g�y�}K�zԤ-�)�C_١(}�b��,�9�ʲ�Av��B�4١0}�e��(�Y�$
�����W��h��D����I����u=j�+�6����V�{bף��O�o�]��g�P��>�
���ߌu��㛱^��؃PO�]�A�"�Z���G񧡖��37m�ݚ�GMۃ`�kj:v���f,8)N����������>\X�rj���;������TG0�9jb��7X���>|�BM��j�/��5�* {�a��X�-='�����!��g��g��J�f}3��8����kd�S�Q�R���?~|os�����o}�X�Z����&��G�G�?�pD�n���%8�;�]��lx@sv�@��O0�M��0{��F �2~I��d�B�{2��_%�1�&�˂;
���(G<cׇ�f�'���� ��|�O�	`�t�'���A�S�|��O��>�W"&�,SG�6\9�&�+��pU� �2L�$G<	�'�ك�O �7� fGn>���|�]�w3���Cvs��7D�����٢�k�$D����	�>���9@������wt����$�E[@pċ/|�����/7��ong�M8�A߄���5H)�CB���x�6�
p�a��1��l7u���E	8�q(>{��G<�'`O�􈇣�d�O��	�$ґ+�] ��Z�F ���~�
��@ߺ�M+�O^�F ���~�"���@���p�|+�W��p��@��}*+�>�Ŭ(�tԹ-":=��S�
��֍1���|b+J�/m�7����~��n�F ���n��pE	8�1�x��or�)8�i�Q�]q
�x�k�����EL@<Y���1
@y��"�b�*e�8FF)����Kp�0�Q�D�I��h��e���5C�ɂT ���ws��g� !\��l+�W���%�'���9Rkp�;�� ��]f����^f�����~��PJ��	�)��Q8�EL>̇1#�2��y|j	�x��O@�����v"W���Y��8ʢ�x�4~�v�C�Q�xϔy��(���鮃鲴yx�îL'��s� �Y>�wfwrR��
��`w��_��Ј�7�0����(�Y����K���I�]\v��I�<�̷��˰�yz��~�N�3�{�iͅ>�8� ���˂��x�]rS�8U����P�Z'��HB~��s�H������0�9Z�ѝh�*��	'��}�
�[+ۮ��+�YO�A��str2���ߑ��ⓥ!ꍡnD Q�uQ��v�S5��8��F��Oe@�fYb�T�l��L��=�39�N�  Kܒ��rI�r`i/�G'v# ���(���E[��*�x'��(ߎ��I��A*�hW9ڇ��I�lgWY$�/�Yn�Y$ow���r�!�j���i�k���7��k��=�V��p��� n���v���� n%���},�{��[�3��_P��c�r��SnB��-Xc��8��
�G��w����rXD�i��ډ<�<X옧��Lf���Ky:z����@���z�\h�	�^�	�^�	�^���^��^%V {t� ��p�|!��r�%��x.����]���&�7��?*{`��	 BW`/�p:B�m �m�� �k)Y���Zʞ����rv�������|�P;D��R<D�l����c���ae����g?��35�1�/P����}68���LN���������c��`q���g�>��i�����s����`����u�7}p�@D僻?p���8Q�=�UטN��(�
]ʾh�.���[9T��e1  Ե��q�+:���o�q�B�ږNԃiE��(B �B����CNa�[�
'�������<?�! �s��-�� t�$g	R[�	1�Sp��(P)6�B�Q���g��]�rEyZ�q(�Rx�:�N�@2}��A�� m����pZ�b�;թ^�Υ+�  FL&pbP�����@�(��
�OvC	� �j9D�D	P�|���s��G�m�)�~�l�[k���E]��hE[7�-���]�t���R`��k�a(��O۰�t������5��&*D��&j]��ub�@�إ�ն*����T�m{�<<  �#�&*@A��j �$MT����O����
Q@=�
Q����K��.��D�T*DA��	��JT�(H�F��YHa�m��cڷ'�nT����ۢ���ݘF�Iq @�C��v�� 
�	��8��6a�D�(H�f���
� �Q�LT�~�m�|��Sט�Ҷ�q8-�x�9��x�9-�x���;`�4���_v�F[��n��E~�F[{��n����}I/���+����7~>�eC���<�/���@�C��_Ժ({��!b�]究CD�X�i��w�t�ح��a�tsu�axk��b�+oK�H=<r@�i�U`~�Z�)+��'�̏t�$�b0�������������������������������O�݇_�/A�<�2�}d�K}�+��pr��q��T�8N��^�#8C�=�[�"�Si���,��ǫ>Y��TӬ�����y��1 s�V�xi������3狈�B��3H. ��� ��GX.���ˈ�ˉ�ˉ�ˉ�ˉ������2���`��ڮ0Z�E�EEp�5��������lh~d���-��Gd4?"
��I ͏p4?�@�����fΏ�?��͜�h~d�������s����X���rh�����䤋��N�?д�<N�X[�TJ�2�����׶:�]_�T0u���^D�b "V&�:f%a �"Zn���C"7B	�R��\�"h��$�	h-�@����Z���'�
44��c)1++p^}!� p1��3ڑ���� ����Q�d�Hlh~dw�Jz�Y�����`5p��b�p�EV��!Xj�ڃ`�j�E`�5Vt�� t�a4��9?"հ����+
͏�1���+
͏��`*(�j;TI�%Kx�S��*}k��8Ւ����\m���#-6\QE���7ꊢ�ب+�������+��G����� ���pE���s�Ä1W�'[�
V�����nQh��
��p-�%gC7\Q���W�z���6R"V
T#`�!����AT+����R��P���*,�C52X=+d���X�0,Ȱ�kX�`����J�a-��m�Mi�t��XW�o@���,d~�̂5ffA bf �d  1W�! 1C
�! 1w�eĨ��8.'F~ �c: �6�2t�V+�,c���@�";͏�����A�"rl(��pC�6t�o�w��y���� �똺��J�}��nԯ��3*��>i�d�!Yf4������Ƒ��}�.>���G���S�z
�L��)H<��s��B#r�1��L�c� ȂJ8V 7u�~�8cj�$���ÿ���;٩��6>�� {��"����h7���}@�"lE =r�3��.�K���M|}�_G��&��7���/?9��kb$A�/��Z��^ޠ�\�r.�7�5�HN,k�0��0��q6g�x-˯�8��g76�$6�+jA�!�W���C�����j���W�Tj�M�W�85܆�+j<�n��%5�:�4"_QC�9G�_QC�9��_QCI�Cz����T�!}�W�P���+j(�wH?�5��;���J��ayI����!ݖWԐ;uD��5�N҅yI�b��#�JOҝyE�ѩyE��i�����zr(���|�C�)�����!��W�PZ�&�+jXZ��py�5y|��_�R��;����!���﯏���4FN�Ţ�}������gx�<�$�?��Oz�Sy��\��N?��O���Y�dO?��O��j��;���?��O~��x'^���Vj�T�}��z���W��g��u���-�.�?\��\��X�x�t��v���r����\Ô�0��z���0��z��z���T��T߸h���}=�z=�;��5����V�V�k��k���Em��;>��'߿=�G8���O��K_w�s��=>}�?=}}�7my��o��8��^�uQ��X-u=x�hգ|�ϗ��E��?���(����k�:޽�:�����/���S?^��<}z}z�[>Ȱ�Ҙ��}a�~VT��~������S>��kѸJ��.U������C���ۻ3B���:a*��>}�?�o��k���痧 �~�����/?����^�O����|0��r�����?��`�y8}���Y� ��Ij�)�9���U�0�T�4L�k�>N���^���s���mE��C@�,��a'L�I�>�p�:�탖B8{��|�;5t��e!��9�P�Ro��U��Pv��v�%X�r�����&[=���N��
K**�1΄�4j>��M?j�Pi�G/�ُNo�g�<���K� ρ�s�n`0�Z�����@f�\-�I�P�'�6��IV�\���&�_c��kN0�C9qN�9|Ċ_����\�J���6����_U����f��G;�7-��@�ؑ0Κ�a�v_���uMU3⌷o��r)����b)�𧙦z��XU��R+UޅM���*�%����<��O|yT��:֋@�	r�{v�vm���ՙfP�ko\[�ڋ« J�6u+E۴�ܔDr!����$���J�>����
���_-����N��r��q�K�D��x��tP%U�6�9O�{�D�:�>�m��ں�7�)��h
ݎYr�
�k�M��� �);/��4��\,�$'��]����`=�1.� h���rN9NT�8��� (�0�drF�TG��"�6N�{�@���nhU`��,���>Ȋ`W[%jٖ�W]��6b�6PR"0��#�R�7u�{�UM�kUn�(�Yz�e�@-�*ٽ4se<��{Ѽ�M� ڵ`BV3��6R��o�����Y_2WT����.�hQ��Z}��@%��@Ks�90>d�w�`�`���/��#-h�o[-K�7�K��J��C9��,=R���X�#���GJ��}jd��bd�@��*<ziJS-�5R���K�T%�1lL�\����F&�9yc`5"mpv�2F��G`?kG㺴�4�"�w-b����hk��!؍��u8)^J߶^f���@�-�ܤD*���uTf����I��M a����&����^��ɼ;m��ż�r�!=-�d��M5=���5&�n�gA��k|A48��"�f^d`	@��=ֈ�3�!�プZ�d��m��Ծ�۾/t�3�ʲ��D���`�H`G��j�f�-|�1���GY.BK�?��Y���ϛIg�{�H��?��M8��w(��\ߜ �Jz�6�|�o��+�!�� N��ڀf��<��J��v�Ƽ��#���h��G��ɮ����xe���?��Y@M2=w@�ڬ��V���	�̨�o����3��6꧁�t\,��&�)$8詁˥%.�5.�8�+5έ����41p�O���@�X��=m�B��~�y*2O��1Jw���� �8�)��n�-��-b%��7_���b,�)5���O���q�?�-x%�apy>/�6��Du��������~���o�m���ol�t����}�g@曺��*d�.�
/&]j�tT�������o�ζΜ�YV��'��o��s����
W�Yt��(2sqJRdW���;�I�WJ/c3[w@EeV���;��_�����	���æ����a�ք�!��`��%��˛��K�]??��t󳵗�GYo_���޺��d=�������g��8�ۗ?��4�f��|��O1���ۗ>�ְ3�7@oV���է+�7�/��
�y ��17�����T����%�$�Y0FSkJ`6K`%��ha��Խ��l�`;;����O7��h,VU���_�����9��,�n���"��K�����z��_O/�h�����������݇�{[����r������ꦟ�.8�����((��t�R��眤x�3u_��>�~_��4�����3R�c�~��ϯ/O���u����A�3����G�C�qff����7�f����~\�`��b�Vg�H��.e)��fF���}ǆms��;AG��9���]@�N4�ܘ��M�9�a۱*�|����~i�4��f��9|�v��m���x�m#X2a-n�D�vS&����u���?aMLn�A�vSZ^m�	��㶷]��A�n�CP3���N�myhڲ9�ǩ�wj�����YX�st#�
&�,iΏ���GN+�����dFM�u�������k�y�8j�A3GP;8s`m��|� ��F�Y� �����陼m�������n�=X϶[q����=S���x�[IX�m����3r4�������W��f�ti1�0���F����kJy&����2�2�3b���Ib���
uc.�ړކ�p�n�ESnITg�o�3�e��8)�>�7ҏ0i�eJ� ��b6p���l�ENcL���dnkLeu��u�ج�m�-�m��yv)>l��I�G�L��9�#��/Uf����Ȼ�=�<�M��r��6OLƇ��Q����X�|�.�^@[.�PW��v+3J�e�����aZo��|��a({��,*=�����<�h��W%"N�~ �Xx7�zna|`�`���Fm��|F�rA��ڲ)����cG��l�(�X��vط�j�aQM)s�G��=.HR���l�qU��ؒj�Mo;8�a�o��Y!<�����X|�!3{�q�KȻ�=*�b����jX�-f5l�0���T��=rz.63{d�\�U���*�xKz,�mG>���0\�xU��)�VI>������bq�i:�F&��GU��<�) h^����12�,���ڲ1�U.�1��Q�05ϫ�A(cxѕm��12*!33F^�r"�R�p�Ę�ھ Z��� \b�w9#c-�� Fzm���"E0�*��m����m����܈\@[���Fd�A��Nq������R��y;��KȻt;t:�U�����������'�<�)����]��#�T|���J#>e�kyո��T����p�|L�;;L�F��]�$2uG��jN�6���^���o��u����L&X�*�@���33����wy�a���~{ q���U��[_��9[�wY�������$�e��]�$TKˁZmK�y�,|�$�C� ��j�c�"�Ж�I�� ��>�}cL�8O`?�|�`&pqպ��v�ĩt��2V��=Ϛ���ʼȻ���:�Sc���y;���K'��Z!b��ս��$�������I`���.g3�4�,��SW���qh=�w�`�<��|L��[�#^�wE1���o�L�XmK�����PIR�Pg�����=��Il�^@��&��Gt�X֋���R�RÐ�M����ܝ�A`7��2n�kH��#j���{�0�W@�|ފM��\`���f8����.2� �q����W;�a(�4]k���}�Em���s3���<v��d��8G
�k��Ҍ/nde��ځܑX��\@��-�R)�[È�ȥ����Q��� �,Z��/�-{\ד�W��X#n�WRw+�mf5gjGv�9��ʻ�ei��]5��.'YvǂF�i�U���*&g�Hv!�9_�:)"��-�Xd1�()���0�I�' �>}��������������7_��y��}�o���O����?���:~�Ǒ���<��}���k�������o�PK   V��W�vh� `� /   images/360150f7-d3d3-484d-baeb-b64063d02086.png�zUO\�%Z���kq9+��R��
wwwwww;8)��]��;�d�?L��Nv�œ�%��� ��@� �,-%�m�����n� B�_\T$E�jg�N��Ƞ�ńՀ��=p�v����by�u}.|�ǥ�Dzh��YщScǐI)+	3�!�xu�(�� �S�aPZю�X\�����]�?��I�����}��u�fW�<��̰m�x���'�����_|�~/���H�eB���KzpBZ����#4��
<T�Yį��Qy�?��S��t������Sم�i��[�s��$��պ�v/�r���.Y��˳&��G�����Dԧe�9��ܽ�����&W+K���wU�6��*�#��iə|,/����/2�2�ɥ�:n:���-}��e�[^H��"��o���
$�3�Ɛ���[�����@�!���7w��9��%��YlC�Ah�5�r/BP}��Q�Ӷ�ʁH/i �%��7]T�Ǿ��� �3�C5Li�7!N��"?�O�w���.W��Ƶŏ�x�p>���VH��}�}[W~gO~��~s�;�>`��c����V��;W�z���Գ`#�'"ɖ�Y�r�:&>y��]��M�l�'tk�&�v���m��w�g�:	e�<JZ����%u��n�o����R��" �nz�I`�t"���S;����2����kI�l@�r�-�[q��%b����Ԭ��r$K� <�R����;e���t�zm��i�xX[���E���Է]�t4R�U�Ӆ���-c:�pź9oO�,Y��KV$��M���,�?3�7#�lcU=�%F�����,Q1�� #���%~��[�X�Z�Q�X'��?����I�5*i	PzA�[�8���x���C�6:8�a��xvc��k��Ne!�����9Ϥ��V_,
�	GU�S�Mt�F�2�����db�zN�Hf`J�O�Bw��g���5�����m(20�í�Tp6އ��a܍��!+W�q�/4�܀?J��nd���̯f���MvX�.��l��Yh�z[�������ja. �ߤ���ρ�^s��Y)c��Kg����B�]��)Fu݊E�"�g¸�X�h���x={z��Y����-��_*m��pRq��w �vΫ����}��ʜ���F�f�/K�!:ę����U��x6�l�2�&���*��Z��r�X�xE:*���b� �"�RJe�D�j~!�Nb�\�Td��*��v����Y�� D3�X��xJY�z�{�LaG{�4��c�H-�Nn"Uϳ���"��O���j�a�AtO���M�?C&�5�4��dǃ��������Gk����z��>/\+
6�R�C���@+Gt`ɣ�6x��3�3]��w����8/d�[yAh�L)ٿy�5.Q`��]��?ߜ}��l��{�;0a�BT��K���Q�8ɑ�c��z}��S��w�%�Ʊv�Aş�խ��m��$t�0�B��OPp�ϗC!;Ҹ��I�����z#-���(�À�W&�J2�|� ��k���tO����{�h�w���F[W�ݜ������MW���$�KϽ�T�G�UF���V_,�n�\
�lJ�r�zڦKOCb�40z�4a���e�1g/V~��r��+���	ή �k�\ʆ�w�ښ�M������h};�?C0�S��W*�����461ށ�q�����2�(?Z�ݾ.;!�<��N���Қ6��RS��7�}���/V�B��̬-�l�M���ի�i�|v���D�B�c�g��\Ĝ�%fݴ�\��&�2�
.)%-��i���"bq�] �m�q�M��V�EtueБ(�$�w��8�X;#?���ώuf?��U���0[�E�b͛l�*�^��>��/($$ԾM���
�4����0�eg���d�l�s�i29�J3��9����d&M+w���:T~��Ѻ�;Ӎ�*2L���EX�9�$�5�$f�����VI)fs�.º%
m��'o�H��'o(�w�'~iSYZ�}�A]s�H����3�6��Z o��gf��vr0�O�pK!`8��狝_�ӝ��-@x ��J2�|��s�x�E �c�i*'#k�������ƺ��e�����,����֊z2��w�V�_�Q���rxUn���.RrÒ:���;Ǆ� ����$����d�St�JǴ^ޏG���`"���� �崗�Y�t2D�2L��p�S��6���{�d�HF�2Bn�V2���5����~�N�+�Ѻ:�����`#"�A��OS'$�]X����^޽�.�`�����=��|Z���j��5��Ș��͙�c��|����1�$���|v-�rc6��.\7Y����&D�����5��z��%����?9�n�kg�.|8qA�P����Xդo�2���;�%��*+�Zw�;��r��$�Z�qu�C�5�c�-<RӉ"������C���B���Љ�A�b�'t˃��GZ$�jl�G�V;����v�-�RH��$�x��6��<���a��4l �VgT�DU�3˰�"�p_�^K���w2�8�#��*�IJVv�[B�B�|��A��W�M�fA���*V)�K)�q�)�Mn]��(�X�C���2U�G�?�Z3�24B�+� �K�ǚ�О6K�K�:�g�@�	�����?�/'� � /4hިHv����HR
(�w�M�	���xfS�Ya��w��vo9�l�hh���޺{�S�X�^`�3��X���0���\�3��&a�Z����cFPC_'��iI��c�#��%p&û�B$���]mr;�{�˃�%K���#z���̃y8O�������v�Z���u^A�&m7��ݮ��ܻ7Ыn�g�vp^�a,ƻ.>>�m.�0�r"�9,3V^n.#������_��o�2+��BV�ΎIc�ن���!� ل2|C��ڠ�;�`A�v
�G\�5�e0d�sz��'�G�ɾ
�-x(΅h���O��9V����N�,��@D���ʸ��vdQ��[m�l|p`�;�~&]O|�8�~��z�{N!t�t'� a�6O-f�d� f���Á�.;�ĸ![&©���J	��G�'��`�(�]��تp�S4�e;a���腝�0��ITT1�4��� �Ȫ=Rخ%5e���V��6��E_�C�Z�{�n�����}ͣ�����@�ΏDF�-� �k�
N["Iח��=�?�pa��]--faCVm��:�Tk�����U�n`�(d0C��+b@2��Bm5KXj��qjM�ۄ���"���Ā����"Z��W��bI��5Ty���˗����F\�3� !�{�V��JϢ�[�sn�No1Zi�Rs�[��j�ҥ���(<�T�ģ/$mQ�ۄ?�������f�'_uI���2�::�=G
#�bݼ+%p��LPI#�W]v�Q}��8�<J�7��=K	�0i�C�1�� ��^E�I��a�������� �-
Q�������~����I��/]袵�A5
�D��5��z�{��Є?1�S@�d���d
/�e�'��C�:���+�w=�42�3�`]�95��2�@�[:�s4��
�f��2c���t/�'��i��>S�X�	�ً� �l��f'=�8�iJh��bl�G�8�j����r�'�����f2�j.9_��B���P��M*Wh�s��j��K��	���,�2%c� Ͻ Ve�f�*�?�x�?3Xo8������3����$���uj�ЗL5%S��fԴ;�y��
0�j��-U���Dt�ȣma�F�1n��r��tɶ\UQh������뻰��%Z���=c$&�̊!M��R�U�DQ@�a2�;Z*�0b^Vuxx�Rbu��y�h�z�y�><7����h�	�|�FWWwecC,�l� NF��1L���9�-��Cg�v����e��~���2D�5��VOR
�]�As�����@Q�_\�EA8��g���Fp�2<�3��"�KVV���%T����+b��wO4M��
Ǟ@��J2���9*�B�� �׬C�e���>I
��A\x�>E��NA<&��@�$}��u��i���>/�i��9��?rI�Ye�l�o�,�Y
��mf����{�t	��GT
�Ϗ$r�tGF�ʣ�/ڦ��4Ԣ�N�Eq����[�P��ɲmqN����q��EN�W���z�A�ȯ���_Nh:u�-�i7�6�Fŭ�^%����~J���,�ĸ�|�!<#�z-n�%���zx����*�c<Z���?堮[C�C��r�hȍ7�ڿ�I�ĳ�S�(0�k���"DC�M���[���M�x*��w�m���,�!���l8�@;L��0�D��W����ӅKx� ��u*U�
&Ѿmɞ�v�Wg��9<��e.��,�����J
�8gJ4���rnS�\�ɗK �g��^|W��3gM�/�6��w��yL9¤,(HA�V��Ƥ�6LTs�l�K�X#�b�yM�ٌj*9��gӃ������ۆf�~[Zֈ?�_SU�r����O��:8L���o�3V��j}�,9jJ��P�5V"=ת���9���%��s(0�ˇ�>��9 `7��e?���p�c'�D��O޴�1���1!�l��F��8D
D�,Z�%�3R�tˁ�ʪ���	Xi�;ۙ��.8�q�?�m'(�2҃ㅩ�fp�g��k�vB�m>B����'T���sȦ)�q�|#�i��*H"JZ�T��J�_#�J��h��L>�V��)1҉��X�x���t�֔�/21��r
���aYU��
>�_�`� �8�<q4��1�����-��]jPЏ7d�`ۜ�1���i!���u�5�\�8�F��|�����9m�Ƒ����iݒ��j���� ������!��htT�uۍ���<<a^W=�ד���ב3ʤ��H�.(΢�
`W�v�F����8|������~�,�82<�4ڈ����m*jh��V�
�_Q��\r�.�s� ��k�q'o����R��8T��۲�Z�J�TJz���,�Ue;�W�מH���u�5���Sɡ��� ���͊�$���_5�����6g��Y��3Y���э斴 '&k�#�R����LN�\y�h����q��d�� �!�ܚ���ex�٠�2�y�/xuU[��묝Uj�R�����.]�7N0�#��ؤ÷e���6Wc�̓����*�f��(7�H�L&�m޾AB7���C,bف8��݆G�\#��yT(֦�:#�㙢{�te�`�߶�"@�����g�?���X�k�0����w��R>]~	ޝ�ɼ��R~����B�F���˦y�7��e"�F�	�XO�l�\�s�ks���4�j�4��U��"¥�#�=�R�}����G��[���A�n�T?��B|t�11�7c��׾&�\8�����m�֮c�N+B,�eݏI���<��C�Sz�"��%]����cޡ��n4IB��z�Q�ط�,3�H3�F��%)h���}����n��ĕ�'ѕ��]Ӊo=�JHR�/���C�r�sF�����7��>�ߑcX�P����-��
�L۲ �ݗÌx��
5v�pI#���n�l�I�sO'�xi*շ^\��+L≱ԇ�qy�ҷ�x�j{`a����`Qc�� :��S�1�7X�y���*��&m�X�o�p�f��K�aP<b-��a�^g�1��M!��pm��b�f���|\�0P��l�2��;�*mj/��nm�U{��TOM�CZ����q��:�t4�ZD�lf�p�]KE��B�-k��Em���h�\������HN��=� �вG:Ά�]��~��qa�+ʡ1��D�%��_�ٔ�K��#�Q8�t(l�d�4X��Gn��Ƞ�`u�%:I@�ؐ6#i�8jh]i�
6ONӯ��Kw�O���Ȼv����<�Uu:�튼S>�0a����T,靟@?���ֵsĩ��j�+.f&t�n˦�9�S��a�qy��߂�:vKD	IOx���� ��A8~�F0qs#@�;�������@��XoVV��Bdn���3�����J���w��7��{
d3�It������RCIc�P<�
�/�HLP��Ԥ����ꨌ�����{2#�Kt	�,
!�H���$�p���i�IR�%+�<9zG#��̯o���!<�u�Fx��>���JD� J�oB6�mێ^�o@�7����!"��Dϡ�[J�����/��������c�5x���<+�ceV�6�`�_U؅�ȍ�Q�o�o�g��eb��-��,�pu ~�x	������E��e��e�Ob��i�3�yi�����Z����`�_�/�.qj$odXa�h�%S%D������N�����JZ��
�":��
t�չb�������i�k��|����Rq�N��9fI���.<��Boy��`"l�����8�$�%kC�*ш�'Jh�"��TI!S��cVX�"\���~�}�ŕJiT!�"�ڨ��}76� ���p.A���H��j�Ă���J��*���FcI̟1����Ijf33Rm��촡���#u0$Ǽ(��I���q���L�4���̂x�'�j6�l�T�M-4$�j]s��5�ʸ�=����n�����he��߰BU�F��c�K��*S����+� ����y�odK���-�;�X�����L���V�/�"�vKv_�H�~̡j2\��PAm�l.�eG{��N���^��v�0�j�~�ֲ�$�������J�p��d#d���#���L5��ܸQ�� �C{�ZU��+x�t����H�7�%��i��C6j.���k��r�;zC�,���4�JN��b��F��_o��"E�$��˓�9 n+{4�J���̀G���$ry�t-����+^��햎�RM�Ğ;�ud!I
��kU�H�
������5�e����QCGo�n9b��/�PS�v��R��u�7#�O2��ӛ�F�$2��n�;��{�/4tx�qg�D�W�&OO,��_(�	�����#���9_��54o��	PN&�g�'��j	ߐ�zf�J8��р�{f�?��]���Od��Yd��g���}�Z�F\%��9�wM%zF�E!�A�߮�=w��]gP�Gn&��ݭ� �.G4�P�Sq<�z�� ����Y�#�w�MnR������h�k[�G�d�0Ե��pK��d��X#UQ��\v���k��E9���Py7ۺsTW�>�ֆ��#�ԭ�7��-NVE�6&�-G��.ɑ!��X����,Ǘ&��z��s�Kd>��U�|Wa���z��~�ǧ+����θΞ�X�7sf3G�I~7k�\ :�D�eP�rm����PD�V�6pY�u��(Q
DG�Va�qS� A��~��U�~�O�~d��h��}��j�}_�2�a�K�d��lt�iD�F�_�����T��}�������(l95U�����c�L��˸�5���	�g_�]���q�P��������nd� Q{�����I$�cJ�z���l���x���ӎ�p떐Fg�48+�����V��o���{�����Xp�73#��͕@��\;ڈ��sd*
GZ�͊����|�!�Aa`�ڴ(�Q�|�[������AY�%�z��a�@[U��:�ퟥ:P�
9��*N�#�Dr�M!F�,��Y�h�1�@S��J�c���R<�K�&�!-���/�c��H_�X�m"+=GX�x�](��:���L��A"U-PC�pN�AG�ūR���{�)G�P�H�g5S�m=+�5��� ���x3��7��3�9��J��0x�
Z��D�2j͡��TήqBX�b��d�����,�(�q? 6��n�5� �f��z�$ފj���L��z��H�9;:�}M�G�Y���G��af�\����	�X�F�DN )!6�Z-�u����PbWZ�)k��/V�8?V�&f�'��3^�݄~ZŏO!/����n�(�u�M�9+�d#�ȵ�b�t%>S�w�M��(�Ķ�8������+k��y��f��ȯ?3���[9�]T�(f@�
����U(%^��P�oJ,C����	��s<꺃������p�le�����4�H����i	졁�j������O=�?Z�<�(� B9��f�=�C3+k,���&�Ǳ}-�|�>)-%�&�D[L��Qy[��ΐ2V����5�j
��/�.ѥ?p�� 
~��Y-T;%!Dqw�u'��N�
k^�14��/���7R��9�����=�����	C��RىX��"g����'�0�*�&u<�53�9dHu��:Kr�A�:�����jٕ�H��"Z���W?b��.Y����zkhD�p��Ӛ�[�*s��R�[4�W�DZzZ�-*o1�౟�+(3%\��\6�"1T�&TFs�I�!S�k��R����r����E�7~>��ϏjEA�XFȆj��d�BI��_3Q�,7pU���N
1�90ڨV͑.�Y��ۯ�������R2��/`ȥ��n'y�S(dTS\�A��MK1�^	�l%kfpo����ЃDNdH�$��VF0]�y�s�\�pqV�i��ްR��q+h�'��vTh���&
����ྡྷ�gM���8ntKh�X����b�5&�[�	Ϭ����R���@y�fg���Z�Q�AS�
s��Ja�Ei}W^��$e�.K/��k�{��K_`[�F����R�O��0VV�o�&�^�/>?�ե(�X٢�i�.�#i�0�SÍ�_���3���CC��5�|y+h',VН5�`Z��pw�&h�ݿo���Ck�݋�WE��=N)f�^��x��#78/���qQ���	g�����MEO�s7Uq଑�G������}��k�{Â@7�ՅՊ�)�|�h��
ʾ�D�$�!.����'�;�5�\R?PF�ʟ���uf�c��ɻ(�t�K�g_��z�y&_z������$���H]�k����ѭ�McMx4�'����j�յ��;�z�W�uW����B�ý�vO`�r�Q�� 4�q���!Gg���}^	������,����~�5�Xm~�BhN�/���,�/���ù�!T�	���S�՞Ō��@�W �������i�̇P4,�t�KC��؅�����|T��jML{@*�we�ҊM�e��#���+PX�������Z鿱F\g��7�'��V탳�}<�l�X�^����S�w���D)���?\� ǆ�A���$���~s_Ys%o4)8`��P��_�~���4�R�7*?�7���&��5��FߔӞr'�=mz��L��� \�"����0��L]�m�L"ށ�X�jU���E��6ku��Y`p�C���X5V�x��<<��",)�V"7���$�ʰY� �
���{�zdb±���MM%DK��(%\��Yێ��cxvZ�F+��(:�c$�y��Gr�Ĝ�t7E�ӈʧ���STC����~��0��ص9�B��B˩x���lw
�7Y�5V�L�6՟F�X 0W�C�N��5���%2�6�&�u��|4r�h��M�L5�ғ�e|iD��L�ר�S�"y'���k����u���{HF�	
7���ɍ�{͍��?Hd�	�D1%����'��{i�$�jYx:m����]?�MJ<K|���ٖl��ۚ�CW��b�z�3 �b��4�����E��FZC�^�~`����6�_����o���!�h�ד���)��+����u��Y�P8�+�_F�Ѕ?���`������C����0�a]-���/���s���d��]rc�6�<���Z�$���y��(�yH��1�����p`�f�(/j��p�d�Z*����5頣c+�|�GC%'W��&�ۊ�k���j*���d~�<L��%=Ή_��}Ζ0�"�s/��i�Ti��"��6u���V�3Y��\! 7ä0����6�S1q�4��Fg7pAa�k�!
�U�ѣ�%�^a��t=v��W�Ik�`/f��xt)�r�k~�I�_,B���T���FR6&ALnd�50w@=NY$�eɲ���I�����cQ�'�Ln`W���(\7���[e��[+���/�����VϤE�A���+yJ>Z&k����M��1>�� n5�}�g�d"h��SW�Rp��m�z���~�*�5Ud��;d���4Ǜ{���.�.�̀4��ڶt�"�Mz5���q�j��m&ln�f�OɘP�~ZHu�_z�ݠ�&�g|�����]m�)J>6�$�}2u�.\�^O���*�z�(�����l��q�l�}�;�:�����T�a�`{2`pwt�N���5釐�|[�jv��بF�:�Z��~�đK�h/����K���W�7��(�8Y��4���T1�3��c���|��R�sx���uK!�.ϙY�o⤚���PC~��K��l@���cE�&(q�=6��C�������?L�H׮�S���E3���_�.�s����O2S��;���NMP�N�ܶ�qT�5��8��K�@���%�B��:<�k��	�{"�Ѫ�k0�k�����p
�C��6���,��w7ȝLI�v 2�(ˎ�ݥ8҈v�X{mh^
ѵ"��r��N����+b�` �T�˒���HW��"7�-�1 W;���=?�
��]	��������������o�^���7��]���&�dZ�"Ő�:�e+�^s� s+'[K'�~��.�֜�4`���믢բ�5�״:�ѝ�@�����St嘼�����:?�ˎ8C�s�ij:~���U���:����jAtL֢�o5��T��Yr"O�dr��|�?z�ݐ��B���z���j~�Dh�&�{����RѺ�tnM,*���N<a��4�v������0��R�uW�y��)uc���%eyp��zb����#�f�_� +M�s[��.���K#�F�U����fUzbդj�Ld�*��2����q�	W�z�4��(xUA��e�ȂbKS��K}~��Z��a�Q�CF����wքO�(��̊d�Ǔ8����`�.K�*9o��39��1�pf�I4��F�!?ڕ+���kZ.�d5x,._R=L1*Ui]Nû��֐N���
����ݡ��KO�_�Rn8�����ҳOe��Zͫ�K����4B�JoG��sF�}�V]�T|Yh��`��4'e�_���W�^h6��!�p��r��2r�ӌ��-<���n�����}z%^&�=��z9�j�[�3���7/�b���wIpo�q���Y�Ƹ�G��Te�(��|�?��#%I����w%���4�N2���~t�y�e��u���b{��Eõpb�E\�ߛ`d�2�F��f����QNAd9,���S47G���HU�I��������Y -��`����z�b6�:Ka��fV5\�T}咛��黃y;��0�]�c�Ǧ0-t������u�ֿI�~lz�ܫ5�g�%z�b3]
⏦jޤ�������f}�`�����9
!���z+�,�������/ܴ{� dt�>������]y����)��:��%��?��|>��C�@��,~�2φ-�*�B��\������Ⱦ�N�z���E��ՆDm~ *���)U�CB[�0��[ԋ��<��eN�c$
�J�wu�r��k'rM�9�M�
�Q�+�#�X�[���Ԩ�W&_�=��#ͭw�lU���I�Rȿ���Q�1/�Pi�.�e����l�ɎA~ ̙����X.>���`�zk¾�W��3�nPΈ�TK;��Ң-���a|��A�&,�˧�.L[Le��f[[^׀���s�v��iD�
q����jJYL�M䥳=y�W�l�K�B�F<
���|!���w�>������7���W�T��_J)�bk��b�I�(7��}�׫�E(q[�6Μ��:-�C@�z�'��a�O�e��.-�u�
cO�/�8�?5�5�58���ۏ��8u����3y�dƏ�=��,헹��o~h�����\)i�it6{$��o]t7IA�K�Ύj���j�"����.@�۶�dx�q�Vi���MN��vU1���pd�W�Y�4�6��y�'''˗	CT�L�`�GUĚ[Z",��ѓ,}D��h��r����#�[߯�(�gL��q�	�E%K�
�쀅�������4�vF�n�y�c����$f��n��j�l���@]�A8%GCռ�^P�ww�����fJ��/��M$jdb�ѷ��c���,��o�9;-/-!�%WP�~�W��ɇ^����sg>��ݜ�U���	Rk�XPXu9��Xf�:-�k���3���t9�nxZ
�s{!}��C:�Ak@��ѺH'm� ���it��sJr�S~�D:�\R%�3Fb���$Fn0j�a��������m�7�'��8������1���dOwG�i�
�DlRA�L��veJ�F�7���8��pi�.�����,��`��g�!9/.;rͶ�ך�:#���xZ�e�0�2T�u��ʿ\j~" �S�����߽��Ǌ��˖�/����+�^�@WCkCl��h����Tl�������n��F��Ô!��Rl���*Tݿ\�(�^���oiLI	���~g[�	j���p�f;�7mNT={��z:L*�9��yT?|������r���h5*O��2	�?6�7ky���-��S�jT��4���U����S��L����#��)ᚯ�7=���|~�Osć���	�;4���G�i/���U��W�ڃn`�����EK����E b��7��y��X��i���;7q�x�6sW�&���e���2��?��7}���/����L�$��գ4��f��|f</�@ߺbI��lIS���v("�3 ���߷{N�,����ɲb��k.i�[y�i��x�mJU�9/=�����ޕ�?��!��ݐ���t-b��	�+�!�	��cD���Ά�������&kuD=� �Q�V�>\�Q��n���D�Ig��w�`ϑ������e
�"��c;{�{<�������Տ�\-�O�Wq�<���b��T�Uj��j�H^OS�Y��nvLɁha��#"b��֏6H�AɨFk|�z	��?����J�v�������qw*-� $�7�9o���F'))?��f37#�F_�W�>��'8�'�O�x�����9��Y�A�z�d�$]�"�սѣ�މ�g�y!���/}���}�+J�\*/��C, ⧍��t��!G��%k����}�^=7]�Z4�6�B0q�T�U��9�c��ʐ�q�.	mz���sBL�`�D
w[������V���H�Q^Ĳ���q��{G�>��*��q�S;��'+��>BT����	֗�N�ڦ���R��4�[�#5�C�vr_l�����b"���r���ݍ1��*+n��(1�#����a��_"���7�;]�py�2��^�P�)��Qɳ�Ž�U�d1�J��S���xXԵ�7g.��h�3v9H*�),�׸��z���G�C��8����4 �y�w��@���aȏ�>#c����W���>�r5/�O&�Q��Ņ��zwH����G��6��I���\\����#��܎���������-����.�#�y�4U�V�y ֜{��k�%����/5��������h߮Xx���Vz��+��`��rL�e����q4\�9���2�O0�H8ЄI}Q��{��D*C�$G��_���B����/#��������lc���W��q�O8EC�������<F�S�'�ѳ���Ѫ7�W��=��&5'8��(�q��M��(�7Z>��8�n�����2v8����X�2$��s8��T�#wyT��D�ܗEڈN�;_ؠ��*x�v�qy�������z��
�_��+��[����c�n�%s�o����7�={��}Ki�� pR���ĵ���濹~2�0BږFϔ�~�͍��?�>v_Bk��S��"��H�'Y*�چ�u�:x���W�Wࡀ��|���ǀ�`�D	p�� ������Zk#�W��p�e�i��i��v1���OT<+)GZ��?�=3�Qp�%6����*�
y���ۛ4��S�����hi#��4r��×׫�&�	���
�	*����8���l����x���G�{��^0�?��b�f2��������"(��Z�T�KT�҆`�c�Iz�օ����%RȒg}3ŕB�#�FJPG��7��ܦ�џCQ����^��9r��<�@(���{5}�|� k���$����p�B%Gg:��l�ⶖ�<��Z`��h[a�ffJ֑���gn�<}.�ݔ����d��:�Pf�;�K+BA�G9��s�95��"fA���M�u�V���[�0�+:ҎP�H���Ӯ�o(�_fx���2A�$�t���^O9��ݍ!^O�v��E�-��#˽0���DM���	`X�R-`y\�����g����t5q�)��!��]��]W�=3aV�"??3f�݄ ��$��d�8���@��w*�W|�);S�D�:���P��5<�?�&��P��s1a0̈́��*~!KV�f�����\qz)]��/��9\�s�����E(�M�!�&-���&[P{y��9��}w�s�{v��W���\��H�i�0u1x�d�}݈R�Z��icD˿�^Ml �IS�
���fv�/�hE*6�-z��Y�������C!֖,ҾG��D�P��i��C��X��'ix�$��9J�"l�	1
#���m8v�tz[IxŸls�-!�"���I��M�&t���`�a~VQ�<la�fXR��e�~Q����镮�^�^�gK��Y�K��罢����譤X+�cD߶�����2)�{��xzDA���0�hh��\�p�ʥ���ͅ����g���+17�A���`q�Mq^:����������Y����͛�O��������f��ָ�]�����������ޫ�sd.DnS,<�x>�Wl���p��I�7k��9r�GZ^���EL"HH�2yU�U�-q�4�~zD�	٠��Ϭ7a�}<��SV���\��11_���۽o��?=DH]^�wFw�9r������y7/��	�aӉAH�O�7� ,^��q$8�g|�,�J�N��M_G���ސ�@>�u-g���es��Mƥ)�S�$LT�';��Y�Q�cj�tT�uI�N`��]�m��e��R#b�!��9:�������Q��5�N���޴5$8��˖#C��3�^���m1ӃZӭ-��'݂�;V�z��={#����t�e���/�����z���wq�n��r�>F2�{�%kŒN��c��}�>4o��<8W�ıh.�?�᩸�E��~;�*Hd��,|���}g�'�Cr:wy^l��n�F)��W����b`����v����#4���׽촊$�O8CLjE]�O�-����=��t@��%�SL؆M�vCr��?o�ύ|C�c ��Bޛ�ۛ���'�<K�"�O��2�{���Q:��]�δ�'�/�=���"��Ё-^wJ�4��ԇ-+iR欨wP��>8��PM��Kɪp1}�����	Z$���y*ݾ8�1�>��؋��7�X�G�f�N��n���Bc2u���}��~��NG����%��p�w��$^�vb~7!�='����?�{��m��hk�JzY�,o�"������H���ů�9F��6���|��}Y��K�͋yH�yb�_W��4fTB8{��o�h?ϛXm�"%��SE����TPnJ
�3�YA��SYk��>Y&)�*y�QoY0�͝�負j{��6&�G��W�S���cY}!v9~hC(	�6�όn ���L�a�D��y6��V��˃������
��5��=3�Re����<��nD�������(�M�i��Q>��	�D��)$@�!��ř��k�^7U~����D����é��X���[�ц�[=p�zw�NՇ8�{�W��1��CF�p�a������t�UW�JʶY��st~��	s�o��P;v��\㦬je[�4*T�T5��Q�����C,�k|n��B��p6����{�M�0`��HH�(`�o�Ѻ�~0�*���k���N��A���|�_�mw������;�d��S(4�w�︳>ȍ?���� �E�C`�w��w�� 8�A��*Y{M��*��q�T�0��/�3@̿��q߶�	z�k)$���U�t򞢧�&Dl�tIxofܮv����Ԋ�bzْӚ�RMb��H�$q��BZ]L��&Oa㽢*��Hr��X���l���#u� ����b��]�< ���ţs��2�M�!�ٹ�?x�{p�u_��}�å�x�o�c��<:����^��kpxy��,i\Q6�%��jJ��s��4���Was}Ip]�A��>
*�JEE~�K��~��H�*��!��	k��Ih�B���\�׿�����kaV��K^�K�|�f�i��ڏ���mPAC6'�^`��h���CxN��S��?[�+�G���=xSB��E]�Ʒo¯��{эr	xHcV�U��\*؞��'	9�gA�Z�P�CG{s\����F2�A�G�4��W>e�I�@ᡗ����+�|d<�~"�/U�"�����8�x�/��Xc�o�^0��
W�����=3x�{ފ����Y=�OW`L��T<=�9SS���� �u�-PG�Lz�<�l����yO{^� O�R,���</��i�$��38t��w������
D9$�|�s�`�x��/�����r���� Y�38r�0��7О]�8Q��y*����ā�M�,���=��D�nU},�]|����ݬ!���&fg���azj'����_�>������a�CTCv�ca�.D�ԓwH�S�'��rL����VV�p�Y����ߊO�K�>�s�?�Ԫ�#s�r���=��ؽ0��s:�𚫡L����j;�q�ͷ�s_�2��4��v�w#�7Ǩ�v������X���׼�x�%gbm�t[g�bE���D�jxASHا?w-��� ����<�9W�wށ����ҫ������H��w������n�T�����}G���t������}�tԏ{=<�iW��\���҈ti�:�-d�XH�8�Ts_���?�����+G�+o��	��`.�����Dz�h)`{�_9�t�^[��8���`��"/
��u�>]bۙ��"K��Y����o�e�^������Е�2m;�|b��!���W^�*\��K�k�\�Po�HO<Ε��6VWW�~s�;���;�#�7p��p�=ǰg��t�?�!}d�輳q�ݷ!`u��g7��ɾ�	�� ���Q�Qi<yV$�-*�ҳ�( �wf�ZE{���@�IՓ��6%�M'��}�������_�⏖��c9��߳�0%���9x�o|���8�"�4���PɈ�1���<���Ϲ��ӏ���.��������1���#>��a�Q)<)n����R���I� ʻ|�%n�t�1'_�d�jG������ ����L�^'�>���'���H�B�&���_L�u�їi+����cN{�`Q���+���*�%|�JڐP�PM���� ��t�����y���Nރw��\���������,Ӈ��zߪz+Ǯ��=ӓ�$#"�d
�aqŀHte�+" Ie�i�a��a�����9U�9|\��5�����s��;�uΜ�����繞���S�����+�+�L��"�Պx�)6;����`6�����4�4�Y&�R&��?q�>�ti��t��~3s�QO*W�$w�?�{��z;��������A���]1��M��u�Ν���B0��
���ŧ�d�L��O_�Ԛ���EVmh�ZA.��e��?�|�1>2�]�4��q:�x�#��3/�����#DI�2Y�8�#Dbl[ЇZ%��9���K1:��!��>ik���)���������+���*l�6d�9XL*�f3���<�����嫯���0�V�}��*�٢;� �bY|�+�"Ul ��A�����)�<��]>��-�#>3	���Z]Z�V3�T<Cux�Y�����K5���c.^�#+��Mh��U.��98��'
��4V��$���dsоÂ@������{Rٚ�H
�6[Sz��pډ�/};wl���ť�aE4A�TA[G'2����r�w�*PfF�ho-�b��7�����MȤ�P�Ee2��葪�t&'F�K��?�Ͽ�*� JM�)��.�7�s����<�6U�Y��X�Hg280|�X}#��[o��t��/�T�'l
,�>*�4ڼv����a��W�`�Xomۊ�y�z�_x	^۶O��IZ�* ��Z�j-����^�i�v �3è4˰�58�n��n�43�2N��Ͼ���ۈ���l���Ʉ3�9����LJ*7m�N��O�e�D�H�@���C"���O\���I�R9�%Kbj|J��e�����HE�p�-7ḣ���E�GO4.05�*����A% �����K-�������p	�D=��f�U�JE�z��O�`ppX�2v29�M��f�1��% }Bv~V�"�b� �+����Ypɥ��އx<"���s!�s0i�����|�+���߃�k��I��_'��sp84�Y�w��A������?�D&�EKWO��Y�N,T'�	nfSV/��=��� �S�Cf�Y��2���&ǹ%�*�2���J��r�o�g�����R]�	��`"���x�s�_�b�M�|�r���E����=a��1���x�������r([_MJ�Q�b��@�j�Wt᪫�#��q�Fl��&���(�<N��Y�J�V�8!K>����[o�%en^�����!�I�i�.�&,]���Edȕ�a�`2���WX��Pd4b���R�T��!��yr~�ԮC=���
	=�Z�1��,��$~�V�}���������J]"n���XTi#P�W�&�$؆���}L��b��=X�|��̜r���0�B�B	�~������0[Pj4�t�0�!f��|���e8��c�<1���u���t�ֳ����÷p�T�Zt2���F1��G��Q,��c��>�S����@��cG���#'Csz126�+�����ɯ1[4���ZU�7�8>{�'p�E����ZL���e��'6=�������܊d��B�w��l>�$�d363�8�$\}��L��a5�E����<U=\�N�.�T?|��m�(I�6
�9���J�s��.����E&ഛeb�d@��d�����ŗ��]Ĳ%(� �X1А�b� 趠�̓[n�6�ٔ���E�>�h��f��=���w�m���X�$���3��NM������g�x,RɈ���4��$W�m�J�p;^�H����G�E&/=S��'�}���W��o|���Lό#D�QUA{g���|����r�R9jMXliQ�4��dH5�5�v�(f�P)&�
lV�R��]�,P�%,^�����x��-�w��H>E4�
�a�?���S�RiI�齵s�nd29Bmp�=��n�	���
f;���4B��p�L8��c���X�d	�� ���p?��ߋd:���?k�:
������+���On�]lrq�ԋp(E|���qĪ~L��IS``K٤����*�V3"�.�?�3�4�g��������NC4�k[ސ���f��QR�"����пd	4
#
�t�[z\_f�	d�)�;b%&FG�0�8\HNO���N�wѨ��/&`R갻(*����h4j7�Zh�?��ؾ}+���?��s�@<2%���_-�/����*�Z�n������M����܌T��Ϧ���/�c�X�̛t�qP&�
E[�4C.�]�x�B�v�͈DfDQ�򁥂���`�vy�n��O?�ˊ+>s%������鲉����5�f28��S�4Z14:�]{����6mޅ���fW�0ȵ+
۳s,�9�4��b>奷�6o8�/�b��e>Dk����I
xl(t�}&���My����:���yԑ?����g0��W�?���_�����^>�_=򫚣{]SuI&]�\��4# t���9	�j'��4	�1l~s�yg7�V-]��"��瓀����9�R���z_����� :;;�͚1>\��f�"o��+��b\1��{;��'�ZNb�a�R� @'�]W7->١�Fވ����,�K6o.�{X���Q*���`�I�U�Й�V���G����CH5��g���سg�������(�
0Jխ�[���?!]��dhb.��j5�n��Nj����o��k��f2�j�8��u��X"բ���Ï=�ǟ��^L�b��6m�XAG��r+-º5+��������+���8����969����:<���Ū!��J4���@jv~�C8��ㄟA�*F�0���u��/���Ex慍���?C[{�'g`��(0]���A�����_��χ���y��d*.ו+�G�d�����܂h�(�M��!��B&s�
I�~�Q��ӗ"��fѣ��nwz�v��^+����(����1�Ȣ��D:Oo#fC�M�\*\f����J��xə�Մ4\���D0D�^÷o��o}Վ���x�R�{v� �����N:�t�}�(�Y,��V��sz���q��.��S�B$桭�C�uk7���r�]ai_S�<;3��'�/�L߸�;88=�t�,VM��B���'ׅ�b���$�լx���q'�-+��%��/��w3v�E����B��˪E�u�p��7©���
��wb&���q�TE"Q1.%������dM&EX݀I��d6��X�ש�K��,���ѨT�=�,��{Q(�hG�]��[~�c�ص6w���z�4E�Om��PJ��U����09y�z��M��%�+�}�ٗ�y�u�)x�����+���۠q!�4�ae%�X���{�r��Y���n�OK��nu���x*oȇl*�ngL�:��(��|��?F{Ь��T����|P�o2+����n������kW�������0�%v��S�s�#���L����8�g��RQ����%���OEz[�yi���O�E)�6��633�B.+����z#V�Y�d2.ti��"�&|0	r�ؾ�-<���غu#>�����H̔���D/�*�R�V�=�don{w��w(PT�Рj��n�^�4�\��0�����I`<;�e/�y/Kɘ���GQ��`r<�����\��ML��oc�F��\�����Th��<���Gu�/>�я�����]X�?�����������;����ŭ��%��)lE��`���x)K	C��Q,eu�&ۉ��:,ZżT�����Y�� ��:��c�1=N��lQr�S����&�31�c�5W՜Jt_1r��Z�����!Fy&E�D��9p�l�u�1�Zѵ2%�+�o<褼����~�/[�lU���T��j�Q� V��RR�Yl��v�Cx���f����=������+���pz�󆄃��177#Ys/n~F�T�f�Q��%(���D����5������E�������_��K/���{p?:bxv
����\���-�r*�(Ԭ�[ԋ��~�]>QFq�E�mh�b�a���ظi3�:�����B��D���炎�s#8b�r�v� ���h!�8%�]Ni9p����Ͽ�;����,�u���9dJ%x�~x\.4*�݇E���w���a��2�J�:s �4�����Dd
�˖c��}px��O�Fq���M!���e�~�ȴL&��n?��6�61Sn��>Dcq<��'P3���и(/g��Jy,�	
8)&��K/�Iҵ���@0��]�w������`hr�7 հZ]A�-�R;6m�?~�b�~�Q��k��*�ZKLYP�bEWg/��x>�(���4(�ç�mh�����|�:=!�+E�Rq9�իVb�%�}`�s�02A�~\�����4j5��'���W������t�y.������Ũ��YT������,��V���
�F��$�,ďn�~�^�W��2��p��q�f��O�X�e��C#�/B�\0��R=�M"�L^-�7ވO8�\QE��=��m(�s�l��7�s��N���@"U�jrIԙJ ^+�e��_���W`rjF�*٨t�ؔ����l��D$��~�S��163��HT@�����s��]i@m4�ؐ�D����ty����G$�G�\;�O:�d�RI�ϰ�U���@a�Q�*����>'-�
0[u~R��\H�?���xD���+8��c%-!�NH|۸�\Z*�l�3�H��I���)LNF015�s�4�Nϋ�T�4?���V[���U�8�G�IPF��F�r9D�MS�K/� ��!LM��N�tׯ3*�,�cl���Dd.�'"��O(|�����d�*Rc�.}�
�:֮?�	O<�<�Fg�e�nT�53�g�:�D%�ıG�]ۥ=�2��J ���p���r����,Wv5,L)!�����mN��p����R&ubhpX����O�Z�B��(Jk�{�ؚ5k�����X�oEI�ܡ�N��ـ�@�����'��������GG�a��ȝUch-}��%���0�)���a/clr>s����`��0��|C�+yTT�ɼ�[I��$��8��:����yr.t4-.Z�j�gt��O�b��?���/c��%�g��
o��M�=��d1n��ӄ� �~*
�#8�?�+!�J�C�|�$M�$��zF
�=D�K�l��iZ-î����h�28q�*���R�!�����~_X���2cll���7<�{��g�.���i؊����aL�aQ{�g�t����I����w(���n<��G165������XX��n�g�1��#���.��,BG�v�&����iX5��Kv��>	k ��h����
p38z�*XN��]�k؝~�Z�1_U���	毻v��;0��">opI��b.���ņ\4�훶�^d��J���?�M��+�db�\�~�lX�^�M�upT��d�{��2�76�C����S�
Vt��(5
��lh��b��r%Ŋ'_ވ��(��24�
�f��\D>��lX�v�Ua%�,i����m^���5��Ï�l4"S����l.7�+fzn�"�8v�2��,X���=�rI��"����@_g7�ڵ[�ٍT���x�r�LnՌ����a�+��w`��H�38묳��݁�}{;��(��Q����8��p Ŏ�a!;G#QE�w��O��1,X"��Y�� ��b��A��'��"�Na.�Tb�F3��T�Հ�������v.��B�>1������]Ӱc����������De^�F �{Ӯ�r��G'�ሣпh	��LV�L��r	�3#�z�	�ׁ^{Ǟ�A�B�̥Qa��YEOЋ��A|�����k��KO,�����"�U� ���q(>n��n�32&�V���z�	��~�Ϳ�5��D.�B1���G�l��ɹ�F*��Ҷ�F�6�Ţ�T6���+�[��s��������f�z�@sZP.���+ƙ�{߃���3?���6��$bs�ڶ�U�9}�\��5E�����q���f�]��LC���-H�x>����)i�	 ��    IDATk�jGnA
��L&�ˎ�������W㳟��9�T�J ��?�� >�����G�Ú�+�l�2q��������1
��/�s/o�+�m���,,���H��p�"i�&����rx��'`|d��TJ��E2C�u�����j���&�l�Ì�"o��t��l�.]�T�k����)������AYdF�����q��>U5׎;�ـ��m���x�Rux�)��RW���$TM��UiZK�Ҩ�MMk#�N�N��T*Ս|m�RQfs�^/�v{�Ag2&_�[�'�F��.Ws9S��l�G��hԋ�f�b�4�0�J�����4�ah�s
���5�:M������&���z�D����Z12zt���\�Z�9��܆�_����1������ͳhm�A������6��4����(�g0���݁��4E�00����b�RFz5���k�߿o�p�	�W�D��J+^���Rf��۪�	��]����3���V�jW�� ��A�]�5s�׍`uR=�Ѹb20̻�O$ �Wڇ�y�1Nz>�|�p�$��Υ<��z.�~�Q8a�Z��0IUВe�������

��	x�Nl{{'���,]�-C��p@�e�i�6�q(%����փ�`���M�A�sM8x� �ٳ��Q���r�\#���b϶-8���$j�iw�+<���x�!Q�ky4�i�mF�*y���p�����Ř˕��ghfQ�ۏ֯A��}���tv��
��g[�16n��c��xu�v<������a*G"2�ٌN�s#cX��3~G�э@�B�N�J��P���0�;�����g6���͌Y&.0�\�5�F�ڀ�PŢ��l������`CG��zn/�1�F<��M��Ʈ�����Uh&l�p��R��jvlX��p���駖e�t�۹�
�.�3/��{�!W�#N�����6ܦ&6,]����y���FA��<^�R�C}&��={1�Ic_lV����l�5[��b@)]��7���h�Ca�٦!S����R+�g�ú#V���~[�F���Ͱrl@)�����M�ؼ�SQ	F����wc�X�܏l&!�.�Ê��2�}pf3Idyx�v�L��NX�F�|�Ix��g���K�![��	Xc�9����^D�T��|��J/.���*;��V-^�O⓸�a��ې� ��4�.��ls3;q�E@��NOO![����������^xUvoق�N;������d�PE�X;��M*�ۇ��؎m�)��+Uᴻ�d���DC�� 6=�*2�I�bI���>�Q�v�iȤ���/���l5��Q�����ֱdɑ�OG`*�a{Wp@sc��  ���#�z��4� 1
��b������������1�z�ih�]��$E�^)t�:�Wv%Lp����x}�V�wt!2G�.�� �@��	�K�}�X��gP�.��:M�s�m�J�d�BZ�(����v|�+��e�*+Jt�V�#�
��� `�1��=X�n5V,_.9�m�����)����</��&^z�M�?8�/��hRڪ���{Z.d%2��������#�bjL%� ���SRh��J��b�8.����U��!z�#@����6M���"R񔼗�E~;+�6�Q,��͆!U�5Vkը�����y�:�6�5�N
��7�Z�ڴ;�uL��]�dR<Y�)��Q�������V�J,�uvu��O��}b|t���x�����Z�f�UEI�2�Q�4�=߬Ռ&��D$��LuEU�&��>$UU��z��(JU1�r�јI�Ӿj�����Zk�5��X7�u�jm4�ED�(��X�F��o�~M�M�(Ĉu�d��mZY�9l�b6Vmk����d�9���A����=a7���;TG�Z*��$�J['�\x2�#ظ�yd9L�#(20W@#W�R*I�US�y�a�<L��:�-B��o����/i;�Z�K8�T�Zٕ������RŃ��t�'	J���b��$����@}�juqK&kE.�յ�m-'x>x��F���M��(T�.j���L�]��s�]��}x�����wvb�E���Cgg/��61�c������c�~�𓟣k�잜B��\.��e�E�����-�O>�ݽ��Z�z]W�9�����R����K/��?<���OD���l�TpҺu8������/!�/�-Ѝ�ݫ�پ &ig1<����P ���.<����\��$a��5
����1t:V���E�	����b1aA;*���>�:��я�y�t�X��d�l�TBZ��a͢���[�R�؉JM������j���߻���Ka����7a��FFQ��d�����A,q�X���TB^á%p�07T����s�H�N!�I��'���}C.\�%)�42�z<nh���a,Y�\@t*[+�}>N�Y$�	�=r��~��/�o�
D�ii��+t85��%���X�h5�{VCsxQ5U������B�O�Ӊ{gg0W��P��b�o�P����Et2�W7����~�5I(��apd?ڂ�LLO���?��e���������
�h�9��A1������0T���.攼g�^榦�ey�E���߁�_x
�"�v>���T�@{:�lX�'�x"��U� ;�98vP��Ӊ$�y�y�u�.XN$�i��%�6�lW�b}�N�}�Y�����Z��#,r�S-P4�&&�tQ7zB\y�%ؼ}��"���Qs�T�C�^c�ZS�㌓O�� �l�z���J��,�jMX�|9���{�7�F��/�k&���
YTi����`r��7�;q�qG#�aA�b�w��18�ֿ�EӬ��ލQVr,~�M�r%Բ1�<�vQMe��g7cْN�1@0��<*V�lvu�f�1������#N9�,���0��<jբ,H�.�MR���Z&lڲ���fw#���g��A�Xli��C "�w���.�t;�z����y^��f��Ԥ�0v86�;;�/_�rٌ�0]�N��n�MO-fSҴwbb��Al8b-V�X&�_�=e�5*���p���M;�e�.O̡�w�DI��=�d�(��>�'�Ã����HQ�o�����_��N'�<�(Ip9��0|p�X}}=���A�T�N�4<&:��e�N�����(9�5;;�bA4g�@�P(4�n���h�Nb;�5�<Jj���f�J�mXkcvv�Ȫ���0�<�:�ĉh�U�Sn��t��tVk��!
�gff�.���i6!Ɣ��F�Tj&H�)a�ۛ}���Z�f��4�FV<(�oԉ���J�^*kF��f0LV��ȿQ��h4j�L���ɳ\*4M���J$e�Xo6
�mL\�iH�Uq���'���M�T�Y�՛&�������_�y][�N�t0�h��=�3&������fO��ՅL:�1�fmW�2�,��-�`��l>�<E��&J��2le�� Kk�IꔼF#�Z�20R��������fP��HM���_b�:o-q�26��%���t���S&��a�Xh���M�M��{�Aɘ	
gK����JWt�/���:Ʋu&/7(�[T��\vi���]���OCk6����o��0��;�'�JQG�_�흝xk�>|��[1��!�S�p;P�����GXk%LA)����Ux풁h�����z	�Ͼ�2~�ǇX��3r�\f��Y��{�cn�~����X�l1,V':������� I�i�����ٝw��o#�x9vOL�rLͬ�TH�����G0z`��������KVN��S�{�J�=�<��_ۄ�L���qxl������cd�<�g�m�.LOӣ��H�8ܳ2N��#�Z����1��C�뉿��׃�\A�\��B�5k������ϼ�B�x}�pj>��L��Zn���R�=�4{�u��bxbZH�~��n�ǬX�#�.��/��+����=m�܏��6Q�y~t,���݆��wcņ���B>�9p��sO>�r��,�6mK�	��d3"����mX3=�v������;a����Ć�T� =2�sN9�8�x�/�Oo7��/�Y��fa�cø���w~q�����Ȍn��u�NY~j�2����0�*.]�|�*����m�F�X�_y9^��6��1X�^�~"��?ԁ�lao �}.��"�lQI�V)�=��~ϥ3�5߽Nb}���1x}n�#Qs94et��0z`H�k�׸�!$�X�.X�i��.���v�ڎx���3�H��d*��@���\vdg���م�/��RE wGOL�*�8<F@SL�9<��[���Î
��	8vp̠k�M2��Bp)tzC(2a�����g�yF����ǣ��G��L�/v�=��&2(���S�Ș3s?���X�v@��[{��&j�T��#�I�P,W�����ׇT|V��0.M+4w��X�н_��Ͻ"a�Ӄt:���i�Hլ��=��39�4�=�_�,Ւ����02:(����6�]�����`vfZ�� �yFD�#��t�'��ދ��b���bDA��0�P,��`�����۰gp���`��U�����w�IȷD-���z�"L�"��q�mGZ���h�H�v8E0�r�!�}��طo�p]�~O����&�b�%�Nr}�2?�x�81ܼ����ف�^݄��aa�$����ţD��k^	����Ӭ��^Oz����b4�	�#&���'Ȑ�155���zaA8��&�Ê3�#�-�[�������sF`��iu}X픶s]��lYE��X|mk?���Z�F�oa��]Oy?�l�r�\��utt5�^o�\��A-����b~��#���s��a��������Ѣ���x�.��km:W��*030"��7?	X�x�퍘��)d�Ԭ�N�%ch�J0���^��Y�#� �dZ�rTh@�E.��29�g�yo�݈A�S�}��?�w���j$��H�9a����e���7Eyɪ�j6��Y��>o2�E�ȿ�(K0�4�,4*=ߒ���/8��4]I�m�d��\i������_��ͮᬓއ�_��!K�GhC���r��9L0;-2@��}n��vh� b�,l��+�N���_��Obr,.�=2�@2�C�j��@ς~=�X����om�W��m�V.�h|Z�1~�����xǝ(M�`h�nx�>��XM~��mpK�
M�ʱ.j�{~�;���m�:��s|UC>���~s�wQ��C"R��D� ɯ4���/-&��n������{�m�����0�0S��"��o]�b*��;�A9o�֭{18C���i�݃�� ֬�������ˣx��7alk�D&+m�Z"	���;��W���3(�+b�	��������B�X��m�ӡ �n�<��N��އ�dsS�hw۱�Ç��y���p��V �3 ��������
��:��%�;��0В�b�կMQ������K���A%��K����	v�� SH
 �����d�G���{�@�c���+.�ꂷ��럿
/=��ܼ;�"�n�a74�3��XV\����O�57\��͂�Ɉh$+~j�^+�}��/�׷��>�=��tw�C<a.\����O?߽�\��/�`���M#����&V.\�뮹!_�L�SڵL`ӂ����q�8TU<��Sxg�nX6��S�`@��1U�Ҿ~|��	{�����uR{w&�t�]�(���Z����/}Z(��rM���Cc�h�����.��چmon�ş��$C��0��\�M�p�X�Lf���ް9�;�b2��&-u
�*�^7Fw��綺a��Oe��X�d�6�{W�\��~�'��
��04�04i0�@���Ҭ�Y.����۾�#7,��T�	��d��!��*+f�Ia�����=�9�\x]NTK9�LO�uI��y�*�o�F�5�1�x�����$Y0�mu1K6�&���B����!�"����Aݺx��H��������d� N=�D�s���@�W[�� �����q1����އu��`��ŰS,d���6���n�ҕk��o`r.��^z����2�U�Mrcs�,J��H'gQ̥��OMc�E�(�NXq����%8��0>>*�d��~�o���GPF(�o%����H#1'�"�ڵo���|�����ݻ���) �6D|�OL�(݇M��b1d���~�wdL'���t;'���^Q�r�h@�y�s�� �ń.x�:����y�F�%ݛBA���U���Z��sz�$������^;��-�@Ҥ����YsW�>3L]��Vk�bն�x�I���,�m0��=x�g �w[G����G~ݴ��O�2��F<����ð�ˈ槰gri�y��p�ٌ�5�T�������t����.�V��1b!����h]8�^��E(��I����U���	�*�aR�ʠ���#���O{���� �m�V�?���l&鞬�@Uƪ"�:��ס�a6J��=�F9�ۆ��x}l�Dd5��A����RP1����=����X �3�fF"U�jQ�6.EE5W@��D.OՔM�Fl�ɪ�d�L��C�x���^�3����N4�b�����179���4�*�P6��n�>�K�ϼ�
������hT@]�m��_���9�
r�Rɢ(1��Y?�ǎޞ�ܜ�t
/oފ�،�j� �\2�JvK	���]=.�Y�+&LL�1:�ƾ}����>��6;�.#���p�-�1��ލ}SS��Q���_1�_܎r*�h2!-����L���ݭ"���Z��_���ضoe��3����'g��=w���`vb�T�����)m^�Ƙ��݅�ـ��	����ʛ[PWU$�9}N;z~��/Ǟ77�ި���C���*�h1�\%/� ��C�<�{��(Fqt/_���R�[��f����|��w7��z�Ξ���+q;����*��;��|_�Q<�⳸��ua�����9���]��<�|<pǽh4M�=x s�T�"�(ڼ~�"q������]���)<����{j
���b,\�
0�ŇN?���7�u���de�Aa�ö7���������(���R�-U+�eG�V�N?�\����76art���1�<~x!�(>���	��/^���6|��_���¾X��]*����O�����P�\���P¡3,v\63����d:��doL�c�R�D��9z�զ![)"�s���A-���m��J�l��k֬����ݍ���;l޲Ꭵ�7���N���^i�Z̡��yEA_O�z��jE?,f��e��K�R��P�R���}�(���~����BD��W@�La@;�h��1�e��u�Nlڼ�]0**���c8'��WOf��L�-��&��*q.�o;fH���d�b\t�G�j�2�R�Ѣ�4���
A��Y1��{p�1Ga��X5�Z�
�&�n�,���oB*[ų/n�T
f�����9lva��i
Y�RL�\.Hh������JHVwI#��sq�m ��~,D!���p��b+�yFDe�@�������Slp��P���'���b��(�"�R���Ֆ{��m�&`j�5)���id1���糲Պ����.�V����@|A?������yO8X�/�$���E�C>����V���XE���hJ~&�F��G����Ԉ�^�l#�fv��jR՝�w�W�����mޛ�{�6������j�<�����,���m��c�?5���)���j�t*/��z�~��V
�'X��wK���[���Oš��yPt8\��-�恗�j���9h:�(ת�&�B4�y��
��V.��F]T�U.e��;ɜ;���ml�1ԍ��I��1�A��WD�W�Nn�RQ�XI��n���le%�4��TQ�.���YDShU���~��;To�<�ͬH��r�,��Tff��y:B��-�5�Hr��fU3�C#�4b�Y�6�.�%�xFQJ.��Jе    IDATZ������dr�a+%엪4�j@zbn[*�U��2��&O���"jMp��ךh����ؔ8�+���:��h�
(�rPV�{�T/�EF�7���
T��tb
�U�Ն=�2�u�<��amo�1P�]J���R�!�#��@��B��"�kl�R�ˏ�XRV�����֭��&��h,��AE�ebZ+!򣣫S�_ټ	�����y0�����p�/܆?�df�ao�P*T��1�PU�/��ݮ�e���I��G�gbM��LJ�!�p��]��-ߺ���S؝LN�adt�R={q�1GC�Ꜯ�|�{�a����
��:̌�QKX�݉k��3C�0�V�Q�MN�
�+܎s?�A���pZ,����_�OLe�((N$s%8�6!g�t��������m���N�.�e�;�$#� m����3_�w��n�o���(�Ę�{߸���a���H%38p`O>�j��N�ڧ>y	�����q����bV1M ��6>����K�~Q?^~�1,^� ��3���A!]���gޢ�d�îapt�fg��ix���$f;�f &@ٿ�2�4�m6!h��ؕk�s����>��6��`����`㫻�G�B04 �=���Y�ý�inLMLˢ�@��raْ|���`ْnh���i*�]����М�H�2��{�����>�f�"�	��S�4�ۊ��rt�O�J���߉���F�X����[�-%��x��c��9Kd�(�LV��4;�SY�K,Z4���
��fT�eIB��F�ƱYr[[�l���W_}g�q�K�UBF��9<Z<X�z=�{i�fSغc?̚�SQ��*Uia�i��f�.a��y�-�ɺ�O+���rH%� �ݑ6�F�f[v� lŲ凪F<>$R5���|u��$V�v���6�n�*`��� ��cJA+g�W[���#��Z~�Oڅ�<&`"�XEaL�Ŀe�`�!�V���[�|=?�e�K����VRLyy��l�� �;����-m0Hu��Q��>��lM��#��~�3�^V�@e����9�Y�{�q��z0~���J�=������x讦�s}��^sF����lqg���ѽ��
���B>�B6�hA1���	i5��T^-'D٢Pc��[?������ٍ����­>����d�VU��@=p��(ݒB�^z&�>�-���:�#�b�ɬ8��, ��S�����tT��萹�\�ͻ�Pd�w06��88YŦ"���N�Ь� _Y�N���J����LA���H���HR��݈ժ��4��5'ʕ<f�s�8��6�~d��X4�*�u��Hw8�B�-J�0�j�#�l����:�9��+�9xl6�2qx��Є�bU8t௕3"u�wU�^C&��1	�ND���� ��*
���E���/+F?1��JV��&�E_[���p�f�i���BV���YȠ\���a�8�-"[����OT�ss�@�C�����8]�d�kV<�N7|f�=d�b������`&`�s��D���f1bvjn�
B}��.�0���f^�j��\|>�*L���Vm(P�=6�]�v�Y3#�/�Rg�x�ͺL�BʵZd�eLu-��ɞʴ@�G�R�|Z�{_ �d,	O[�B��>TU��+c֬K�46;:�N�
$2���]�R��c���y�|�"d�N���� �/ �ʢ��`���#C8i��(er�����2�/	��2���������d�}�����8[��QC��F�*���;	�xo��Y D�j�_7U�~�1�;���lzi�4�Þ�k�U�f�2|��VҚ�4V*�D0ԎSO>Y��G�bbj?��p���&`�h�@�L������*�ڼ۷nE�G��P� O�U5�\��$76=�s�(x��6:��fC�Zժ���B@Sa�'�n`��<��h��
��B8�>���;h[�ZÎ\�Q�Q���,B�-���IXM&�Z� W]�1�[�����T�:&!��5���bG:��7��-���G�ū���>%����y6�I�(˰9�������ƛ~(�/��+�C:��牀��YN�<_[��,Ǉ/��gt|&�����E��W��7��/�� �gj���Z(���w�q��atvzq���b�>��p{\B�z�:�JŀO� ^ym6m}�����oG$�G$��jۑa~�M�1��4ʥ�XyHA����v���r8��81;;%^�|p���+�j��C��_�I#�C�gEj.[p�{���H���XB��R�CI�'�=��)�I��L&5|A՘3�-�9�1#CÇ���-�X�-	 YijEM�M0���'_�"�����(��Tӳ�������(�;[���;~���"(㢄`SVL)��u�/�#��u�
�;�09��iRL�ׯ?���C潩��-���	�n��w�������*�����:�p:��
hԒ(g�ⷣ6�[>W�����4��ר��V#%��?I�?��*]����'��?߻n)��А�z*9GT���f�F��mW|����gT5�PhԑCCZ�TB.N?9��u�O�-��Br�PI�g�
+e�MȅɕC*��k�TK�*f�5��ج�bQ8�f	��:�����x����Fdj�ha��y� �V ��4�����)~ a�p`pbma�<�PA�[�ٌVɄc[�QI>�G&Lz����$󏼞"e�F�ҖD#_r�h�jU!�3���p���XD���������Ѵ��'��ٞ��a��rx�\A��(�p�5�.������xdp������(M�����/8���֔����@��[
�y��tJȽ�JY=��U���.'l���t �se�EH��	�������� ��ܺZ�j]��R�E��/�о}B�R�����p�F����v��	K3���}��M�Uq��`���'�6K�`�"�rV2����1)Go&&K "�`u�F��b	
��D�8.�M%�E�:3��cg*�	�fi�y�Uԋx�&��������
vee�Qhq`D���Ea�	�79��+(W�	e*�v�6�UxdҢPu��SC��h]���L1;yc0 �ʄ��C�)�$+�O�J�>�`���C��[���Ǌ C�"rc|fMՀR��t��l�$����Oxc�J�r��8x`/�߇������@"���{�t`�K��~�� iV��ƗakcT����މE�~�,��C)ců�|��a�\X�f5��y [�@[h�����nڬ`�i�8=05UQ�QC(��w��E�p�:�ky�v�#	��S�d��j��i�*"�\Í��,H&b����cnv&�|�d�����[a�8�\�����O���>��"�c\��D�!و��Klё��q�-���K��_���Zؾ����u�@Ӧ�!��/Ɔ#����|�R���xٚc�E�Oy=g�Uy��xi�رk[���\4Us	���c|�+y���t�09:�Z5��"U{����?���b�
�^�[��Dt�����P� (
	��?v	fgY)$Q��I�EI��qBO|�[�����{9��ļ��Q��J����A~f����8ɘc4��Z1S���a���'?��	kq�Z-�Ýd>=,��uZƽl���ժ��:Z��_�&S	���}�}lUЄ�'���Y]��t��v�}ς�K�b�Z��_	���4����[�z�w��a�[�����(�h��PN��i �7,F�^��g��j=*J�h��[t�:����ɉ<��OY�[̇�][���ۘD�<��R�K�4]mɥ���`��/!���̠H�]�U1�e����1���ި�ź���]���d\��b��qN0�	�$%�@ �X\J�JU"S�*�OGs�	�I�+ex�NL����*�*T��s�X�a����K1���0kȣ�B� A��ME� ("�����,���"�bA&���a�y=����� +�C5 �H�Y.�i���/JLN�h�d9d?�
B媌�:���f�c!�9rN���������g�J4J;�i��$�JE@��5�r4��"RmUo0s�%�g%�FU�Q'wt�K����V��`�v�L;��\EӤ�P�i.�̬�1��>KM�:���<IX@?�&:���(2~�50E�N��D��F���l� ֽ�j��^}2�B�yr�^��.�(V��S�Ҁ'��j����B�lF����U�U5M*jeV58ț�b��$f��=^9�'�`�9���,��X���{�(;��JtW�U�n��s�э@$� �$R")�
$�d[z�9'�����~3��z3�Ҳ�h�T6M��42m���T�HR#@��@#4:w��s��}���mj��֚g�P�E�}Cݪ�η�9�썼O].����ZmD8��*k�_G��E�"Qէ
�+F�CF�)�q[6��j]
�L�x��FD<Ez�IC@b�����w l�_Z�C�I�Fӊ��x�m�kI~[���ґ#��/�d�ޟ�	�ဉ�@�̪b	ղ�|V�m�)8fW�ۅ�ʢ��O Z�K��|��s�琌��x���NO��qL,��ɦ�C��<��E��p��ݸd�i;��Ϟ���
2�>��ana�x�;HgG�89�w���>*��l�L���,�uE�O�,�w������hV^��b1R7�K�.�IH+�>�q:t��6��?��p��	�q��Ɍ�v,�F�E��n�w��8��կ���z'JS�·��tb����'����]�`��1�אI�M��\�[o�E��x화p�ׁ�IO����ǕW^��C�8"��1���%3�M\��J<��O09�ǃ��!񞥴���| ��"��bx�3��V�y�$f2�L��x<�s=J�B��@VI�̴���D��TO�~�; �9t�Z��#�#��6�Mo�EZw|A�{4��5%ӕG��(b����^�۝�ץۺa�5?s=[?_��������S��䗂?y���\\�����'�sDPK\��t�����!����=���ݶ��P�W�������>tǽ_��F��k�~Z��.V��� ��]d��0�G�e����M��N�XVܔ,h�ؚ-A��;JB4�X��#��T�?O�U`?^�:#�!�Y4U��:]T�g�^&3����  �:�ʶ�&N�����4�mX=Y��/I&K����nS	���?��p:�)6�-7�v$}$*�.��>���₌�W)�hX*q��r�XLDX�Y��9!�jh��1��yů�f�Qw\�,�?:��Aq
p|����i�du(n�8r�J�K�Kf�!�n�,��Rï�0��Ь�|"5P�s��Mc~i^Z�I�C��@��G޹�[0�m���O�ԫ�>�
�`�<:}�2P�հR*"�d��E�r7*\���&13?'�45�FCM�pf�t��Y�'%&��obi%�����dˈv4��#�*�C�X�1p�@N�ҽ@�˱vE奀Qh�&]7�k�U
Q����$��Qo�I@����<�\`���D�s(ϖ.̈)�
h()r^D �ڮ��j�ZWU6�'�Y�c�@f1��U��E����j��s"Ry�Ģ0\K�t�xZ�"3��*41�8����-��,W�arB@�D)�͟W��rE�	��B�Rpˉ[�DV���@Nm�|?A-uM�Z�k���t亱rN�>��몷c�����&�}����ٙF���{3pQ������	�Ù��pZ�
R	�K�b�M���T���
��TԹa�>4]ӕ"�t^6+V:�Fej��G��݈�ҌLY>t���j�%�8}Cè�|�z7�R~��SXZ.H��r,Ij���6l��&$n������Fo6����(ҷZ�7p�ЋY"�Z�лՓU�'�'Ҧ�x����'�t�9��rj��+�2	᭼�\F�����5|������y�YiO���?އ�q�� �Ds�X�`2D
��ܴ(���[���9��*;z`J*2����ż ��ø�˰RXƞ�w	 $��/EQ	�H�#�5����S��ґ�xv�a,�KH�{�_.��V�/�Y����N��Plh�'6w�"�֢�E����)B�
��?�x0�;�oX�WU#z��$	��9���m��E�[�l�iR�"JW�cPU������y�I���Y��.�Q�1�ʗF�
�������+e��V�`���3���y͸���|�Z�D�)���^���d���%($�@�A�\9/�f� ��a�_����'��_��;���Xz�b���H�P,̡'kb|�Bܚ�U;cx��!��C�XFy�&���B8oJ��/�.e���c�ր��hzi��/����	��F���u��b��f툉�ǖ�2�%�j!��j�y�Y<v�|��MC�ؒ�3ӧ���S*�1�-�Z���B{Ʒ��k�Ŏ�[�Ph�DcӉ ;؃CgN�C/���CܸA��TZx�^�������gظaT6���?	)��o=�-�q4Ѳ=t�.�4F7���?�z��r��do��"�H}�L<���3���>_ī/�S��k�)��z�0�����Ml�|�k5�;uT�6�Te���iF`�L�_�/�(�ԛ�\����dЪ+�@�bL�#�(n��xF�7�����c[��ɠ ji �\!�%*��s��\s<���6�?G%�-����{Q셣�q�� �t:�J����i�!��Y��\j���rXy_��	mi;�V5����H�t�MX�I���K���f]@���X.�l�� �u�ֽ���Y��z�?< �|�:�������@�NM��	7�Lׂ����i��J3���:�� \�'n]��ևGN+�l���'�%>\߆��/�@i� U&��=�vh�E.��+z$"�~n���$׏߻T�J5��l�1�9�)Y~ �ɿS�X���Wc���0Z��5�B�J,�V���`�r#�W+�V�b쾰��64"^^���8��f��LD��M0�N$Q-�Ѣ�!5#������A,��ߨ�+��]\>2�kv]���i\��l݁��!�׏�>�(.�d6m�.�Hr�>����Vz�8j�&f�q������mv�zߗ�JD�ϓ7���Bi�]�HTt��j�������A��NNH�`%� ��rr(g�*�+C3^���:1��'@��&�lقk��V�9��,�������t�r�jk�jr^���J���oŖ�MR-a�����+��,�V�8�^S��O~�3��w��.�&�p��;��#f�QkvQ��x�g�q��94Z�=�����/� ��QT
�رe�zI�#+N���`��Q��#A�M4��wA���J���'-ٖ���ѫ��#B��" �b9�����'{TTU����ꀄe ��ii]����z`v`|�
��i�����W.�k��0��1�=��y����31�{<����$�g^��P�Uڥ��p���i��aF��B�G������#�쎯|�N�^V��p�Ģ�Y��������wrVt��X$��5�p����jԪ/�^��S���lDx����~\�\�*��6�GBQX%C��^�}3�m��'U�QX2�,x��?5����	�g�0GAZ*�Seɨ�j�p��1Q���	�,����2�����)~sS���O~�TOc�8v�4�9��gOcx|�S�hj��W�}�z��}Z���ʙ�s����zS�� �ʎÌy����q��Qky�1�(Vh�n"�b����־aL�������ב_Z�K�ݰ�Eo��^���8I��P����>�es�5L4uN�v�����Ͷ�G�yaN��y~ԍ'�&�%���*2�h�REla�6|�6�����Z�M3��˸����gP��e% 2�1V#ӵ�l"�ސv�C��4j�p���H+1��cn9�Vց8���BkU��L}t�����6I�\��D�䜰r��$U �	�`]+��>ߗ�b����,+    IDAT[AI�W�], ��R�2j�����El�C1���sP%��)19��z�Z�!t��k��Rԑ ���Z+i��<6�RGu*%)�@�Q:Af�-|��y�{d��-�@��l Ae/`|��/����a"������ے�g�XJ���z��E��K'�P\A�\
Z�Tr	���pW����Z�R��6����J>7\ݶ���ڳ�a&$�6'&0�p�E;��G1:�����+�v^|1��6�?���MX�06�I���T�������?��H'�1;5���>����p��l�g��O�ѱ!�;U��Y6
yU����WKےհx"���,�+��Q�nD�g���1��h��RיN?}�g����S�Oc���ry��J0��(�r��5��w��W���kC�"^��t{��ӛ�<擒������9/<$Ur�{<�{{���?$C�<w@Z�����rF?-����T SC�ݨk ��Kq��!4���l!��+����^l���	�=��٪lR ��� ���
�`1f��ʎ�,�-7�ғ�R	
*S��&�.���nG�����iФ����{�a��~�z F��A���i�&�RN�v�~̪�~��UV;AeQ�j���Ϛ�}�a���(H}�+֎$����Ȏ�4LDZ-��@�:���6Ɔ;p�3�����`����S�kb�J�8G^� ,\���0�E�.�/�j�+$�*z_�h+˿��H�^��J���mײe�IqJ+0��um��c�k�K�'~�g�O�O�D�� L�A�â��ioD ��]l�-���[ކ�R�jS��sg�"�����iL�q��ǹ�E�s)�&{p��p��d�It�m4;���'��~U���".[�I��6l߈�p˵%�/j���S��5\�����Gp��f8�&�x���d��vb�MO!�/�I��sR�x��1�����M��Q%p���>��2�Npnjͅ�Ԅ�Ҁ_oK�GԦ	��ob�l9��-SAݶ���	R�n�\c��+��ӏ�������w�M��M�) �6�^;�\W�ۜVm��#A�b�Z ��B~��>���*"�_ge�a)6���IJ`80���<��Q�+
�T�*�*ۢO %�d���l=q8E�虵��C���3$�
��0K.��0_�6ڰ�轕�F۵С�AD7u�"��&X9㄃A�$^�`5;���*���mN�s����[��3"mN��XU��gU�g�B L��!��k��������E�̫|�d� �5�*�T �d&8W��Ȼ��7�+��	�`#�ː�D�[�k+�4�.O[���#����-�9�����B����jŐ]؈8��a�L�Qn�m�\#1��Yx�x?b�,6��q}tOhw��T�U`�P,����E��V�J同�b��<��ܽ@7�N����[�ۿ��q�e���=�Pŋ/��?|L@ضc(�PX�����|�>��o����P��G:��0;b���l{lp�"�ĨҒX�E2�Ȫ<[�������7�R,�95c�Cy���z�}�v\q�صk�PT[������҃�`�'g�kK�L�TF��?�/�?z�)g1�i��vVXb�4��.b�2��:;�7��0-���13��ޞ!I�L���\W�ݍ�gN�c*m/N-J��SrZ�B�*�3�}��(�'���"�+>�B]����G�כ^w�|F:�Z%��LM�'S�Eо�n=Jbh�I|
8��A����w��F��qkB�/��Z{l=�{j�ǿk��S�z�N��z��`(�U��5�� �L�k�m��g�P㙯��+¾���+>r��>��l��J�l�'�A�>��t	�7u1�i�������t������w�(Ljm�X^[$q�?�ףp}�UFppX�W�iE|��RD3a�٪��:h٤Zu��@�A��`EP�d�?���8�f*���P�3�.����c)iBSH�
��H4L\2�;����;hkHEc�W꨷��t��w���JfV2&�P2�;��ؘ�o�ӧ&�s�b8~���ǱP)��b2�H2�'��#H�fPh-��K4Θ�u�&̎���N>��F� Y��w|��JG7�j�\@������/,`���%��tL�����0h��u�k!��^�����kđ�\�ȡ�;U(�V�t7:�t]jVs��4���QQ8��d�b�5��-��+��䉙t\+L�C`�ydƮ����?}:e�HPb��15 ���g<fV(^+�F[�IO�������H��{���	�KJsuU��!�&�#��G�������è5$�H)�2()	��!y:Ғ`;Vއ���2r%	0��q&?�2AX� ��{�Rzs�|��ڎ϶�k�mg˹Ձ��@W@[tі	�҆Ul�k[0���B*��1����9R�40�5�c{Tt�h`��S��>���ҲU�M��.�W5L"\PVjİBm~jc�yQ�Q����D���u��$d��^oz�dc	B�%�W�S�4���h���Lǵ��[^�$̱ܩ�f�f�1���,5W��1�M`��`{"�]c���'1�q+�GFQ�T102,�m���x,'�K�)�d�)�͉���E|�λQ��H'������=;1:6��><����JNd_6�
����q�W���߄驳HR�,�b~aJ*}���\��i��X�k�|T��S99O��Ze+�ׇ���ɓb��*��\�$es2�v:�pC^%���*�X���t,V'�X ?��Tet8u�<���/cjjF�^:���v��I������˯�W^���q����(k�\R<J� 9�a�/#ڄ�	��'G	�C�Dx�;U4 i?�W�=�: ��<h	��4c&�#�G�m����Fyo�3^�U�� +պ�0�U��	�&��1 3��0���3~��Tk '�ڗA�-��@l=�
�N�6F��	�Z�sm�Wq[���/�FQZ#�w�Yی�c���a�����+���wR�.�5,8aq�U9�L<���"�9Żo���s�1�H�Z���ͬ�^��2��r���E��S�Ot	2��+�G�������"��O7خF{�JwF/V�H���ږR�oY��u��M����(�{�	��0�j,�*���A��w8��(��Of�vd��h�;�FP��ǀ�?;�����^Aͨ#9܃�y	f6��i�����M`$�B"��S'N��R���iU1p�^X@�ZG�M��e���0�k��)�k0�&��6��q+���Y�~�E�ݸ���/��\v9���z��
�:NNN���s��d�Lǐo�`x6��P(�c@�⃱(�Ti�,/א�F�i��vY��['�M\G�d)�J��^NE��#�\�l�VC�.l�C�݁A^J�%Y�O� ���E��rn�܈�)&]Bg�����a剭�B3p����V��mEԆ�b���(�'^�%k���j)���ilK�F�:(��ARG�i��&��vb(qb(���>���*�����Qi����ϊ��B��(���~xT�-`%���Ҭ��tqzv
�nC,�Fb�C���Ꞷ)]N�%<�>lue�Zl��@�T����X�&b�*5ݺ2��|+VH��X��ԛr�b�T^�'�&����J�$��*�iV�r�Q�UQ��d��*�:�K�3���*e`l͂��Է����̜����H�T�p�Z�GH?$@sh��B�r�l�$�zk�ZpMQ���̘����Ly񴅸�F��1b;x�uo���+ߎD*'�+�Hr�	Q�cY!�g3=��>/f��6���J�c����_B��E�7������st13?ǋ�Ҩ��:�LcqaJl��9����M������#�ɒ�MP�	J7W$.�)*�ј��X4!�Z�f��ϰ�zt+����X)k�@���hN>[���(�򹬈r��1�nK�I@V��Z�a>�P�$�#���u�ؾ�E�R���Ż����	\{�x�����{�C���zS��E�[$&ٞc`�@M��b��SH}.�8���w)�����*ykkDvE�WR6����yn�/(S�J���b6��@U��[o{s�<�P誖Aʸ[�'y�9U�s������ LW�t�"��N��V�Zh��w���;W��5��g�=������$��Z�a*��I�
1L_Ρk�c�Ν�a�{���+��}�������G.ow�8Z�)�\:���6�m�`SO���oFm��r"�ӆ�FQgFJ�ۘ�F�.�$Y��Y2ce�&!4�]
�BK@6�i��}�ѼZ`��yI��1�4G��Ѣ1`�J3g���N
�ꏟ��zը�z�a4��X��P�E��ْb�հ=#��],bk����۱85�N�)���(�s�~ّ>w��>�/q\���jSn I�EO.+��r	�~�;8s�,�XB��K$�'�������َ�hE��r��B�*���r&:KUL<s;�FQ>3��o{~��_Gai�l�s3`���?���p�=������8={]�TP +�ɀA.׃\,�Ak���\Y��ϑL�u%�K�%����n;]%���Qo!�ʉ�%T�J�U@�9�P�+S}lq��-����r�6����0��Njs8��.������=I�>; �jT`��Z���[Q$'hip�\�
((�揪����C8P<���eyd���j��*�$�ӕ�j��f�Μ��c21�xD��m�&osnⴜ�2!��5[B�O���H��]�Q��X�!Z�$d`�L��$�Z9GM.���>?;'4�7��� �3��I�LJ�R����kIYI�دV��L��:�El�]]?��i�</Ș4��H�v>����
���*���ͪ7��I )�͖��
tt\�V�е���FS��lC�IJ%�o`�JC@:�^�b��cR��/sʐ�5�D1�X���~:tG�@o?r�^93��pbQ,��Qi��a|HD��eN&�D���{;��k���Ԅxq�"����P�K�S@ 'ߊ�J�������¢�&rC�@"%���+��QO
H!F1�چ�ROW@�*<yi�H���uq�r��ۆ�1=qw���9=���Qi/�-,���;��KW}���8u�vIYpU\����L�Z0:u����8��S"n��\�!@I��$�25�����Vabkޗ���:���&�9Z�tp`XX�ۼev��&@,�!�R1��x)�F��Ɂ!NY�'��F��	���0�-�o�<�Z|A�C�NW�t��{0��Е2�N�N�����C�Ĉ�	��R+�!z�|�����5��5�g̛��v�/f%���^�_��ϵ���kM1�� 6o �2-��_~�K���\tV��B�O�C��Oښl�)���w�ۑ>��u�M��`��*��	o*)iR{����R-)_��7	�Rʥ��`���<�T�I��d�3L4�f�5<v�E���Q��y����l!��Y�V�FjSd��@l��Fs6���pn}�kq��q�y�!�Y����0_^F���=#��e���p2����(.-�%K��s���ѓx���Pl�P�(�M�qWT����"9��r�#�a���ɭV�!����K8��1l�c�I�ݷ��x��p��I��n�J��|����&���G`%��q��-���H�X���'C�M�]i!�v�\��-���D����3;�s�j5v���D�E���f.���4���d!BM��R�ΠF�ZQW�ށjA	�����-r�9d���֎�Q�*�+�v�Q��&KH�4[_�WO�[���$"X/�8����������-MYڱM�dT#'�2��n��"ZU��i�E��luYyyn� U��m���l��C�M�U��o�UT�#�&�RG�	D��|�H�M�i�Ͽ�n��Rb$E�D��rMΥߡn5�q�4gO6� �{�ɚ�®�0}�x��qe���������Y
,ȵ�8 � k��ڰ��M�9~f��p`���Ӆ�vql���PO�������M�Plv�؈�ͻ�ƒ24�%H��E�d/���P�V00؃V�����U�&�zǏ��J�(mi/��Ra	n*3F�,�|�b��]h�J8z��.Л�p�MW��8+�]E�D~a^�n��Ғg�,�0f;��/x��*�����d��Z�-�0�B����*���*�H��׃�``��S������覍�|	_����Y��v�B��B�2>���"'w�Ң���+$�M$�)(L��ģ���?����s���O~(@� �֠�RY�h<7�c��`
��s����Aα��A>��cǎatt��7��^��kQ,����Z��ga�2�$x��F1b��TEL�0!>\W��W�I�Z����5�0�X8~��KM��a}:.3��*����$�F��6��-���U¾����|�������kvl$��|�P-��� 0>�ŶA��~���;�^'��(mӔ�{�Y|�{��N�� �ܶ��eA���ߋ����� 3��2o� ,A<����m��/�^�Z���B�g����հ`!=���
�:r�f���Pg����HUo�<��AuD�İ(ӅKF����c��p��=0[\�>ʭ�o����#����=�/��i�.���Zq4�E���7#??'��?8��^�#�~K�"��@Y툻H�eK'0�mn���jf�C�ے� ��Jb��<��P,��o����|�0[*Q�^��񩻾�G���1ԭ.2�YDc��H�],7KB��X���uKڑ��*��#�d��.e;���x|+��"%`I�^����^V��3�_�0GȺB �ꈪn�:R���>	�z\Zs��`a-�
@ͺ�\�W�
��0j�I�MG�d)h�AҚ��,gy�����X8����j�I�j��
��(��LL͜�<�`�D�I���qӴ]J��qt��ك��	��%<��sj�^L6͖i�深���%pzMչ%Dچ�hк:T�h���V��7��X`���Uૅ@�*��+��NU+��0wD��5�vT�W�@o�:>�E�VUS�)�s��@oJ�N}O�j�D�6XpHn	�:�|^�$w��S��K�H
���m���9���G"݇��;����T��LE���Z3s+ro��m���i�A"5������Ph���3��6]d29ikF.�Q�F�C=��˰8;�C/���C�����^��A������݋�������T�X�f;�\1���Fm�F���#��B���k'D�%��D"(����(R%� '�4�)�T�:AK���r����������ܬ豝;?�r��E}��q$�ēYL���*+�MQ��Q0[o�@� ���b5��;����⮅���G���8/@�q$�/~�LX�桍�uB����`J�K��;�5�,����'b��Rl�2�M�8uꄴg��!	���]�L�*�E��*1T����/Zuz�(�a��wpi��r0u��I����[s���(�x?�{�JD-�p�3�����<���P�`�2�{M���a�x �·~v������"ٽ��%zB��@�2���&F��x�����7�p���Q��0�(��"������
:4����A/4yA��KK��-�+�W<3P�a2�)0��(t/2A=M+�kI fu%�RSjl:O��(�K�\~��(������c�
��d�M]�)�U]��T��ڛ�m�Fٰ�y��@2�C����ch�R���#(/�׾��E���_A!�kNF�o���������P.�������=$�2H�f�q�FI3�yd��i�V�<s'���װ��&�0�1O��W�W�܉�Ǥ�À�c��?>��>�|7��P?��m`�)�+"�l��I����'1�GΏ��PD�񂍊�Q�xT�.'���P��@􋣈�˴�7�N�+G��Ցpucvڪ䭕�}��%�TS������H��ɲ�V�A�bt�[[k7�
n'i�    IDAT�ɼ@���L�<c%,6�;�$��	�0�6X�4[mG�+&O�X�6eMV��� �c�j(��ݗ�֛nB*{�k��F���ߏ����r�V��ǥUtbr-����Z�YFܰ�W���p� ��Ť�A�@O�����(��,���<�6��kch�[ORj��>��L] o��@M�o4ј�-gG�2[��u�s��k+��*�l��NPh��F>c�R>��&����h;]�g�	ǯ!i�xӫ���@/^8t�A*5������⑚��E,�A�H>��H��N�O�0�V�����pLG��l��k���\�п���]�뮻3���]w`����b���3���r�_؏={v�-oy�x�*Ζ�V�*�	;T�'���V��U��_UH��G�ir�(����x]Xq�-<V�hU��|@̺99ȵ822"zd\\��5�n	�r��D2���`%��d~��x,-y]�`3E߲]�Ky}�a��05=�{��?��UG�B�"�N�f[j�Q���:��� )ҽN���\Ǔ���7�N|{z���+�*����FM�'V�U�K�0*�ў>ˁ @��^�z�K�,h��c��׃ǟ����F�W\/��h@�?_�3��iR�+͋��$� ��p��_���0-3r�iڟ���}��^�?<�׭�Х�bf���C2�26orЛXƎ��WnF��qdIF������L�#��^,TQ�=P�!�ޘ�X-]� �����-b�bm����]�¾ 32C�Pm���A-"NQQI�^���噪��`�%D�+��.'��+E"��ǉ���x�/rZ��N�0S���u���g�Tf�[��޻��&��4/�h���o>����
�΢Ш�޾�۱kd���cj�,"�+FT���g����<'�b|�1$�3�璢�x�0�c�'�_~;��N?%���#g�|bR�3������l���y�, �I��𩿹O>�� ���m݈�@
��'w��n�*B��zͺ��/��pj�nv�G e1��m~ s�l�I�$���L[�"�#����r͆�li���!��E�?�y���)5i*v+Xk�D�lNo����S5��4��ƫC��0����ᠣr�O?���t!�[e�h b��͎�9 �ӑ���u���4c"�J����-���1zY���I�q��q��ΞG�� |�[x������Mb�]��\��:��^;.�|U6#�xh�ōJ�D�Q�>gP����¬���`]k���[��ҩ2q>_on��u��#�A�^s��9cՁ��c#a��_��jAN�����ޘܑ�ɇ(�L���0�;�v��d~
��0�U��p��K�}|�wn���fg��,4�L� ��yzY�J���^$�e˽�$��ơqL�����GP(����I�n�tE��i�\/c�U����Ȁ���xm9�/bc�`~�.�;i�Q=��_4o����b��u��J�$�M�聾^9wuZ��G�#��xBp���y�����u�ʿn29�Պ����Q�����K��ĉرc��(�_�0L�SQ݃O�쎅L�_\N�>-#�3`lqݘ�5)OF��ߤC����߇�z&'��������̴j��ղ�N*��ou_��_8iZ��\��j���i�]c[5���k�~R.�s�v��w)��4�ł�މ���?d���h���9֜��P���=�Z}o��AR8���kF$g5�j�?��ߩʠ�h�X��=��t��9}>�݂�1�m�}�4��8k����<�����X;��>y�������mؾ�X�è��Y-t�s�:Eþ�~��7�x�0r,a�2EΏe��<���ĩ���J�bYZ$�4Z�ie�Y���J��-H~+A�Wʤ���m���Đ8�J�BЈ������F�}k�fbPbLB������b��2t�m�1<�8`�RJ�~[6
�P[i��8Z�~������0��%Y���#���v?}�1t�"���h鸵6~����W��VL����xf������{�ԧ�T-��V^�E$E���c'̈�JX�.ڳK�X�ϞG�O����M�b8��[o�Wlنv�����{��񩿹/>�n,��M#ذcќ�j��l����>��ګ�|������߃�M`Cfv͂_l"iFE��c��m�! ��Q�w���p+�2�!]	ܙ�ʍ�j�oDnҺ$..|)�Sm[��A9�ן�e"�|>.�A��U�&�+����Ѭ�CmE´B�5��
5Y* a���]GJ]��na�nu`�W՟�a��֑�;��r	G��v=83�4���n}����4�C8�.�Vq|�$��:~��qzn��^��	�(�Q:7�,\i�i�+�Z�'�}K6A����$"��?��������w������3��� �����z�)�hhJM��x<<>'7F]�����uxAE6�_�AO1b���gk�����&�B0{f���
�햛���*홳�[D�\����GǱ�ҫ08��Tۻ�TJHg�P�Jx���3_��P-7��j��eQI8Yi���1�u\�w/�x ��q��T�ї^¶�c(�,��+�[ȁJ�r�\��R�`Q&A��)��*'�k5i��1>�LBR~���h���Ǥ�M�_N["�kU$D(JlZ�:��"�ʪ�p��\.'�8t�b���Y^�l.����u�'�O~i�V���1��
STڐ�o�-	jܨ�:m�ȭ�pM<��71��� ���~3s��FȎ�{��*�����0����EJ5^�	y�^")�K)�w12<����}B�+��ĶG�5��q�E}�h-1݆���w(���� �J 5E'\�^�� 3�dtB+�5d ������
����.��\�<Jz�����0�D��S�� ,�i��j՗J�k�P��æ)wW�������G��V�z]ׅ���ǿt&}�gdB�7�i��Ҧ���I�Ȅ�gMRj���d_����|(M@im�7	..~��2���%�FL^�L�b�_OMV��䉨��m#���Y.�5Z�@T��J"���p&��U֬*�Vz
�"�J��y�Q����#h:���M���:�s��0?=% ��j1��SO=�O~�3X��ъ�J[,�!7ԇ�z	��킝t��-��Ql�P��L����I;r��)&����܆=���E�X(�Rm⁇�O�yV*���/���A�-Mcd(�7��
d�&6cf�����=X.���-����ʦDoQ���Q�$E:��D�f�kf;
Y�V�=I���a��Wi��q�4�Z)N���U�@N��NI��-�6�hEi	-5-�2��^UT���j�*�%�Bb>'p��W������"m�sBO�[��������0��}�EeՑ���ʤ�m�	��i`|`P�#n�CCC��� J����"2�,N�?���`�{�"�#!���Y��0mۢ+��<nݎ���\����Q�p�_?	�!	���ZѢY n�`WO���i�9����c�V��I<U%0$��w<.��3�pPD�V�������F ��-�WUp�0�0A���Ȕb�V@�T�;o����ɥ����C=���{��ah�(��E�/RѝB�Q5�I[,��ce���bn�W<;5��j(�a��7l��K/��cG������#���*�Jn&��ȥ�ur,�&N �I#�bg����v��&����k;u!���%«"�JAW�1���xG�s9�妨�3c��M���J����E��l�6�㙧�����5ת���ZYQ뵖X+y^BZk��ʲ���Q�@���徧���m�]�FQ��'�|C}I<��G�innF*t�ލ�`�\B���T�+Bdw^+�yݒ�)������0������I����?<��4i?��Z
C�3]_�:� L'���.z=��y��^��{8�]x���#��{�S�H�{O?{�zLKrmPJE}��w�X�Z]���0
�L��g�7��u���c�?7�����+V	�럟�<rGlhǞb�T�h2=��ƣ�YSxՎ~�-עp�z9V��(6:�(��L��w߇y���3�1;;+ecV���j3#%�����f�A�L��"�����	�͖�FɺԯO��q�J[-���u�
-W:��1����h�dq������3#���Y�o���<o߄��Jf7,��/�#}X^\B�T�L����ķ��=�4��ˢ$U��M[q�u�������~�)���g��'>�)!�[}i�,�Ev�3�9\rե�21�4��RQL�?7�Q�!���I%l0�vd�z��x��{�tnZ��33?����8p訴�����<��_��O�Po
�|Í�����fF�<�Hx��v��V�k ��,u�,F�K8ۅ�^GGU�x#���`�*�g��)�#���Q-z7�U�*b�dҶ�DZ.�5�D�*5k]�WՔ5�ka/3٨�[y���-�<D��AL�p5�4��uA4M�]�-��^��S�Q��r��5OZ�g&���:�w�er.�g�����HzQQ#g���I�*ed�{Q���&'ӓ�l���k�@��T
~�&��v��
��s�t��$�iv�XX	�ky]�-��y�ޙီ�l>����k����H��U[ym�Rg�|ݞ={�8�'%Sj
t���Z19N���nB������Tq�L(����cc�Z�=Lm��2�N��Щt����Y!�w�8�c''q����ܲcu�H�^Z,"��G;b�R��ǣk��W�l�X7��<��'��a���_ݤeP����쏯T�1���Ȟ��\�6�;LTԴX�/+,z�CA4�.�M[��t����㵔X΄K�QU�� ������E�B�ť<<7&\U�vEʈ2�+K0�tB]j׹	����-�N�jCZ�̻8I�Z�-����z�V�)��*2�����ї�#�3y.�P��!1� �b���p�R>סN�=��i�G�.����]�e�4��?�AD�B�&�K�A�Zl5��\����~�����z�N�nGj���Q8AZ�>�7�צ��DU���?���X�x>4mD�N��V�ց��� *���������1� �_���_��+����_���3�q�%+ņi5؎l�R���6��<�ؚ�o�vO�p"�I���x���#�%#����߸@�-n֦�Qp��Q}x VZ��X�j�Q�II\qJd�c�1�Ҳ��f��L� (��dܺ���fE���q��ͤѓL�]k	H#�#H���(�YZM��
�nَn����?��lV�tQjb~nN���|���wÈX�,�[B_<�[���}�����#B�\��E�v���~�����a$=L7j�h��k6y��6FwlB<�@�UA�]����[]��1����s�ۀ�������!�A�X�f�������qd��t�M�oȢw� �"��<^{ťx��W�U������gav�����U��j*�&�&
Zl�z�=UcSg�b��C���?.\��q���6\�L���2�0�' "�i���#��SMܖKU���=W2R�\�>���T�jm:�\��l�RZW�n�6�ݵ�W��A-\I���[�)��iaCM�@���z2\������]y�G��t�H�?7EQ�.�E���K��W�t.ٹC86y_�Z"���S?��}zqV"��@f�%Xv�N��ed��xK�~V`�cԛ��6J?zd]&r����ɴ��0x�b!T����т���zc�A��4E+C�4(�㜚e�k�"���l���ߵ��J����5yL �
U?��@OMr���(�NN _\F�Q�+�R
�Z��]ģq4�6|��ۍ�p�hw\4�`8���(�B�qCt�8n:J]��숍��"z�br���16>���i�-�+jB��J��D,)k����W_#k���9lٲ'O���s�i)�NO�^aŗ��m���ާ� )|M�B^^�2��?��Hȭ l��FP��&��@�׉��H
)�H�|�CZ"�+�e�tQ�^a������F$�oR�,�����J�<��Ka��乎�o7��ɏ��4+��\<�y��l^9	��ӜG�Y��TX��U�"_Λz?�+�Vk(Cuzi�����������`q <���c���6���u>��`T�C�n�y:��v%��[���c��:>��O��`�R���t�4cC��>��X�&1e%<��W����aX�� �o�s�՟���r�7_Z��aԪ�9,	�bӨ��3�}[��7_���)���T Oe�\k O�s�O�:�Kˢc�- �7P|�d&�*s�LI*b�L�i��`�y�,.ѲQ�tU9Y2�1j!�븨���X��Dc_2&�0V�,G�:���T�M���~��FM��,//NOcfb^����b�g _��gP\��#G��c��j�����<�XOF2.���[�؎����[p��qQ%��^,㙟=�'~�St�6
���͛�����"��&�9Db�[e����&F#Qt�u����p�.ݴ^���o{.�	�T�v�r�����G?�q�sL�'��@=�1�k�V	��Y��`г91�/c!_C���{���:Dȓ��)J��\�E�=湈G]Ѭ�&��lH;(G�\���ii	�A��E��	� 9����e��M0^����
�9"k`! �]�z��O�Fٔ�6�C�i����:V!ۭ�ٞ�O�㔪���+�	ω�����.�B�V��j�k�J�#�i����Kϥ%��]��g>���S��/!�K�߱�i�ŗ^wމ��d�F'�8U#�:�*x�����$Y;���X<��^�;��K�����H�-V��8\���H��56xA%���L�-j�����>���|?W�aFV���|\�t�g5����AWp,��s�c;|�V��b	��[���#aE�n����M^2D..W��7�d�_�pҺ2u�"`�*���h�vI8Q�%z:�%^0^u:�:v��a5Yg�H�S���>}W^w�9V||,��I{,��$dq~gv�hV�<�9#�l5�h5��Wk�aF� �+m���r��iR�"�n���I�5Rm����	iJi�
��'�7���H�'�$E�`Չ�TNB&E#�2M\�Nf�튀�;6cin
�"f��7Ծ�q�x�΋E��
�G�`�?����@�j1���v<ה�!p� �`_?~�Wuu�
��wޟ��$1N�>�Z�$PO#�{���a ~<�������	o����±Iǫp�_���{
��S��x�����:h:~�dU���%D~ه�Ϧi}�q���p��{y�O��������Z݊a��s�����R�ͷ\��"Qau����������x���'\Ю��hG#��u��u���H��̌���J��h�L\��:cPb��pvn
}Z�����ۍ���b����X���$��H$�B�fI�7���[� ���[T���������XZ̮?��O�?��ق�͵+5!B�ŧ>����y�P�5���[���W�{.چri�޴�������<�T8��L�gl6l�,@�X/��,9�j�*�|yE6-u�Rչ"J��f��o�����7^v=N;*��ʝ8{�������#H�"�eHF�[-�K�V�#�B���m}a5lX^��6���h�����[Ҳ�E=x����*u5���#��	�y$7M��0+���/h���]�6�a�>���	��� ��^#��Bc�E^�D��,���R���`�2�@Keh����T��~|t�Z-	H��f���� T�4(ԙ�� �毞/L(EM�\%�@B�~[8a�g�L��7F�?�o�7�x�M�����(csC&�;ڏ�8�;��,�=�n:��A��*�5�P�c��Y�k.}���9������w�m�^��3E�D��בHΌ�L$0�W��,�BN��yJ���e�|}�V ��T2#mGm�"����뫕�An~    IDAT�/�/�����e�>h7i@΄,X�ꏐ�A�(U8&N�9�B)ä(d2�c��eM�#�an<7����
��O��:�ǥnE9vR���ʼ kgV�%1�eZ�A_/ZuN5Vts*�	�T{mGbB��{.݋��Y������qͳ-���zc��6��Z)�#1��,Ȩ0ONW%�u���|ip"�oHŋ�I��@��L%5�ʽ����rurY���S�4��B0Z����;�t-t}��i���"bG�|Jy=ms��*��!�0r�FF�ѬḦ ,����z����K�y[�r�z�*Y<&��0�&�bx�ʬ�U�Z�*��{��^-�y�=N6�}h�I[اX�(��kT�<��m���r`�����h�0��kܛ�D��$��d�~���k�Z]	ӕ/��+���ۧ�O����5?�F���ݿ�?_�v����;���wu�{�m��RD�b�]��񘀰�vd�7��ɣ荘dB����J�\��^t㞴��,n��l5!��"J�)VP䂅$5y��Ѧ��K��ʼ�*�R��L����1(���3G����SXa����TM�U�����ģ��j��?8<�J�&����P4��h��T>�v%:�X�\�q�+�>:��t ǩ���ѣG���󥢜�"�@�9$�v�n��M��1�	�f��<��Ν9����X��Q�[�)��0��{.���jK@�8zn�FU���b݈T�"U�f��.�h~�ַ�3m4kM��<vz��O�/�q�d=[7��I`���z��d�7��z�,7��0�m�'�5"H5l$:�hI�=@�Ժm�ṣ��L��-Tx)r��C���4?x��ኒ8�zQ΋�������'-O�pD�;(���td�����:����DI���Vغ ��ƙڐd�B�"U��B������X���r���)΢��逤�K��� �7�}I��0���J�����ݧF�ˠ��?�I\}�2�5<�AirJ��Qa�����>��=�(�Ԏ�Ƕ+�	��Y1D�I��`��(�4���>��h0��(��DkcmV(&�Lʵ�&����{��c��:Gj�Ӡ��dڤX��EeUeY�ZW�
h�yp���T�  �����R��e�@�O�Yƍ��]�'X	�5O�(igO�XYF$B�����C1cj.%�I�x�#�U�#�$��wg�U����-�]RP}*����k���O=)ߗלSv���H�ύ7�,U�cG�J|$����yҙ$Z���;N�sj�U�J�^E�������ɭ��* ƪ�ԲĜ;���Y��,�V�!�@�Hm�:�����������6 �Da�t�`e��0W,�h���$�FP�e���0��dG,f�RX�J�%d{[�bi�1��iʹ�A(�A˯�Jt�����	HU�f�!3F~�c�瞓5���_��_���Ӑ��$-�8���וs^[��i �c�>�aP��1�w��S��h ��3�z����X���Ճ.:~�;�w<��	���J_��W�m��ip�}r@�0� �/���Ŀ�Z�A������������o쒎A�X�ѭ���1>E̝b��q#�>�4�Q��-�\L�A1�@I]�Syb�f*8�!O�E ��*��̊�Bbf(���1(+E�Ucm�/eZ��
�#�☮������*j��z�F�J�/�ŕ�/o�x2�r�&U��U�A��b��m8~���}�XX���,�[�˸xx3���<��[��.��/���S��ɸ ��Z��+�@*��P"��C*��[������2܈j-�8wFl�J�b=�h�nD�1,VV�B��!��,�ʬ����S���]�]�#�
41`f��
����UǄ�"�`�Q2ꠣ�D�T@:ѱ��r>ur����w�:��x�{�����EU��7���׳����+d����m�j�k�(T��X����{;P�K���G��t����0>?��D��6X#^ �5�A瘟H�:p �QL.���E�l�U�`��(��!��6x��T[�"E�8��3w�t#8�7��4ã�j>K���--4��td�N�4� ������|^IC�s8�����\\�����-�c?��&�.��ߘ"c F����(�c��W�o�SQt{+�:)���0�xXtp�^?�i[���J^�}RE��4��(/,&'���F2p�~����W\x1��8�{{�yWj�� [Fo�k>y~��#�W���u�o�j�Yr��pV8�J`��O�#u?T9����f������M�bd��T`M_w>���x�<w�	�xL1^6Y��yޚ"� �@R��b7�+VȳР�U����L�M�񢗑,�%y?�>M�̦�ɸbTLH�ԬjF=����!��)x��A����B��G��@&[�7�&EI�|��Eґç@��*� cW$3)/�LOO�l�0�/�o�σ�p�t۶nK�C�����5p����ѧ�@,�жi������dR,#��?�NͪF�55F�F^�A����jvOQ~�Z�ݑf�8�[}�d.4��5Cz�rQ�6[՛��tʿY�lXXHʦ���4KJv�f���O�%�,Jb�����kU�4�'��Q��/ݺG�>�z9�R3�r|�:�dE�Y��xe>��כ(V������|FZ�,i�x\�g��8p� zz���#�-[�7���>a�L�%�4�ћ3]��{�����n���SA��G:��㌎A�@�צ����3�
p*��~O릓�����P�5ifPb�Ei>�S�� U��{tu�"�S@��sV��V�����L��@X��0n���n��C_wG�n�.�H��"
�i,[��9�m���/Bv� �|.���C�JU.ev�{Qy�;+ F����}�j"�"�ף��4mi�{������T/��]���=���7��d���)�LGr�dȖ��::��{K�!��;��b:�t:O8(���}6�oHR~�9�b��W��ƭu����X��c�-2��62�(�F�q���'�\j^v���Ɓ�G��0[�
[�ynҕ<�5�Y�
i��yD��e�Т�Rnh80�D�#�w�+A*����#���eS8>5{؋�׆L�$`����ǟ���� �B�B��X�m��j�(U���
,sdşMy	5,����C��eR��J2Qeggn7t)��򻤻�E��(���^����R\��hH��	p�UYt��PAKG)�J��_ZF� ���R�1�-�8Zӓ� Lο�ij_�V��@�LL��/V}֟�0�Nx����U�5��&�������*���N�!�_�C:�ܻ�q��h����G��
0ǳ���.�gxvf[���d��n�,�t$��A��$Aݥ�z��I����%̣n�M@�s&���lص�� �$&E?�ǤҎB� �#&�J1sA1qR�,iQ/4p$s�/��sl�|6^S(�R����Ӌ��ǆ�I-����ZÖ��p�Y/����?���N������8x���:b�2������3�°.d3��%��d��������ދe�K�������Q*���T�w������'W����w�K�,�SO���<�_�{�-l?�l<x#�G̔'��V������96�����J��ŮOj��)L��!2�=D3<z~�Y,�l>�v*�l�m�M&�H�Srш��"�w8<�V�wP� X���J��ZY≌c�!Vh���زa��c:R1L\�T��L�*<��.գ�J��V�>ﵮd|����ݺu���ɀqL��O�׽�url�O��j��ʐ�t��(Sj����AR+���Zo�ZA�R�?G�0OW[�c3�@���9��Ws����{�X Ey�L��3��J6t���U}����ٰFØv�|ߴX��{�������[�{c��;��e�SX1�߻�Ӗy�7�����^�yp�Y��IY۬h���G��Y�8���.�d4X��=��pI��0 �bQ�����&
WM բ���{�f����礭^<xh?��N��!O&����fi�z���Ŭ���z\��1�hw9�|�Z`c�9i��&�4i��g�H����/Ҏ6o^��t+���G���>V��A�+e�Xn�"���Dg(�����<�g�>~�xRv��F�m���q8;#X�e�v�b�#W-J (׊����������Q�eAa6��H��Vgo؂6�ɹz:�0��cza��A�f g���`<5���!N�F��R�(���tN*A�l�
��~�aG���b��H�nk�`���XF �vB<?>͊�U[S�j�i�m�D���]�	Jr����r9����sq�8ء��6�N�E���c�'8D��D^��c�`�I�����Q�/�
�*8�@�@�A�b�NN��Y��	n�Չ����@���Z��ʐ�4�/z�+Ph2a�E�	�M&,�J(�Q�t����K6SS�L���P� �j_�'3�,�:�킿3��ukD7�*4P�䐍Ǜ�|����h�IM�Ne�\���ML����t�P���	�7n�(@����=|"6�*ƒ�D.�d�+H/�v��Tp,�O�oddD���80T��fbtL@�k�u�T
��P��D�M3f��c��J�$��f'ƐJ��뢵N�����-o����\��v���CC��س����:�b��E"���� e2	�0�kXlnT+���b�x/+U��u�����Uh�z�������
���t��\,!�%=]�8:t=�}\ևL�
����_(�����Sri�A/l;
������b�uf؍�"}ZU(6�d�[z�Rv��D;1s5�R�f�9I��9tRA3}iX�%���}&3,��v'�{�����n;P&+�t
�KfK���6
�$�Bnt�����؝@1�*�"2�kMX����	;fz�i�)_�MOk�n*9v�ʲ���?�l.��kժ5�4Y��)�ʦ�xz���������g�̖f�ylv��OK���uT�0���PQ[�����>6Ǭ�U�%~������3{��8��.��Z߭?S��V�X&\���,���0��
��b�����z���n	�n�c���z��8V��#�O`�R7>��ע01�`��ŐܵsWᲡT-�^� Gӕ\݄�4�ƚ��y�E�,���b/F�����@&��χK���]"���rV/:2�[w�G�@��{r�Օ������K�"mth�H�Za����*ҵ�Aib[�aad
�C����ۜ��~��b�����o}�Pm?7���%Ț�E���]�6�ߺ���J��r��B>�XAln�?�fr)MN��&���Q��s��!sW,��b�Trdc)�NL�%�7�6��?v6�����a,���C�f��ׅ��w�����R%���dT��:<�>9:��lȗ�j����J!/v�X�j1Pci9�u켿��}�+�ߣa��h5�}�ǅ a��r;e�Y*��IU��Q@K���Sūvitw�b멹�9���L��b�����sl�Ν�o�Xz V��Rr:H)���sj�Z�S��J*�-f%9U�7��,�q�OͯS@�CC��N�BY������6a�F�G`�;�r�Q�)͓���9<���J��t��@W���vzð�kp[�C|�ÇO��엚&���?WZ��8۷�E����}���/��@ͤ����{,� �ѯ�y��c�LW� �����g�ɦT35�8a�Lk�)-f��jQ%#[��QR)�8S��y^�T;�z����QdS��^+�p�9g���5�(���q$RY��̓p{7�-[�J�A7=䋦�l�(���X�w½����$�N�*����*�oXJ�����Y��r����J���Q�y+e�[H�����ϕ���p��Ã>�l6/��'��jF�˺aqZ$�Iְ^�KK�5�t��qT�Y�w�z���(���w^C��T]�>�����j �)H�jSc( ���a��`���D���n�҃9)�'paz������ �`���Ȥ����8�{8�50cV���z3%?�% 㳒��1?���C"G�-$0ZS�P���,0ӑ�(�%�a ��� �7�k5�[찰��ꐖd��J��\�b���f�q�)D'̶f�h��I�f�ZS9~�{�����C�OY�����ꭴ5��^�7?�����F:����]����y~2?P��`JUl@�ҋ�q�L8^�8�1W�{Ɣ��4`�����xۓ����a�m.���tGu#�p;Sj)XKc����	z#�:k�*���l[�`C<e�a&��.��F���K�7;���HR�Ʋnq1V�L頯�ܺE��`au��<얺`�������_>�ɲ�RC	`Y�l���f�V������h��	Ha��v�{{�c��bJf�P�"6:���hs�`�=�ʁx�[ފ��.�ݽ�w?ƇNH��|)���y8=^�\p5��{�X2Ї���"�Z���q�:��y�|u��8|}t/_���Ȧ�
D8�9Y�X�3z\��������@���{�|9V�,��e�D&V��7�<�u��h�Έh�\3��GF��e�Uj��:P\H�+Ԏ��-���ȳ�%�&��̲0'mq�]*Z�r�[wn��۬���@5Y��:��n��U�t���.�WL�p�|	�|^�V���.0�����
�a��N������W�qUŗ>W�pҺ�RKB�~��T���#���(Y!mi�,�[fJ���tuW,σ�o�LBҲ.7>���g�vltl+�hP8CG�V?>�G#�/!�F���\10(-pj�� �T*�R���5�Zdl� �)k2(d��Ʊ+�V��q�a?I�Gk.����d|��ɂ�ؒs_R?�����ɫX���<wǢ+?sɒ%�T'Q՗��4�6�<3��3�?K�On��G�WjL��R�D���᭑�7����j�7J�$��sOǥ��������ҁA�u����[*WD��C~�dJػ�����**�+Vaד��뾮������ֆ/\�9lݶ�л|��A{[H�|��L].��w���f���}]���
������~�;�������G�7�J"u�� �l#7�L�xR���P�\UڗF��,���Y�����>[5n�ԩ/�K�6ǔt91�?�)��519��H��>��������C�\G�T��B
3���@��H�Y�H
d�ZQ��VB�mE|v~�S�m�7�~�L��,
ϙ�����!``i	�g@oo� +���'��'=���zl,�P�C����|=�Yb^3�jx/�Z�<��\�Ĝ�B
�X�%L`��W��B)��h'b�y���p��Fq��Q/YjH-�_�T"-]���Ւ�o|rL������Iu.�#_ǝ*A���ϙ����5�̍?y��?�2II�sͧ���G"����
s��D���O'����L��tu{����W��t�g�Ꭿ����O5�}�^0a���|�����oּ��U6N6�D��a�Oa��6��U�/ Ϧ$x��6TsY��Z���G��ԩ]�JGrW�pyqq?(��ܩ�S(�/�
�j� ;M��4%`��f��ø���1Zta�d�砎����L<�Y}h���cw��1Џ|E5o�yyj�����ؤTJ��T��嬗�-������	��-���a,w%[���ԧ;�¶3� ����������W�Ы�É��v�/�sU
��L�RK��*�N�P*��F�P������R_�v7�|���30еDL9����˗![.��!��%�������WmT�J�X]X�хz�*���|�l�CX)���V��\|ޜL:��'ت)�%�8�ʴ����Z-e`V�
�'?e
o%��.��b��45`
imP�PRV&3��j����Pͱ[ǮfYD<�&�f��_a�#M��`L����u�MK%�������f��6K�~��;vT1aAAf�p�W�q�'��r�\(���GچY>r�R�
)Pa    IDATu�̘�$n$8=8��^����WUm�te#�(�0�=W<��l uw�����	��
��Yɸ ��N�vJf�:�����	*��@yqM���s~�jXI����>�+�]y<��daL��9M��:�N�S��=G�y�=W�ZA�`���l`~v�t�M�4Jx��o�_]�:\��/�e���W���;����Awo?�bI�3���E4�&}@������#����yU��}~����8{�V�ٹj'���+*�+�R���y!�C$�e�:HZ1��P̂�g�ݏ��D3x�w��G�( ��2�>���>��W�� ��% �Ҳ[�i䗾�|V�흨������n���d�K!�G͋�a
�x+W��.�}2vK�.Ömg`�3097���Ǳ�g��&fb�ĺ�D;�D;J϶F9�QG<6;dӲ���](s�PN��//uY�=2�n�$@�c��hՊ�D;�� �֘�
�T6%�P,y�i�ڵK��E���矏��q�;7$�"�^�gn#�0r9�]��c[UP����P��E�����V�.���	yY�u��	�=t��	nB�Z��s�!��i=7	�ue1�ϓ 3@̿��nZ���rN162n���O���3�*��u96S����KutP��V�=>�r�C�]7{^l�|ތo����ෳ��F����%�,E�k��^�@���5{iQ�a�}]�px܂��x����jz���fCQS��zPe�|0�N-DV����C��?t�&@�6�8u�ڵ0JE�CK*�N"���{7��M&�Ϙ�d/+6���e�9ȊX��ڄF�Nַj�jWD[�J�r�xB�Nfb
��K�5��R���q79||�D�R�h��5�0J@�+�p( f٫7��+h���4R�4�=�\�{�@���e]�e��u21�f�X@2�L#=Cblv��h8v�d�P/Cp�s���0F(��d�*�x&�d6#��z{��mX5Wƚe�(���:�Z�&�_)]P@�.�Q����*��f�Z�j�� ����?L5;�3S��c��a�� �4n6�6�N�j?}���A��ZK��*��N�/2a��x�:��SZL��d�0��xOx�r=�ɒQ�A�B|���"8�/��ꫯ��F&�i@z=��-��9zBGI@�֠��]��?����R��b�cQU�� �i:��G�&j�LƋ���EIWH�a%���P �?��S�ކ0R��0@���sQC(���3VpA���������u�<��f� ro�y�#NoZ���T����	Sv5T-e�Jf�5H�x��*�4��2>p囱��3p�n�>���vt"����g!�e
��.��6�Z�r��h$�x"��Wb����/}G�-T*�L�p������Qm40>>*�h/��o~˖"67���.qi_��B�!aF��Y�;ڢx�k.���Z�ځ�{D�B.ޯ}�q�9���_�gY�)QP�k�RI*`Ԭ�#+�Һ��TVZY�����E���Ǐɘ���g��R��7��R�	cOG�����6���ɏ-$p��q�����>�)\�W�?��;�0O��}��u���P��6�qZ�lT079
/;zs0�+3*8t�F� �M���p]Rڶm�6����YI�v�ja��:t����Ue/�w,o6�����|@���q�S�gReII	���kO0�p����i�7��-�>?���b|+~F���g�g�9A�X�C����lbB����s�H�,�[��s�{9gxn\S�;�A�i�-٠&.
H#���������l(��5tjs�u����K�۰������F��%�� ��w=���Ϳ�X3`+#�|y}+���t���!57�Z./���j�x%v�iUM�l)�7�ܕk�k��h���R��ү��s�R/I
�QŖ5+�޿��
�4i���\�v~��A�r�o1Vrc���U���4�6جB��0�ހ��	����D�'Ss\8��{V�x2�����_��p�����-�f��N�"3�@y:-�2���M+�����6>�³����JY���@�@|m���(�����-�]�+��,T�r�ҳq��y�2z::����O (�81��Ĕx��9��c�6�L�ٹ/��J.���=��,�Ʀv�a�(er�xCM���S4�|�&�IC<��h�('�f´MK�	��X�&#ƴS/�Nj�L��b� ���gS#h��o1�߷�d9��[l_�N�/�#��i�G��f�;�*�7��Na¸eW�&VyV%95=.��Z]Y|���4���(����fU6���9|tH�!�<^�֮�nx<>�=~��ϗ2\eK��u�'eP�z��
J�[S��Zs7�v�c�����l
@1���sq�b�k���;���2u{y9&&���-�j�x.qv\���p�Q�q�����d���4 k�.��|��x�J|q�_aO���
��j>{oy�%x]��ݎ�~�s������`v7{D��;�DFD��
C��0&.�3��㟾(#U�*3j�ǫ.=O��}WHؕm[�`lt��NA�X^�332Zd�v?�4�c��m\�7��uD�~є%�i����{�n��^����R��g�R�
�0ۯǫ���5�f��D�xTu3����Ϝϒ�4�+��M��b�U�>�Lb!���Uk����{�U�HA�a����M<��Y����"�-���a��բ�̤s�����ܒ.��N�%� ;�(3v��Ǧ�&n<y��Q�ܱ�&77[�����>�_�@XR������Ās����F�� ���� gϞ=�CȖT)��L�q�����k��� �s��m����|6�=���5|�jC�W]�στ�����y�|֏=���Y��|�Z���t��F%��<�n���r���Z8�x�ody<Ͳuu�ȵI�v($ �ϓ�����������n��嫮7#�?��;����#)�����f��P��a+�#�le��F``w��h�a�E4?7czu�P��K��e�nNv��icM�(k!�Z�+@�Z�	K�f��R�-��Y�*L[� g���A|��(��(���k���,N���A��/��MhP�+�\� ��M��ᴱ$�	^'7��ތt}玗�O�|��\�����W6j�8(�V��g
���]�Í�-��d#���'�êͫ�nwa6>��l��9�5���(�z�tQuX�p�YpZ\�9���|<unܭs�x(�,� �˕P�N�L_"����.)����8r�x
�lǇ%������f�K��f��Ax.����z�	̎N��A�T�4��t���Q�E�M�ݠ�[da��#���i̲�6M3�[�d��������������K*�J�� 
�)M �M�%��'1`�q��U��j�L_��&��ӑ� L�T��R6{H� ���R�&;u����3���6���������a��i&)���U�ٷCǇ����Y�tׯ� �V���͓������XmG!Z-(P&���EL
_$���S����LKZT��s�`@f`�e���La��fz����&L�$Ɏ�*Ѩ�G����A�L><m����i���1���.������a5C1aԖ��f�Р�B)��ǂ׾��l�����?|��X��_�~�h�jw�����;�!���B;�D")�HM���'�O}	535N���k����t�0X���'Dϵe�6���/ �?�_�䳠� �S�4��lN�V\�Ob�@��F"۹{�[�C�
ֳ�:��ܵx��]��7��I�G
�E�n6얢1ff�J]��Q�J��9�(X��s숰���![�9L�̊6ꪫ�/����n�|�{��BǇGн��*p��F���D���06>7�Nٿ��b����Z1�F��D|N
}X���K���N~�¼�����FwO��յ��`��A�G����hU+
��Ar�q��~q<�M��$��P+�q�9�1JM�-3����z���vy�}�\����V��E;�-��9��dnN�&sͨ�	�8F8/������&�JYL�9�i��c�M�,�Ȧ��3A�4;F�~|��}���P@�, -Y�{��s.�r_������������F�a��O��w���`���
iXYd*SX��5o[^ZA�I������-�}Á\� ;i����%b{���z����gz�p�18Hr%�2��~�] �����>�����E���ˮچPX�zp���L�u��H&�&}��,�RdB��*aS�N���"�&ub�h������b��q�a���:����)�V	�Uj����!?��'��t�3����p��1��!���h~D�m��?�C��C�f`>��a���3������XJUTrt�B��X�֋J�O�'V,wMB����.L�ĉ�B%�E��PG�nƖ�[��v���c�K�c��g��M����\>�SlM ���te��@�s���X�Ԡ���n���GfS��b�t�L�n�CR�Z���A�A�#���\�*�[A�E�q1�R0��ϙ0�z݀�\8y�S|.MX+�ө2�;I��ޑ�~7��}��1�͋Ɔ1���=�E��jM�=;	�d�-<��.=1
��-j����N۴E�m�]!���	|ս��C�."0�����;]�Mt�炰u��SSr����<�"Q;v���FQ;�L\�@��r1!��5��������	�vT����ul��x�Q"�%,�Yh�65�-a�?(�N,$�a>�Z��^�����X=8����g��U������>؜>��A8=~�
e��y�<~��81,������5k�g�a|�S_/,j\	
hwpݗ� ǧ��u��w��\|�Œ�{��������z9�.Y��x�Y�	��?���p�����g����؂;~���y�w�޾����ص�I�sDQ|��@��2���ݢ�-hI<�����Y2�yO>���Y�0m!��:n&�v��!��C�P��o�����'auz`w{Q7x��qXl�D.��
��/^�z�zl`G�%ZT
I�4s�_5�]���<�������
�����O�$,�2��u�P�!�����-��?A�7�I��{���:Yݭ7{����ѭb��VL���g�_X(@y����s��F;�͙���vc~~V2�^�A�MY_������#x&(�q٠�ϳ�w�X�P���)�:�aUr�hǎ����x����d�Tt��M}�~���A$��48�:��7o����k���c�m?z��[����\��%v�.��F
��$Vm�Eŕ��Q��n���T	2wk�zAZD������K�� ��|�,�� '{$m#��$t�ܺ���JD�
��"�h8�q�om�UNcY�_���a-,�(��ٱP^u�p��G�Q��*�f1��^;�n�JU��)�|nt�����>�dV
&SUH�z����y���1`�><�S�G�;��r8��tG��x1�y%���%cH/�qp��u¾��t"��\.%l����X@��U���c녻�-��Y��Gfz��>�.���NVa,6��K��Jٰ��f�'��W'H��f��G�PJ���V��e���l��u`�uH-�)��� ´p��ӁJ-�u	�M�J�d&0 x�b#�>���١~�]�Q**�ǘf0�b��Ŗ+'���A�~v
x-�К�DfŰΊ��Q�Ȕ����ŠUt�^���ο~�h	���,��y����������Q$N�/���7�~��ˁ���!�Ҥ��s%����LA�Ī2����u��bjzӓʗJ���0eL��g�UF. P�D2��Y C���`��@wr�3���D�r>\�0_���c��K��	´1���RG��~�u��uY �<R�j�P��-��۶l�#�K����>H����Ui*=I]����б�
P���-���ŗn�QґdD�5V�eq�?_�W��e8p�Y�u����>�O�D|��m�݁cG�Ij��{�p� �\����%�]���?�[��&\���pιg��?�����.��Mشq>���b�3����p�݀6��M�Ԉ�QVi0�7�N���QE,�&s�m��1K"�Q����6}�Qd����_ ���O$�]v�e8xt'���ʔkC�P��{���X�#�އ\��b./�|��c�H[�n�d|�vQ����ڼ�_,WlN\x��b��L.����زe36n�  �`����
��5�d}�ܴ f6�9K�bV�*cZa�L�jVK�>�5��AO�L�t�j�A.�f���숐ʈ���N�w������6
�=��p���t9���2X�jɸ�Qkk�!_�I��W�5����Aj�a���8JŲ��˗�Z�ϥ��켴��qx?���|�u��_��Xԅ:���*�ل-�z��xfW�{_�����|� L��p��Ç}����u�/_W*�`)d�F��8V�ދ�+�����F��b����lz�bJ������ M.����ܕ�>�*�e�71K�
�KS��p�����'>�nX
1Xk�ʕ�_�QC��ǎ��AXE�Xj��06��ܷ�;E��귂�`W���,QK��Hk���7`-�Htq�N��[�A5���P�K������5��TC;��;ځ@W+6��-�Ĕ�S8����"�0z�t ����,
l ni�gI��(��_w�l����J�(��!��'�0sh�JC�]�O⼳�p�0?�w���pxݘ��ap�ji�44rB(�@0���Kaa[�j�D�dF��zۻa��´��Yl3��
3�����c�4�L�Ӏ�	����7�Q;�.
lnSI�6��I�hXX�&��-I�'�f�:̴o��M��z���@��C&L���u3+u1�Jߛ�5������;Z�#Gabb\<�V�Z�h$��/V�a��tWWn�N�8���iq"�����B^�I�g����)qݚ��л�;�-b�ϛW��3VBZ�$�����>��Fa��&�ˢoI��_�A���z�(�a3Y6|��l���T�ͧ#X�f~���czfR�6?��5q��bڄ�6Ss�"���@b����v�zR�J�t�=j������f�ת�?��Lʅ
fg&��r!�K^vV� Z�%P�S�F��պvS�^t� ������P*��-�Ic�����=�­?�Cܞ�֐�)�W�v�h����K.�����rC�{H�qrr
�����K02<�;��k�.qx�X���zgo)^��Kq�]��=����o~+������g�뙧����VRβ�1�Wi�*掦������:*��e��`\6�C<����B��A3Je�R]y�R�w睷����կ~5���f�b�W*�u i�#;�����ű�c��๳ۋ����ހ�A?�lV��:%�
On��ib�j�
iO<+�&�UU����M*��X�/ L�n��aqÐ�<e���X�z���%
Sh�0���Y	�$-(�`�:a�kF]WGr�q���H��z������ۺ(���ܴp=֖0��sJ�{�l?�_�M�x������	D5��ߣ�v4#�Yg~�f�fj���cq��@[�[yl^����s��׹\��È� �K�e/��	��'�����~�u#ܿ�� �O�QK�X���-ݨ��9J�9������hԩ-`�<
��f����rPP0-�$���Y�J���q��]6}��qk��������r�k��,g�ii>�W���G>5�XhO��*���;���8���\���5�����b�W���AVfu�0�z�45A�B�$?� ϛ�}�8���,rٌ<:G���P���g�i�-�{��?1��}��;пf��,�+��A�\
��G�ن�7���%p�����2)l<m��-JՐ�I��1:t\��ڻ������a�.���4��>���KP-��[��n�.��869��g�=K���~)���"�f�2k�L����?��H��"�!r��yS��4�i'}��    IDAT"ϕ����	c0�~[H��J!Y�iDh.~����k�P���M��Ё�LWj`�C���4v5w�L(�
���T�hEL�ݪO���{`T�[a�X8QUl�b��ԙl�N�0_:��k�1x>M�Ƽ����i��d����czz��6����W��el۶�x\�St�/�;7m����w�U�����D���/����N�"LXr6f^h��4��HF�d���Y�⢢��6�*� 5��⃯!��s��38oظY���]P{S-��Ϟ�4�WMUFƚͷU4*c�s���¢��;<k�/��L;��V��� L^k�s�VU�	D'F�0?;�J9�����mY�}��/���)Tj� ���	a��-���#�/�-�)c��^~����'��>�X�4­��}�_����?b!N1�=��`/��YDW�Z%����׳d�?s�����Oᓟ���k{{��9�å?�W��b�������հ9m��{1��H�!�)�7��1��.���=��Q���N+ӫuE�s�1�4���� ��Uc	��moƦM�p�]w!���=s&ggp�;0;��+���?8�щy��ٰ��%�~2a�K:�Lw����З��T>��aI�/�f25Z콚N'�N��Kʖ_�@e�L]�i�,�֕73$��3���y��l޼kV��4�fxy�O�;=F�Ѱ��� V�_0�r��}*�Ym4�{��s�������z�Yz�����������%��d���$A�����S�QOǲ��	5��ρu�a5��5��0�s/z�@5a�v���߽�7߬��6V�~^L�Z��T�����+�-+U���<4�s�Q�dQ�fa�(�Vq!�-*�9���>8b��ԠL])̓�i���jX����*\�.x]N��
��ƪ�0>�����RB��
�k�Y8C���;�_=q�S@�BLmlY�A�(zDH�g1k����k\�]9�uF�)�EOe���ۘ�H���0O@�gy3+��9�҈n�P�y�O����ܴP�m���1�M�>#�߉ޕ�p�XX�Ev>��{� �lGg���KQ�60:;��Q�'���ݝ���t�/����~�&�(�r�����֗���Ԉ���,��d,&,[{l~F�'������d �5QO�p�cw�3�%-�x\�I]�x)�/q�rQ*#[�ޟ�'L��O���-B����hL�%[R��r5h�g������0�B��&�%�Y���YԊ�]�H�㨴�"���M f�fy���� ���
�tP��� �VEa����]��Q&��S�����=�s����2~��y|��Ǿ��D���'dW�q�zy��d�	��u�^��a�ZX���m(05wl<��*	��G��RԌ�=�Fa7�h;ɕ�K�9��$�vVl$m�A��p��© [UR�d Tz3';l��4P8ul�4�d����J1���a��B1�\M�M"�I�Q'kQ��z3^v���G#�_��Kр����T���wjU�	;Q*���D�Z����Ń�����	p�m����q��>����|j'I�QDq���1yn;z�\��1��}W���f����E$�!3�����go?���lټV�QbCQ���w��G�d&!w@k���@-����̦����֤�]Z԰�c]m��(�IC蚌�q% �쨢{���<�igZ�HS��q�&���L�t�w1�Ƕ���>�?�b��ݍD�]5�����j�`/��S��uަXp��6M�ucz^�4r^�&�(�ρרƒҗ���ju�:L�_�e��A�^��K��� ;��(3D�o�=
t� I3I���|��|�$�j�﵂:���,@`�j�Jo4�n�ha��UA�b�U���YU�Wv@Z{�s�W߹���i�7_/�ٔ���a����%��[���/Ff|��t���Upvl&���hT(c+ք��f�@{�r~"����,R�קʒ��
JE�-`�
�s�d-�$���t������ۨ����y�K4��pP�O��l/Y�o��Rxl��v*���E��H~p��q���q$m��U��҇���%��%��A�0��-�06��y �/؟�Z� '�������6�E!���3�K�|:6'���ŏ�d�c���Ï�����)=ñ��p���ً��#�׉��b�6]���3�k����a��*iU�� CF6��o�=�6̎O⇷�*)�c�������H{�D� wЏ��R�t^�ζ8�6x�^L��R���*��rKM��&&'�Ye�@`͒�@nZ��fU��zԻr.@�G'�F�ˈ�"e���A���|�
|J�N]��^�8Z�8ٛN�t��fAR�&�Y�5��z��� L�3����0�eb�	�( �Z����w����׈0�0g�'���EŔ����OL�����(SV�ϋU,�'� �*�Z]��h�T�h��1]�q�k'�6L��/}�+�?�#'�������KХ���	��k�E�c����P@[�X�9%G)�E �S L���N��ܤ ����ry�l����ʄ�q���);��Ud��d�N������$:{ڤ�a2�AO�RX�.x=a5�x�a��ۺ�ϕ��W[�sր8�S���ދH0�����}�����[�%�j���O�G?�2�4^��W�Yr����Çp��a��ud��u���\��o��P��{��O}�6�E:���'�(�袋$�{`�!��=�Ǉ���M�U��S4��ں&�5�ik5�t��VI9n7���.J�zf��bQ����7�CΏ��T��-�p��a�#!8�^ܿ�!x|��%KgỤۇB>T��]�	�1�M&�,"Dy�|q�n(&�	�أ֡�De#lW,ײ&3���a~9��V�5��oz�_���W���g+k�H��l����r�R�u�TJ�N�>j��ޙK����+ԺU7���O�X���������(�O�M�)�� qs�� V6�&�"��"��\k�4�졾o���f�lX�������0������������%�tﾳn�����§Uh�Z�I:�aİ|��3	�5�ngg�Ī�.�� ǂ�N��$Մ��U���K�L=��zgu�-�&�jq��9���q�c*���t6��ύMkW�V���^�U������;w��OƱ�q�@l�x�E1aNqy�	&=��td�=�4a���j�ܨ�Ĕd�$�K�6ŀ���b\�V/_��B\��gц�q�vG����~�jX�̌�`vxcC�p~��:�5Џ��z���Gِ�]1{�N�ry���T5?;�����辸��uD{���lZ�V@�C��P6[�e�G�Ш��\|�'~bR]���Za_P�=iM1|�¾�TT��y3tj𥟝�L�m3Ķ0R��U�:�uQ��R�Y�2ZK���sqt� �fU��@��Tn֪
O�_*�~V� �0���5������S��L�SS`��.��[]���!bqj�k��@�0�~��s�#i��s��&�S$&���_�7]�W�J��� ��Bx�|�S���3�5<U�^�_2  �M�*��� L=�S�C�	���3�묪@�Z�*������s3��M��JI�8
k.iJ�sYڿL�+b��i.$\��77xiԘ���*��d���d��3���突{�3:�	c�"� �tY#�M$٣cGNy�p� � ���7�r�c�*@��|��T��l��r|�V�` "@��O��)�Ҋ�֬���8>���������س�)�zj�����/�%�\�{��P��pJ���u�a�y00����;�I��&�b�_n�"�x�:�c��B|^2O<��<*P�9d�	�����9c��Ts#̿�>����0����ϟ����1Ѡԩ�j�H���J�rRm���@�+����)�?x�(.y��aX����=��ΈU~�J]�*h�	x�����ц��"��K�cA���u�PqLU+��R)>ѻ���Z���"��K5w��F�Z3���WHK�Ç�L��Ӈ�Y�㑌��x�8��|��J�Ō�K�3&�,�і����u�f��_�4t�^�r��(P�1Qf��2_+?7�_ZXk<?	���;A�-��/J��{vo���~��n"�k)�j
0������Up�k/�ڮ¬� �(�p4P�����;10s�z��I���(X?LVRZ�p���N���%�%6��?��ݨg�2q��Sa0`��P�}����C8��
��
��S�0�#5kՄu-_" �.e���шV\��d���'��&��~4��Τ�0�U��@u>���<���J��j��@��Cvn��s���ڜhx���}���ɉ�)xmD<AI=��
��J�r���|���}��6;��8��M�=���
5:gS����0>;�x�*D��72�H���
K�W��z��b�H��\�͸��������d@��N=�[uTz��h̪�/v ��b�T:Q*MWt���bA4�&��&�BG���EC1K�\��;R�O3S��k�:� �^j<6����P�b�������W�j���ڞ�����c+2a�O��j�i㬗����ł��y�\̦f�q��1�/,�Ď|�V�TkQ����#�<��Ү��
����2�M�h��~�s�"X�0��Cǎ�~~V���0s�<�lFYM�cE��Զ���7�0�t������xLY1E�ԥ�M*��uRz���_���
X���,���1�0AK�8XjR�]��Լ2ɭ���|U�
�ݲ3��YifC0�������+F�Ĵ$�� ���۩k�P�����{����x����>�T2�?>�;l�~�l݌_�{/�ch(��?�mo�>�{$�Y�\���1�r�M8���0KJ�+e�i�o�1F��ᢋ.�}����2��y\�N�,T����r�t(��"@w�]*]R�&�C20�;���Z*�@i0�uI�H	
��̶H���%K��R�wi?��s��կ�f�F���{~q�}p��8��ӱc�ܷ��#ظn%���Yo+[���N
yd�Q������g�eV����� ����#sd�[dLӮ���t�ޜq���y�#����#�d�4AA@�:&Y�5^
d��=�^����;l���+��W��F��"�i��kk݄��YoP�|ЩQ�^��\���V]�|�Y(u*�%L���ST\T �j5�k�9��0�W��F�a�׻�8�w=|c�ݾ��ޕ���z#�U+|�O�%�¸���Ó_@XY9Xϱ�=,.H3o���LUI�j�-����-�OP�",w��Y(ڕM�I��� �f�rT��څ�!�Ķv|���q���8��!I&G�ӊ	�ҡ-*�w�Ʉq|0juY�38�b]/�A�JY�h�Ij���dUL���
1K���E��@5�Cn4��B;�>t"�����N�P@�fA9���|�1L'sH4(�E�C�|A��L�L]�2�榦�zp�g��gnG:���󼙒a�y��ǥ���4LGnZ��1T�<�o/v<�k<��I	`�bn����8��\�ms�FA��-�XDȍ�;��5��:良ӆ�W�0�7�qsҋ��T��?�U�f�ZE�4����+�:STk�0]�ô�I�I)���3��qY�� ȿI��)�o��cCF��?�c��~�kP;�E6���0_1a|+e	�h.��}���R�ɦ�܎��]�Fwo/
��ɔ4��ؔ����2i�e��	�4�A�~^��Ϛѻg~�٪�J*�SdVo���3�S��� �lw��<�0]AF�%���]&)Ϛ ��S����9�9&�:^7A�T/�����)fF��O�z����4�=�	� �]2��c�S�hR���l�F��6�6���'U�Ǐ�I�qؽp�=�!"����X���h6���wZ���w��0�>'����'��`�+i���=юvic�/���ڞ�����WJV�O#�+��	��㢋.��}�j
Y��C�V�9����c�(�J\�/^-���-1��V���RW��~S�OY�%U�"��A6�U���ڴ�S<�T���� L��2tL��#4�����g�#�G�#�[�W�m��z�d�+t��`|:������������?�#��oz�bQ���$H�g�iC��;s���_�O*���`�U�'��b��dM@M�"e�,J�䆢�����0n��2���!1�i���+?�S�V��uA���t��OR�G[��Z;�*��s����j��%�ikP�5�j憅���Gon�	S_��t���_#�n�j5n���7c�����_� �H�����]��_>�oUǚ��l�]͠V�����mƥ����=�����ѷ�&M�]v�P"Z1�4[�P0-�,�o��R��$�K5a)'p�)��3��$=&�pR�<p�:�.��֍���.ܿ�N���T#d�h�^�x'�� �Kӑڢ��4AS��RQ@X�a66�=���T�$e�A��*͑���ȍ�"7<_�)팸Xv,mömk1�²N���)����͓{�4쨰I4�É�BJ|�6Ү4�������B^?�����z./��w�$ ��6���g�Y)��b��f��03;��}�xl�Ni���z�.ħ��p�es�������n�I�N:�Km����^�$�6���s"�T�]OB=�[u'r_�j��*p	{D��Ls�I�@���C��R�jǩc��"�haO:�<�~��� ���켜w�b�j(���a>����I竟U�W���d�9�sg�mvvFZoq�?��)=B{z��a�:�[�Fz�r��%��!���yn!�L.�]YN�G1,�2b}L3����E�S��E.`���t�xX�OR��z0>>�eJնFW,�	�$5QL!�]�=t{U�̈́�y���W�\�&#��l��xzzVޫu`��|e��NNI�+���������D1ar�O��`1������Ѱ�{B��:\A�dRe_�#s���ç@X��!�$�Ɇ��Tk�
�=�L��i=�u�ۑ�$�w�3ؼy��֙��E0��}�3�&g��g�/�r���+�����-�k?��>?v=��\s��.��b��Ȥ�\�m.?vX��GdD�
c�S�/�D[4��+ϗ��cMo�'��zCL>���L�.к��h�X8�|~�̃���r��?}��3l�,�K�����pbd\�I�pP�]
(`�!�Ó�=�{~~7�>*��9d�X�Jk	2ad���^���P��PX8��&�`Cr�γ�^Y��j�I#s�yy�7�j�[��&�(�̓5�����x��s�)�7t<��PU�z0���c��Ѡ�����5�I�~j`|h2_�����a�sJ2W��x���tu�)�9i��n�U`ީ�C���>�a{gf�w�8x�Ow��+�`�*���l�[N�T�ř[zQKć�v	V��貕�,fP�daq5P��P�T�p�1��f(v�?����/L�[(�Oi�A�K]*�ű�����%v�r$o.��1ei��ދ���n<��(F�u����#G�(�W�J{��Q��&F�2��V,Y�/�92aY�^)夿"igi�f:=3��#�	��Ϊ�J	n��lsϞ@y,��H7�v���4p��[q��gbYg!�Sڊ��l���㷿G��B��B^R\Vx�.�x�|�7o�_�Z={{w?��윤��~ו�̓�Kc�e}l��N��``9ۧԐ�d���+���b��(v���>.i���^� �ގم�%e�
�����H��e�6Hu<PK�	xOM��@�C�;5��V�)oM�����QmR$1"U��ހW�Pl�]?'��Y��9K�i��א^�<z���p�;h��p!`��bfG�|Nb'��Ea�~��:�
�t'�?��,)ߢXl�GNHi<+���9txHRd���ַ��5��T�rQ����ɋ���H�n�)�`���E�i�	D��5��h"ŋ�dƿIj��v9��d�:bs��F��~.�^S���8�Y׷�W�.|�/���=l$    IDAT~�f���O��z>>���.i<�ry�)J~�n���f!�s�'ap�-�>���	F�)zU�q9�B�Nˈ(���M�{��U]٢��*U)�,���Mp �`0�1n�h��t���19���LN&	���B���ʹN����k���2����w�p�O_���9���k�5�c�	�3�|1���dea�(ȷT��x{�VT��i	�;eP����D0����+�pL*?��S��S��{��-|��ֆup����~��r/�DT��/�"�J������u��D0T���.�w���X��V$�e��ߎ�����N=Y6��<�����Bqz$Fh@�����8x�u�r/�>�q0;�:�;�xdd��&SIx�x�X��:&�����"���2�1�����>�q�7�U*��.ߟL�O�'�]t4�L����b���v�������}��{}��� ���1�׺R����AaT�D�猥L�<2_Q0�Cz=ѣ��R�]���F(�א��1m.��|Y�l���y�5*a1�q&�Ы����͌S0'�~���5��9��y����A�a�� �̆����l��͠K__-�ׂ}-�����n��K�X,ޞ��18�c�[�}��w�p $@ۿT��,V�(gr���@efx)u᫧�y¶�4��(�ҹ��:[ɅlZ�h�Cj�v5O�kT�+�1E���2���2�5�,I#� x�s٦/�D�C�
��85'm������o}��bV����gW��V�hgA�bE�*",�����F��f)G�+%�
9$q�'���L
��E�_��)���Eab�$��jaˡ�w1��޲~�G�\��Y�#�/�{o��#���M���?M>��Ӄx�)�RQ>���C��=Q�ٟ�>}�	p�]Bo���G�p�E���_C��tU��i��Υ�<�A�*`������n�z�|�m�I�bμ�2�e9����@0��? :f�sS�!ฬ��޺� ��Ԭ�:$'M��1�92��jЮ�8�!�)-��b����qR��<��tW�Yw�����{��U�B	V���A�����_�w�Zs �ݓ�)uBo4���́F>�<m���#m<�;;�{10ԯt-�����8�K�b���رcN8����{������F��i�������F�M�~w,7Ϛ:]lx�E��_�L\8D,�ϡ���]4@,E���FG�"�����=�3j�ds(A4?vt����F���y���XtDޟL�b�Ug(���9<�:���K�3$�^�t��Q���y0�8z3Q��*�,�Z(��x�Ir��~�t>sNa<1�H��-�3>}>u�q���v8�^lڸٴK���[���g=�
�st�f��� �|��l72;�����p�c_��<�{�x򩇱~�kȤ9�ٍP*-k���`%�Rym}^}�M���1O�։ ���.�g�~/���h	�FDjq��w`��7$�r�%`��b	�<�M��뮻�h�<i�ؽ�S��2��ڻ����cڴ�U5�<Ͻ�ر�9��y[�m����je��U�uZݨ���_��,�s�)�4<�R���%a�|n+��\cL2�9T
y<�裘9�/��<^}�e��2���4�g5�� �����d�Хm�_&�2��}�x��^]ۀ@(,�a21�����7���:��r��օQr���`�ɐ�ds|�3���򟊍*f)Vlb��d����gצ������eQ���/?���Nf��q}<V��R�߄������*RFC�A%�	F��ۍN����]9��Rq�q��z��M�/���+NT�$_�k� O���ԉ?w$�D\�TRpXҰY�p�K�q�6�8<pX����Q5{�E��XT]~Ѿaz1���2%�i���>\�&Ŋp�0[��VJ���;�ĕ�=�=#q�i3a�+٭�;9`��́�Q�[E�����pܨ�R��Y�~\* S̢(�'�.V`鑓W%Σd��,Lf�� ��F��Ʈ�!\r��.�� N:��|�aȏ���7��V�\n�<�0|�?�c���=��E��F�/�K�mNTY<8���p�c@',���f��q�>����MTW�����Í��CV�E�ޤ<W���
��M��#��y���!�*���wK`�͑ ��r	���k�$� �0,�i�K���;'3H�(6~c���Fw��aC��A�n��{լC�SkEw�̺ E���8̺U���j�#��3��R������V�R�� 6���������k�����sp.�r��Պ�N:	˖,��K-���g��GAO_/��Q�P��m�x{�&i �5��3�i�T�)F۾$FF�����fF��IX�l�u���IY�nP9;���Z�쓎.�==}��&:�S6}]�"��M�4K^|(f�!�u������K˔ir_,h'��t���&�'�ߔQ(�(6"I^L�u�ۉ�x]}�H�ch�����_/>^��b
+;��ta��}H%-x��wa������ǎ1�es�B�p�Yu�4)T����I�H����	'#V��r#l�"��d�Rx�G��5�,���Yc�T�}c#������y�=[0g��#��v�k����/�]���[���d�4��O}�D<��3�Scٚ��\Z��o��F.4ԇ0<�����vn�!,��eC��Css=��������ކ_~Ut���Jp��q5C�Z���N����T�M����m�p4�9碷�.����g��҅����8��Oc��E��B&�L�]�%��n֯_��6�Wɗ�T�ឮ�D�ھ�m<�Ru�+2����D�`�k��s��9�'S�ǒ���Zq����H�,%"NBPMFL�ɾ��$����NK���B|3�1�0��&�dMN����:��c�ʈ����A��99���W�|}���g�E��e+A��Ga��5o��7�/{���+N�Sl�K��!,"V<���z7��(Da)�`��P�j�]���h�����ë�M�%��w9��F�f�RwV��fj,ʂ2F���X����>�K9q�;���K�aC�z�9d)��4�revֹTG��/�d�@3[�ᳫ������b�rQ[�3rc��>LbmP�ȦA�D���k&�jоy0�����{�8r�B�~�'��$��Ɔ�p{�8����/�~��������>?\n��o6���bG�/�#���I�Vc����z@��=8��ӱ���X%�	���c9�SN��+��_�ʤ	�`,Ǎ7܌'�~J@����/���˗/��yP46�x.�]�ф)1�5DV���w윍�� ����1Żfvb"����V3������]ds��:�耥��W�5�t�%�A�8�e9�;����c|&�0sw��@��A���?aeY�� m�_L>th����M�v-S[��l�2l߹��-e%6�xA)�p ��b�X��K���*$�LZY�j�e��6mQa���>΄�ҕ�<�������Y+�}�t{=Xs�K�P��.K��92�j�F`�/:㓽�z2&�8t9�����͟�HJ�ez#��Q_;Y;Fl1oP�Ɇ���٫
���V���@}�O�[\���@>�@��-Sgb���@W?���E��@]C38��z����rHeh��F X�Jَ��=}#��0�I�	���P�����,ƞv`��S�e6oOg�0�C�����x�;�Vaמv�}L�9�W���G	�ۉy����Md��)-¤m�����w��yKf��߿￷���8���ظq#�l}�V����z������>��w5
Y��Wl�(^/�&���ܹsq�'�ͷ6�����ern�L��(\n+BA?,e�4}X+6�8扣�����I3;W9+�MA�WJ��͍2E`JCN����\���a�ܾ}+~d�����˕�J7������f�5��I��/)�r���ҙ�j�142*VLfL��/|�4�'�J�ei�D�Vv'kGz�#��:1�~u�2�G���Mk2�Ҿ~���y:��Nf�b�{M5 ��ŝ`�~G�̺��a 전�#���9�)�fv���}�#-�yxñ�m�MoxA��@9] J,��`�L���O=S�%�y�*�9d�I�<���x��װ��VOH���N'���ōY/ �0Ԣ�E_$�N��ƍաj�0\[ś��v��K���x:������G���H� m�p��f�/��-Y�� b��d(��	w��HC5��0a4l-Љ�2T)�%Qf�ܰd5Z̙Ս&��Pɗ��Yѷ���!�D�q:0��_=��۬X��߰��w%�~��K�e�k���t
�>�W@Ul8
K���;��@a��D� ���ÄP�146"�x{taۖ-R�#v�a����8������h��a��\/><��T*V|��ӱh�"���K��M=K�P�X\E
j(Ҍ��Z+�cKo|�L�~fΚ(�Տ�Y2��#��t�v��k)�U����d�^�K��	3V>G3j��$�J�E��5�:
p��Q���5>،�?�f��� a�e>?
�]�`#9&AX����a@����N5\�|����4����w�_��Ԅ�%��s����>�eV�֩2��̏ي=���&�0�4aG>��r$�`{{�8��<+<n��x��� B��$,�lc������%?��>/zm�ɲ"�=?�8�3�ʰYfb܎�D�&usiJ��`YL����4q%ńY!,�'�G_� �P�w�QL�.���ϯ{��?:������sy��o�5�f*�EӘ�2�=���O�K�M�'z�M�ڌ�H{��ġ+#��e���]���j����b��|�
Q］AX�t��-�w����g��%���Y�r1��7��ߞ}�w �.]�ݻ���.�tzoi��T���<=�)w���]�r�)���2f�ضm.��b��%Ѽ��E��q{,6�pPMH`�c���;����~2S���W}r��0�v7J��*[asx�(���^x+��7w.:�c�;�"%����CV��n���3i�����_����������3G��Y>�N5�ɑ^/f��eK?קt���.�LI���I����f�q�D��sb��Uf�J�4���80��4�1'�����M3�"����:���ֱ�\�ʁ��H����f \&�<q6�����Dg�{����z����cɄ]��[���ٵ�݁Ŋ�TAd�:�%�<��G���*G�r��H�bkG~y�m�X���)L�L	�(�<�E7�	����B��"�DL����r:�k�d(�v��(�H'3��Fa-�d�bC�ZF��JQf��,6��9��Z#v����`��@}�LB@X��MkY���0�l�/ᰨ:��$O��
	���H��0���|u^f�ա�*�S�Y�cW/;���0�_}/mz�6��N`G��G.����m�8
��dE��k��b����5�_�\::d3d�`G&�J�*$���G��W��Q�o~�;<�����9w�
CC�G"��|��r���r!�PY���&�,(&�'3����w������JW��,m�F7,7ڇH3a" 6�3��7g_��]��ٚz�����7Z`���,��u¯`dz�:)��Z�0�3��(� L5�g3����e>)�@��K�\K2�6+>سG��t8���M��G4EӴ�2����[�n��ب<� 67=�\jx�͎"AX��iSZ�6^�����aIb$��ϸ���8���fPWW+�o_�)%>9��&�\(��ze�Z��k�T�1���"f�7�����r]�:*�W����"���,��F��ڒnfSW����*r����(���]ntu� AC�/svq�w�K��;�Õ����ll�(���`��yr�E��u#� e�6B�:t���O~~�x_q=RVW[�֩������c�f���Ѷo��s�oE��<���i���硾�6����s��կ��T*/��g�~B: 	dO8�8��X�l���j��b�&�jnn�������8>4<���;�^��E���X�~#�;�|�ܳL�����}(�����^3m�K���N���6in������B�D�oR9&�vI��	a��kHаt�b��+gP,В�@̇�/>�l����aY�k~�>���0��16�0np�h&L1h4��?�}Kv\�i>�1�8���;]�)���w�*g����Q�c��k����r$��a �̈�9v��F�Ƅ��3�\�f?j�_�er'�0s��;P�!#��I�9�����Y�,�����ч�����+�}�
e;J鲀0�}Kf�)���-�]��$�l�-����Ï��ņ��S�D�<�j<�pܢM�¢9�o$.�
F�)�U�C.:��zK'd��DS%o��g�j�R9�uY�g	�����%E�CN�H��
\^���9�	x�"�N
�z\ldR�XQ�P�K0��7ˑ�0�NX�+%x9�(�G���X��=�[mh�U��|B>�2�<^{�M������Q�ර`-Y�v�������j)�-ې������|�ż�$;ƀ���1������D��B^L:	®��o�ؓOH9�7[KK+�n�%���@P<z�`���g��5�-��5�?ڦ� &b��7�.I���z�����`*�-����S]z"�6hx^/u��<��k�`�&��zLɄNB�;ա��_��lC6@3aZ'���@O&�����Y��3��L���9)}��/�.�"\�ؿ8�n�-I^��¨�D���%�1~gٞ�r�Q�X1n~%6��1��E�U�?o�q����Ym�KR5&�<��.�P�YEzNM�ڊv���2q(L����`,�'S�C
�ݲ��鍍^c�;�g�V���5uD[e��d3x��:���Gz�Ӭ?�a��W{r��1�HUՕG�� o��Z��Ջt2�j��� n��x������[�?�����d-y���G�d�P<���W���;�X��K��]��I��e3)aP��6"��a�t��^�1�Y-��?�+�_�g��n˃��:�w�� N8��q��X��&$�Y|�SQU����(�߼	��{14�/����.N>�d<������V��/���A �J�x�eS���>�[n�CC�i���ƓO>)��l
"�[>G*�ix=a�-����������X���V}�lK�.F0���#~�����aK6d88��&�pM-F�b���q�Ēej�tvu`$֋T:[�����w�|4�Ԧxo�x�ǤL�u�狺�wFLq|����jΑ�6T�)���?CuM�Gd_bY�q�1�/}u���R�y�l��M$�4˦A��(��������T��g��s4� Mʜ�x�A7U`2�����*�����LWc�&'��l6h\���x��a���^=��7޻.g��-��(�(����.u��SW	�.�����^U���1�����s�S-Τc� ��7:甸P�O,���cttXuy�RE{�Y��K+Ƽ+�d��C4���-E�-�
�ec! q[l�Ė����z3>���W��dȼA?�>'�R	a��,N���|!�6s�qN�2�d��r#�.� Kh�����!���, 9<&3��$j�8�%D|>r	�Is�����X�N$��lq�ku��Q�
'��li/Z�.Yগ[��H(���rX]j��'�����A��Q(es�f�l��._��L��0�d�PD�mAf�Cp���w�����&�`�`�1ˆ�9r��|��~/���6*+U�����tW��%eVg��\��da���<��A�Q0��=��p�i�� �:�h��f}����\��t�S�wAʤ��|
	Ĳ���0��0�Bf��QrYa�8�X�����na����^^@�f��e��V�Hi}jC�h%v�8��݀��Sf��1�u�&�!��q��*"%5�;��5�, ���Ki�|L���    IDAT��<�ր?�/K�[�lQ�� ���Z� �eb9��z��VќN�V��0l������r0|YbF�T ;غ{�����o-�8n���xꩧ����~�r5'��9��f�ᦼ{�>T,.T�Q,X��"�,�[�^�x2+k��O#
`���cg�߅O~��}�����؏-[6#E0\�������a�{���ƹ瞋��w���k_��VQ�;�M�I��w�� �?�'�9N�1���&�І�&�sc�1�z�gq��7�P?��=Ř������X��ɸ8Г�9��/�����-���㶋y�N�,b�(^{��@���SØ�`���8������w�dq�����lu��Î��y��cO"�ȢT���3�A*ǚ��CMm3Z[q�m��Ef;1�ݎ�o��;�C4aLD�ό�>3��$�	�|b^,�u��'�
YC�O�ml�?)G�����ۙg�)�0t���U�m��)��Tv�zz�ĬH���5��� �\��06Y��c�8����'���	��h����5�\N҄Mm���CFM��O���U����ǽ���k�V��bņb�74��*MXi?�r�*L��ew$�(f3���(۽�������E�;�M���3R�0����W�R4�W�nC3C=�����QP�M����Aއ�N�%A��brX�CVL���ԣ��_S���(6@�[�����"v[y�0����
�Ơaa\cUr��ġ�����PS�ζH�S��dKR��ǒ���D6Ŕ�:��Y���:�H�(�P�����j�oB]U/��eB58e�	ػe;��g	����'�(�2��8h�b]�h=��.7`:�Ϟ;Gu�+R�"���.	 ġ@S�O���(����ƈ�i���+͖����j�,����$���on�}́a�!3ʑ��L[�c	�4��K[)���t�Pj~�Ձޜ5XS��C{9�A�r�A����L�a:KT�hXSe����j}Oh���YZ��? a|=[�)h��L�Q[_'�J�/Kv�n�[�Q
ahp］I>�O�a.�Otd{R��E��ͭ�|L�\##��c�� � �N�,����L�c�%#4X��#�[i֪6�!�	�9f�#��T\{���z��KpF&������a$����:��3���G�0��d��S��`���/�@��]�Ȧ�*�V���3��o�{4������567ap@��ė��c�<Ѕ`��l.g@���"�������i����Tc���BKk=F���`�\lݲ	��^�iC��%D͛7_�u���71{�<iؽ�c�,Vv�t�N�ъё�޳�}�k�pڬHg�"$W�d^�����`��U��n��f466�y�]2aW^y��ξ� ��_#c�ز�]̟;���X�p>ֿ�":�w��ct��T\4�Y�n��4YfB�-��A�PNO�nى�x�TV:O{�q�mw���o�c�=%��V�8?�������b�Ƶ���/�߾�5�u���*���'���²�~�C�c�"c�ħRuCr�k�"�0��ye��߫8a����֭C�XFm}�Heƫ?v���Ξ3�RN���L�7��EFA-�̟�3�a��$Y�p^�/F��aZįU�f���c�@��A��x�$I$.��c�#�D�iT&�� ��1|�s�^0�$iv�6��ݑw~�4a]]]����z���6��Vΐ	K��~,��7�������p�����a���A	.���?�����]�#�EP[6�7 z��#�G�9l�d��"2W"ڟ���fKfG�e��C!�Ȓ:�SD�bAY�y;�U����$�D�|
�6�M��j�n(;�~/jZ0�0��#f�d�Ȅ�Ό�6;(��gp{�)���Ν�t")��v�ltY�b~Ktbh�X,=2����.��H ��-3Ze����(����J�i�'�8��,G����7n�민��}�l{��-���7/nx�\�����Ɏ�������ߟ���#�����
W���Iu�u�J�1g�0^+�a4�x���W2ï������0-��b����H�R�8���v4McP T;RO�g�0
^[NL�{t�t7�*�M4�ҝ���Z:�e��]%�=��Cf��
�,��2F}���f��mR�����n�9f�-��Q��t�����M��E��G�R��=�M���M����,`��YԆE�:O�:���,$� M�#�����5"��j�!b�AU�����77n���}cѸ}�p・�s�;>� K5(O>����i�e^?Γ$���!3{n*ZGH+
�,�g�
j���U ��F�Q1G�[U�_�c�PAo_?��J�(��2~t�`��]x��-���~)`�%=Z�#��z�b-���с�&�N�Iklh��h
���
�T��BF�VM�u��cx������R�{��'$�aR���OG:�ŏ���7J)��m;�/�#0"@��s���}D�CX0g:��`���\L �����-l��E�Z5n��x≧��Hrd҅^����Ghk? ���7o�*��ؿ���2��'�����v�!������%K9����q�W��^72`�����K�w�	���݅s�clv/>�����DU��c��p���_z�{.���K�ٰ�������L�d���bӿq����a^,r������5��JB��$�M�6I���Q��\���K_���6+��8�e�������+?�F�@֬.Cj��&֭�=�'tf:n�K�&�3�t��Q����s�C��UMt(�ur9��i�{���q���\.�;���v��;�wo�u����̺��=�Eve���P��bAXf/.��Ta�rn�6��Kf��������y��>�k��0;��>z�p��r;���E\o�`�Z)`&��@�d9����M��$��OǱЩ�L���%BvyY�	�/�h��ٙ�Z�p���l���G��PC5F1a6���҇qX+�k�������g��C�gϜ��X\�����Q��S��]�"��ʠ���!�ٳG~V:�[�6TM�B�f�I�R��}�eKh�V�ģ��I+>�b9�l:��o�ǻon��.�m;w!���N�)>�aQ_�G{�9�t��/7,-(v�����D�t�̚�)-�8��C���G=���A��lt��MY�0��r��v�<�w �O��U�F���� R�o�VA�V:�jFUgx�V�ӫ��1F7$�`#0����gbh��@՚�۾j�����h6>��́�wtC���	��e�����hG��E%�w2�w9���ŀ���N�A~�s��ǂ��'W54<,A�k� ���5m��O��?��i.G�sqޠf�~�ۥ��q2ʦ�Z +�WƆ'F���Y���j&�m\����5��yʹ[���N�}��a�ǇX��b㛖�.���)к� �/�^�tx'�#���H'a�Ѱ��b��L��Ӊ��.dq�=����\"���>�SX�h\N����0�
��6GF��8E��Ⱥ��8���z�i��-EKt�'W���g��֭}_���l���U�5RU+Z'��#�1ع�C�6h�AV]���9�;v�&B�H	G���	ry����2��ߕٍ/<�*�~�Yi�PF�^�x�'q��.G_�$y
/���LI�5kvm߁��f�>�0��`����"!l�(�*�*4��"��Y�/���t����V�No5��!����se�U8�̳�̳/�pc�i��&����3O#���O�݋t<��\�Klߺ=�]"� 1�u@ �A����G�}��,T��>dff�,LZC}� Y���sS�l$\{�}Z�6I�
�̈́ac��1�C%��;��V���ɦf�%6^gI�A�~���hm�����ԩ����k}�iT��2�xRnj���!��&� �����~_ t����b��Í���/�)c�^�T�<���<��&���*6Tr�9�(�K������/��+I8�c8�@>+��?A��.����_*vS�=[[�):�>6j8�t~�R�����3e����Œc�a����,C�W�C��e ͱFԻ[���L�\�f�h���/� �����_M����t\uJV�l0ї��2�7�0f٢/�vy7F��K�������Y \%�ks#1EtdTn�`  硶�
�������N�m��1R�B4�f_-.<�K�Q�,�h�F���;�������.�pg79G͢��$���`	#I��E���,���W^�}�>�-۷��e��vN��I�9k�t[���k��{�U)+��$��&��P��M����m�� �|��L̊TԻ����;�gy��W)j�d��oh�j&��0�:X�jތUg��O�5�?a�h)�E����㥱�_|ބ[�D�����h\�'����h�J)ro{��y2a|>A����܅s�e?�c��G����J�iR��#���10��Cvs�����jٴB��<��'>���.�%�=Y2/e ��9����ɀh�;%�p긆9�/#��ev����۷o7���gIR�&��'PP%H5k��&��fQ���9S�Y��R�2��e�Nr�<���mV�i? �� ʩQ��?�+����H��<U�)�6��j����J��n@ ��I~V~�p$�M／_����x��9���n����^wֿ����K1k�Y�&h��]�����j�5
��A���j�sOF�c�����Nl��>Z��U:4ꮮ����G_�0vl�-�0����?���2���ڌ��.I(y=i�}�6,_�g�y:�A�߳C�QW�Ӗ6�Vɳ;d��d|f�\���K�����4L�C>�[��#q�Ϯ8�p�[�&V�<�t[6��Ay�̪C������S�=�g�z	�����r���vD��r�Hw��[Yfˬc53rt���ϭ1�&�d�X\�W�Oˎc�[�����%�s�>K4a�N�M�v62�iӲ՜f��ۺQH�$�P�2�dvK���xd��q�-�����������df�4X��x��:}�fL��ɱN'��׌L���j�s��-�e��"���o�Oa�J���?�y��O�t�#Ҹ�ĒR��r�T|/��ه�/>������a���C�P��@�X��s��N��3�@��Ef\�ҡE�T�%�eH�B������mTݫ@i8��sJ2d��.n����L��E�C��H�}�Z\�<�Ti�^m�*�P�P�	#��!�T��TL@\�%�b�J=�!��l��� L9G�1]ݽ��g�)��b	�b��n�/r�ѽ����[����� D;�p@@`�`�P��t�lU�<9��4bɬ����bth�d�r���71��-#h���O�����I��'�y(&�Y/�'/��wѶ���d�rf0�Ll�'��9�K�d��N;��H���a �|c~��u ��m�J��������byE�+0@&L�M L�]BPHͫ�Y���.O�uz�	�R���(�g�q����Ʀ;��y�_��r��!��L�>���UGF��L� 6c�1CY�|	�Κ���v⢋.�}��+���o������͊T&+��n��[��H�woB���c�0��@kv�V��Wt�,CRH��8n�,��}^V\c|P�C�U]UcL*`Gj	˖/m��ݻ��yo��p)o*P�͞��12�|�>xMX�ך>}��|5r¬U�[����� Ly�H6�%�ي:׉|Vtu�:{D�p[����)P�#S� �+���.�O<�/<�g�U�aU�hlhAWO�$=}���G�1�}c=���:I��N�����p�-7"��������0Z[[P]Qe�lA���%ص��Cc�d2%�w�"��q�z~�^���s��W^xooz%��Q�Z�?K�3��F:�٘����)Z?�OZ�\vٿ��U+�c�,Y�>�����f��%�]�_>�,�qtv|���6�V�d
�0+S睱��_�<3�
F�,X~*����Ӹ���op-S����� E&��<H%X�tK_�j.�؃���ګ�[o�	�����������Z�9�W�"u��87ӥ�%�6�2^J�I��؀����rm�ɉ�[|p� 5a�S��f�\�Y���0���
�Q�Lm�֞��蘢��G��`��F韏c�.mjL��J�(��o��?'��'��{�O�W�n8��b���},ZF��L�H �wy=�9�ޛ,���Ox�S@?�U�u��p���uˑef��(��N,��'�?��L�T���p[J�����_t;��m?<5S�**Gz�C_���&���Fn���B���yT��Z�鈪�ޠ�5�A�Tٜ��I;w�� ���M�'gE�Yg!/���_�*&�}����A]�=A�Z�AX�iV�0.@o�S�0a\Xd�da�UɃKD�@����:��(��0�݇��.ģ1Ѹ�>a��~]WQ n`@�Q>�Gۮ���ҘR��
�ߍ%�Ȑ�\*��ǋy3�⧗_���>�\n�#h�Z jo�ϟ/bc�)�-�[������6z��h��Ī�ܬ�	#p�f-����I���>ځ�L���'-�����Jώ�Ե�"&��ƈ!n�b�í��A�)m�;�%�̘g��D�A���k?9-F�;Ә"�2	�
�
���H��*٘�-�s�@�Nì�M'�x@F|6Mx�c&a^�9�x��Y���p�=���/�L�.ت*�\��8�3�66Kǯ%Gf�К�k�1r�������؀�d��9��ߋ�0R�-hjl0�䀿�y%#{"e�	��4
�Ff���u�u���Ϗ��[Z�+�E�E�G��ן��ߖ122ވ�o�2@���&�dLoԘ*�`~v��T(�͏�1�E�mp}�ư}�f�4 �8�}�X�|1�>�ۆ'�|S�f �.� �h�s1��ԡX��M�\^J�<�D:%�=���m�.-��o��ױt�B�؋7ֽ&��~ޯVU�%��hTٕ �n�n�����=>@XE
��Ξ��>
�{�I�����_¼ys���O�_�ut�߳�CtGGH&��,�Z}�[��W����qtuw�s�M7�g`|Y}��ػg/X��]�,;͓�����
���e�9���_�J��d+�+!�)c鑟D<e������{#cjL��Lj�����y�<�6�	�B��<�}�R\����٧&1���X2���6ʐ�;2�L���}4�:"�R�Py�V*����2������g�}���3	���1�M���c��,-�dV�az��:�C�3j4c��7��R�&"��Sω��U�Nd���l2�4�vKW.���c�tR+�#.�kNv���?��$�r�9��8����{o�X���>�i��k^��i^�/[QɧQ���l���9^xR���g���C�������4�zd��	��p�l�!WR�Z_l�� L�ᚄf ���rS�����,w���G@:���&3Y����mޅ-)��M���*��8��[DMAo�r����yű�c��4`4Mˑ�TL�6�A�KG&L@�[����1�J$����!!	BNJci��!=�������:m�C	�s*�W뾞>��� �Zߌ|"G�{�*�w*����Y3��\Z�i�Z��e�қo��ؙ����54c�<����_����t��
<�,ղC��Z����l3�SL��	81��r�������?a���!�Kw��n���K5~М��#�V�`:(j�%Cx�ńy��:�٠tI��n���	]߃�������M{���"����� �lY��?�A��`�&&D��A�zS�0� ,����B�*"@F��C!|�3����#��/��2����
�Dp�$q`4:&]�d�fN����>Dh�a���4f(�S�RP�I�k��n�Ɠ46�#�{�X�c��E@�I+@J
�=>�i/!�Ԡ��Nm�Ip
�Z���'��0�If_a�*�    IDAT��׋Xa�U�K�]��������:ka�|B�����D�^ضH���	n�H�����c1$3	�DpVr9K����Q�D�O�U�b=14���w�Rq#D�S��ˇ5bv���x�USS-&�ܨ����� L��[�{�MG�L��<ҕ�,�JT\�2~���uع�
�CU�~N��:a5����'���p���`����Y�{�.�{����%�B۾N<����"�<�+�"�jn��&̜9�Tm�q͵�W1-���!��,]!@(:2�dl}]{�v�w�Α*95��q������?�D*��h���G����4�y�M�x����0k�L��bs㤓>�{��3�������I,\1�]����㇗]�����.��rd�C��넇מI�W&��2B���ސ��Y��%U��:���W�Iza����;����W	��x��j6�|��a$�a-5����v`Oi���U�ks�0'��ߛA�9�h�K�!s���L<��G�k�y&=��Z
b~.�K37�	����@�N��,�F�>�]N�窏'[��{�fK�qe�dE9G7�1�փ��p�]x&j�xY���RL�_X����]enPe��)�ˋ#-��6~}%�2�3�LC 6@ɿHe�M�
��YA��-n7|������{?�{i:SD���(��|vG��l����(a��8;r8>zPwd���d5���8�[�M�%(K9�R("5<"��`i��ƠӃ�P�����bw��u
B��B�Ǣ�(
(f�H�f1�=��X>��S��ؠ2|N7�jho�G>G)�Ă�3��CCh��A������&�s��ϭ����3�L�t����ž�va�X���b$:&�/ļyDKDp��[�2��"��"�����QJF9��#�Y0ޘ���8r�7ngg��q������9	�Ę�c�u��j�3��[`)��ܸ٧f:X�!Z�Q�����G)��(\���<n����:^:�Aq23�%�ɜ�	���*d2�;2��R$���<���\��}�3X�p�t>���xw�f�L�a�C����TAU(��3f`���ۍF�� �L�����S^I9��@�|��%E2i0��<�sHwd�(�/7'r�+�lȿ�9�ڷJʘ��0��6�JƌCS=��)��u����:��k�P�)g��8�V���2�Qe#Q�,�*2p�tR�?'V�1D�b��MEQ�!� ��!���|m��׀��1EytD T�\�L��D�`������ǁ�dM�"Ǹ��h�l�ذa=j�Cx](�"��<M��),����.[�/��
������B�Ĺ�^Ccd�O~�8��%�����{�6|��p��w��u
�9�)�����ǟ��/��a���sϽ�Y�f��n_/	�#g͚���W 2A�qǭ��ob�̹8j��H`���=�PW�Fھ�Q��2G�!fDm�/5a�%��G��XΎ'��:n��n��v��ɓq衇a͚5h۷�h�4ˑ^��%�̨C"9�K��5|��/�����[o�A@X(D�<5
K���A��cr��XiI�T��˽�t2�P�54WenՍ�&$�Ճ�Eh��E���1s�?����ThU��1�]zT��9��5�a	��Md���Z�J�$�6�x�~�]�ړ�ϟ�E��9�i�4�SRW$Ȋ���a�>^�O�]�ПS�G6����?� ��Y��O�~K�]�2[�����j�p�!,��'��}�LT��������@��<8���s�$��ʌUke(Eo8��>B#e�=��#�,MJ����e!�D�25�6+�*��r�?�(=�ʤ���zB��M`_<���1�H�'��B�eD�s�R.�A%�g�H�8��qvd���s��H������L����wJK�c6���$�@䅹��`ϕ0�ً���èi�G�V�"!d2)U����s��c��� �p[��1X{��9=b����_���~tuc�s?�n7.��|tv���ys�o�C�����6C���("�OJ7�* ����]���.)��.#�`���WE��7 Z;�A�S4m7488HSe���� �L�f+x�y\dFv��.A��A�������N��+1�]�, �ZZ��gᆮ����|�M
�y���%��&A!� 7|��=߇ݑ<N]���dRe��r��lvrw�d���Lm쎤S��#�|"��M�s8p�Eː�˖cÆ�8��O�Aݔ)��,�,���9��d���,��fs�	Xэ
 �-_M]_bYb�����E3Ա�Mu>�lhjjQ�;�`dOx���gdeɰ����x�$�@O6eJ�\7��EF�N��`�������[���L�����c��d3��R	�R%��Ӧދf�Y�3���Ȅ�@��TT�Sj�H�Fac\��Iv#�4Max�6~8�~d�x�A�����Q.іr/��}��+X!E��6��T� �}Y�<O>/�]T$Y�6u���1��翊66�0M���v�q����'���x��5Xuءr��޲̴r�Jtwu�`sf�G<��ٍ,K�����bѢyr���1�6����>u���� ���0�=�HT
y��J�u[�N�n+�/W��(ǹ�6)�ĊX�b5��F<����Ϗ����W�m AY���1X-.T�8\V����:�	_��8|�!x���q�UW�($����<�k��5�1�bP2CW{�G\Ϭ�Ý���������3���[�|9��bhk۫: ��4@�Ӄ�O?] �t� LO �gP �)l�صPO��a����m�l����CM��JF���{�^�����x�|A�".��D\�r/�$SR�)�e�ۚhTCȯ"��&(6���X��4J/��jj�աHz���o|�q�{Ƒ��!��y����k�ɪR����.������?��Oӄ�����Z|-+
+r�Q��i�؇j�.:���v"3Љj��t+�N��/uv�h�����!�ר�����*�L����8�\"cBh��.1�)F�Zg-%0C�(����Aj�
�j���-]���}(�y=Ɓ�t4�O.>]A��v�Y�;��a�����>a,K���hvx����Y�\pR�.�A�;|��l`��͍T���4�T��أQt�E�U)P��a��Ձz�Syil�������5��=�p��?G>�����y'����#�7�a��9bM���T�@W�2�X8����Ó�bQ1d���?Ⱨ�Ď];1m�L	2�.ļ9�1m�t�_����={�m-���y��b9�hi��{ܻF�f��EÇ���m� o-��W�g�N�4���.S��0��f����2��z#�*�_�s�M�Zs9�����r:�����5� ��X�����(s��D������d��N������>cr���dVQ[8�����u�	1�jٕv�o�.E>�������7_$gȏ��)ZG�;ѩ����|A�x��a�u�k��8�Hg�<�`������1c\n'�ly�(?(o%q�=��pTYX^�Y����5�yb1� M]�`�	���P�^mbи��<.�������ߋ��!��5T%h�l�@�j�`*�N<��%��/��ٴk7�G�ʏ�*/J��L.˜�PDuM�H$|��Jp�ع����U��V�(�x�j�<�`<nz�U�bdJ�/~�}�B����فb!�l:�T͙�~�e���fpp�\�?�0���h���SjS�.��"N��j\���_��}g��Ni�:�Ӎ�o�=��SO����Ck��P#cI��6������E_��� 뇋ɫ��1)C�Յ��E�N��1���F�����P��U�<��c����e��h#��:����r7��*�f�����p�i���I��؈��)j����կ��C]�%�ȵ���kq���{��%{;�{�4��ż�7&��.lN��/���ب�Kv<�L�J	���:��d����O�<�Ē|^��
#��-&�F�7c�rδe��f2�Ҩ�0��9�wx^��##"9�5A��JN'�kj�y���M�����a�9���m���g�01��x0��/w�Y�����������Q�?�\^l�H0p���e�h�2gjK�$��A=}�p9\�TWaldTz��	U����l�p�[�idp{=��i3�=g�?� 슿�q����|k�ۼ4/���c��b�7-oq�Y�':��^lE$ǆ`�זף\�9G�ėDU� #��d�f0� �E %��̏�\�sF	����(������2�L<����m�b_x�k �C(h���y-��\��e���8�,U�yn����
��s[��)~ޤ�������ő��T��Cf�(I�LILZ�+|e?�u$�B:�)��a�YHXKHes�?00��h�L�Ձ��R��i�t�6V-X�}�d���\u|6'Z���ֆ�����1�9��ї(/z._�C�sę�ã#r�����x��װs��Z�x�hs8��:��Us�Q� 3|��5�ͨu[;�A3�b6ο*c��]��I�D�lݞ����(=�Y�2�Yk�7Xa�
����e3�7=��#?��̈́i!7AϗD����|_U�,��8��N�q�w�E��.�kЩ�CͰ���)�C_g貴&L9�^��s?b�\^��Zh=¬���ǯ~�+Dc�b�ʌ����?ގko��r��:T聗S>S,%Ξ2�RN2��c��������i���VV���*	��K���iǶm[���F�H�0��U�D�2���uu5�)���M�睬�h��~�	�ɹՌ��^�w���5��i�#�6A׌ү18ȫ�9�-���y[��$e,\�\̜_X���0�^��r��rZ��&��
�N/rE���Q)�a�xņ�nq�Hz�(Y
9��;el�_��x���R���m��ޮN񻪮ᨣ����\s�5�y9��I��{	/�}�W���^՘���U+1��
�^�U�v�ux�٧p��7��o��e�p�y����_Ă����O�'���_��X
^_X���s���G����f��,�)�TȠ����}H�ȥ��b�>�m6�TQ,������1�^d��X�B����Vtt����X<�?$6:�:�+V,öm�PSW�c�>^4UUU!p����Q�R�M7\�5��x��RP^U��}cv0u�ҽ���²e�Dx���9sg���K�.���V�d��tRʀL*��5�Ub���Z*��]$�H�J��T�9�R�}Ƶ��͝=W*�fz������_x�y=�.��1J7�0����s&.�u�|.(�#�/�\r���cU���Q@��	Yk&A|������_RMm�L[*��%ag,P3(����&11�BV�9 ������\�l��=��~�����Oc�~��G?��������BN{�� "�<f4{�L/Ϭ�e��2�8l���Q�gd!SS�L�\T:�&�����u���NM0t�W�)R�+$K�"�w����e�,��+�p$�\�����]F[x�{P@A�i��W�t��a6�{��#T�#�&���	�d�,E���f�jmnm��C.��;w��?�V���Kʊm�l�m4��ˍ��M�nm@�����d��u ����F��C}M-"�*�~7oz�x
�� �͚�ۯ����t�͵k��'q�1��{�|���`�F:���^nn1>�����{�(ɪ2[|ߘ���y�ʬy�b.e�[[��}���q�v�6�FA�D}j;<�F@���������ʚ+�1"2c�{c���w�Ɍ�W������U+�Ȉ7�=�;��o����چ�~~��Fbf�]8��%�	��wX�eC�A �\Q���](
�Oq�Yd�4�РD���5�~%��M���#A��K��'0��CkȖ�5�ȽЬ���^Y��:^Q����8�ݪT��J���5����?�^���k�Sa6�"i=���n|�Ϭg����&[s L��g��%=�y<|)V|<� �����dIM'0ĠY�`QO/v�܅�mn��!��ҚK�tV���U�J+��L��_�Aܾ�L��~�hƉ��i4�T*!�s�X������y��Uk"�6>6e�|���o*�Zd�#ã�qqḤ��8ǒ�^�g��g�����:����\8������G�|�X��"�j���V1�����J�%{�A�0�x��5�����-iK{�d�>4�v�����u{C
�9����������U)���hnj���+�o@)�C��#Ȧg0����cT.�l�MS��/�o~�(���]���-�1����된���m�{�z�{��x�7J%$��t&���V���/��b�L� ~$SY�]s:�����+�7�Aa�Z�uG� �2����fQ
�
�"?R�	��1��gӸ������g�:��E
�* �W���x7֞�k�o��F��It�'N����ĸ0��\��!�!��(UL8��u���G�H6|�d�8B�	{���"V���,��5kd74F�a�za�؀�㷧�G�"�EnPs(�0Z0��Ky'b�����%��s9����c�oZ�p3�k��8^5��c��ս*�T���j>U8���:��w���U�=��%�Z�l��eft�^�$��xԈi�9�����$�d�T�!�2S�Q����;uݪ=Seɲ����7���YT|�gO^���^��h[��u�QD՚B�_ª�q��Ch�԰q�R,�nƒ��p;���i9�vJy�6��z���L���5�zVƐ�g0yHz��h�h�ʼwM4\�Z��(��ȥ'��ٕN'��
�0�|�q�``�Ȕ�0rornLnJ�� ,��~lj&��I2a�����1y�̩�ܰX��LI�nl����n&SIA�4�%�88���p���T��{if��T*�&3��>��iol=5r�\v�Gq:�oK;�3�$^{�e���Z�q���Ǳ}}��lmk��öI2A�NY�;�TR�66�%K���6㦯~EL>.���4mj��= gK{� �`th�Ph6M�A��f����c���R/�:T�	<�,?�x���f�89���=mЪAU��KMɄ)!�W}���]���N�U�d�r�؋ E�v/J����k���лJ�'Q��,[���j�WF瀫K���(�
�Y�l���q�{Ⱥ���#�026��% �����lF��X<&�`��o����A��FcW;��\$:����]%��g���t�|&�@�mYp�ƅ��8�;g.Z�nmk�Ν;���'�;�/ٰ��qIE�!g�;S��Bn�J�m�tړ�q� ���;��+d�t�����k_9��~�I��r\�Ō��\Zu�����.�~oP4�cS	D�Q�<�K��b.�ޮ����-g��|����x��gѳx%j���xm�^ٴ�r�j�E�� �1���t�$���fi�����ރ�I<�ģR���IE#��n��z�Z�M͍p������l�Qsz0�Ja��5�
��/\��υ��[7o����/��?��8v��j	�o"��) ��7���bP��_��}�X弜+�@�H���9Ew�Mj��R1�t����O�S<�����)�B���z;[e��>x�_���cM�������+�K&��t���qd3JSy{4��C	���mx�G��e�!jZe���^fij�g��MC� ���a�d�-[*��m�>Z�����舀.v���nj���Ĕ�K��Hc����'A�?献�`��iL�-��*�,�z�S�?������t�y��v|^oNԦ\	�E�
��4�}t��k�N�ylW��\��]��8��1UW�0e�~���<W^�H$���Z;�"��M��&�~_9o�����ο5C��Mx�)LX�Vs��Ϟ����_��䎯ʲj̜����I�}��2��y�����z�B=3�+��43�Z�!�>�c���K���6B��^���\]]Q    IDATbC�ži�ǋ���:�U�1*������ ��|6J-�dт"��3��q��p������,� e:R2+v:��w>?�5/�����8��	�XW�i
5
�Đ�T"৷� >pVD]A~e7�D��8��Q,]�)����H�%118W (@���U�?�tj�G�QH� Ps"��"�	�*�%�p����n@!�������[��JH�:��n"c�rx�σ�7o�7�u��"�~��k�2�p��}΁���ꙹ�, \<�����@7B�	eW�͟7�iK�T��K���+Ɲ�Wk_,�>���Ս_�U��5�C��&���`��ǅ�;I�W�!)��I48T�e���AT/��4W=�����\���4��x�B-n�y�-j9�G�p��{GU��n�JUȓM�w�J%�l����cC�,a��g���FDkE�yO[7��*���z*M��$�i����|h�g�f���}^P7�$��<��fS�����S
XQn@Q3ӑ�/z��m�x�x)��`��E��^�n�n6��R5#�7w|i�!�	�� ��a|j\,u|A�(PL�q��DZD����$���".xa���m���f������`Ǯ���w�gQ2�a`�	��+]((��w�قg ,N4j��,_�w�yF����Q<���ذ~��m~���Va��hl����>�U��6o{.oP�<�z�q�7�.�v�<�8n���L ��O�t~�a�v0+���D$��Ȥ���]����(�9��e|�P���;R��"Bf]�	�>@��Tf�X(���&~�㟠�^�	L�](��r�pb��5���D��#�dW+X���RM뒩f�Tȉ�t��9��Js�|�����*}u9gs�b;m`$TT��P���oVd�����]��&ӊ�H�17<�����gҜ��l,�D���&��,���8$8��8��� �c����0��n�6b�m�Y[�S�))l��i�}��x&3�<�w�sV��C4f�QU������\�~��t�>�:�c`�{0��T����D�W�~�/[�#G���R�����z�F�x�W^�I�*ߛ�x�@��?��_<��=���+3�"J�)Ă@&y�n\�|vNg���4�Ŭ��Tk�#��U�$�L�ҍ��*Cf�i7}���o�Ik!2Meq=wx��_@w�*��w^p&�X��#��߃R�D����5?n���7+{�0lq.A� �7 a,.�&���GGa��"c��=���l
�%���K-��8t��먑�e�i9u�qx�T3h�֫���.G��`|l�DCǇ�pyD,���7�Ы$IL��!�����D9���p�=MIs�]�����4�/�E9[@�*sy�S��B��ѣ2Q{/��َ#'��O?��6m���������,���Ěޥ��-8H��i����?���$ VdNf����&+U��3٩&ّ��4@ҋ����w�&'+�\+�ָ��0���N>M��]�>�fXd4��SZ\�������U�A��V��_O�<�Ne����e�̙t��B?�	� �#c�����js@��ě�������vV�REA~ӂN�.���q��x���M�U���U"�ć�ɠ÷7��`5�$.����XeG�kM�vm�+2����eB>�I+�q
�y��M��t\|}Z>Sy')�S_ǀ_�����tW�.P�/�����ŃsA����Zq���L��DbB
l��ݱ��+��[�8�����S����b��v¡ �'�x�9V�o����۞\�|¨���V�\�ˣ�}�����&��3������[���G�����K�:>���ؿ�O���\�f��kz&�H4��/����~���?��;w������������Cx��-����.��bi"�uc,&i�/<���v��{Pl hUA��7|���_��s��rc�F�4��	��T
��ѡ�Gg[�h�
�&��D����s�.���̴*���ʧ�!${n,�zz��_>����9�݋�#X�l�lK�<���{imRF ���d�?�2��|��w���E#j*���H>֮^�L��J���Tb���X�t���^rх����}� ��<�4��MU2ን�!+* �����^�����d�� �\��$3��Ci���P-�T���I-2gd��G���x��\��Km���)�G�E ��EO��Hp�3z�zr�Eƌ�� �b�)���$d#	�0�V34��t������w�>_�𛀿��&|r�Vs~��/���6�j[�"[,�Z�Fs̍��8��e�GQEpQ(�P�(D4�Kg��j�
����Sa�>!�&;`�N��;�u����%c���
����PEE\��w�ӗ�(%ᨙ�e�0,!��Kw~O@���0aa�pԁ0j��3a��/���Ըl�RŜj�D��y��N~/�E(̧���=.͢�EΪβa�G^ۋZ2��p��&a�bN�B9��ȱ!)k_�x�z�Q��Z�"U��|e)��^�\E�XBblB��LP�@g����l����ֺ;�p�-Eȴ�2i4�6��v`xr\�y~�Q���(���P0t��������=�[U;&á�G�TH�G�Բ��N= �)��td�p'c�a[.�\�5�uVZ�ϱ����9�����,uf@�ϋ(��V���N�����uѧh�p���:�)-"+��D?����9�ﯟ�O]&�Y!��;�`F������I�\F"9%� p*L6�ぞ_Q��Y0�EaL� �Si�#!T�.@��/A(B�������-*��j�����퇔�
��k��0�@�>Vq)����Cp�q��M��LNh�LeU �kCtd<�,�6��)��lǆ�!a/�'�C|�?��,H�0(�7K]���$������{�����	�:$�g�)�) ��6p��AlCV����g�ލW^~�<�2������e���Q5��8P*V�DU;62���x��cJ�B$րg�{	7��E��*"/�/Z�;�y+J�4���)1��3�,�ƌx+�J���֮Y��N?�>��z�%Rm�ʎ�d�G�������}�<��r�F��da������ؿ��I�.ѳu�/�����>��O�O|N�oLY���>DZ�wh �dF��ǆQ+[�}�f��\Q�^*J �oL�Q>�k��ҟ� �����H��4o.�GO�df��e�p�x�*��!�b��K�v	���q��碫�n���W���o���c���Y��Q8�z��4ӛ�<��n�U��s~[ظq#&�&�'7Kz	7�XʦB�8������������_ujJZqsL�h�{j&�u���&p����ƪ�<�r�"[#�T#�
��q�l���8gl�zͼivXO�ߞ���r���g7F|�Y���4S�������t��+e���P���7�ɶ,�h8��/[�{�a���x�j5��x��}�{i[�+��;,�7�19t��/@��@i$2c���EERE�L���T(Ѿ��h���M#�+��Vө4\n��LQt�}7��pr���'�`�<{0.�k5�2B�>��w�KQ͍!覠�&��w�Q�F��o���a��� ,�M�a�=�O�`���ʥ���L�4o�����Sr\8�� �
f�ܖ���v�c���H��V���B��#0'2�3��e��p�B��&���B�HM��Ɏ/��� ��I� ��K:izx�L��qD�Ƣ�^���tؿ_EN��Ǐ�kQ�b��%�EB812�pS�0~�XE�5�*N�j.&����6�
u5�:+�_V7BV0$Ȕ���e�-{�B;��T@�o���ɉ�EU���S�%�,&�JL����wiA�_��ږi�DR��Q�0��:(i�Ŝ�B�0�G�v����v��z`RϬՃ0����J�bul�uJVm�Q�Ie��RZ6��V���C�w�L�g�b�_�=Ѿ��m~�jE[+E�=͝�Au�P���.�,zL��z�R9
�2��~\Ȩc����� ��ܹsV�B��YO�����������������u<���� ,�Q��Y=�EKkyOy��p��#SJ�B��n�D�#���B�bn(X�hUU;2ѭ���s�����C��
������w7��N�;2�{��!^ٱ�KW�Ou^�pLD.L��2f�<�pu��3���]��-߂����;(�1�ǽwݎ���F�ȡ>ajhGp��!1	Mgs�76�ΝƆ&�XA��a`lL�
�ۚ%x^{!�[�{����ȝ]�^5�XTlP�6=�n��߂� |�Yg�ڿ� ���b̤E�ؽg7����x˹ê�Ef��܄L:����d ���".�^2/LK��+�T�q4ߴ��n�GĚ���008*���\A�������RZ5�ްg�}���?���=�Νw�{��.�v*�L��G[<^6K��.�u��thko�j˖M2�9&y������jQh�9�X±(��u�W���������}����,W�TT�����Fβ;�06��N�c%�'��iN-��Y]̢�Gx�x�L�&�5��jzVW���gq�h�����1�A+�IK>���t�Pl�!���s�Ź�����<����1<b�6ӕJŬ��h(��0��o��1a�k5���_��{<~W-ܾ�BϤ�$�Fd�~���$��$��
����&\]35Dl��8���'�*x������U��Ơb�&�R�w��fK"�Ρ	�n3����'>x%�8w���R������m7��+��[@؞���#�� &UI�P����	��"�o�nECG�0`�C=�����d�LVk��2!.�BjGTq���a�<U7B��^ٍJ*�x4_<��g��X&!��w��chin�����pl��H@��Q0ͅ����C�S��`�H�).;��B{Vafp+�,�o=WXŇzH�:?����ǿ�)�4��{�������?+Q��rJu'@��,��)��5�*q�^��B7Uh!7Rn�m�)6�H�kG��f�t�O�M�`Mj�y����S���&����g!��1$8���f���^�Ō�V��;2�t�лR��y0���|o=�Y8~F}jL�U%�,3�є���Te}������rufA�x�iZ�����>��:=�ړ	#�J��/�\:(طO�?���i��l�DU�+�<n�6u�K�J
P�j�T�å��|Ĳþ�j�l>��k�N�j�nţ�+�eJ '#@�K���^7�������+#�����y��b�?�n\�y��8&t���~ժUr�}}}"��,���F������Ʉ�DR�*�<v���5m'����tb�JK:#��+_ĭ_�g�C1|��?��Ds�/*pI��;f2��(��H��6&�?<�	w��W��h�K���4p���3.���1��l
l�#�=L�ʵ�;N���~Y($@�I��C�\��%K�w{���Ɖ>Qwө&�&ѱ`!�|b3����`ͪ3���ڮk�}?�~��*tM��G~�����?��E+1<D{��=�����f6�'3���Ї���p�]�ٛ#/�.f2Yt�,B�4a�}X�r����<���"��kH����	�_��ؓ����w���ށ��{l}~��m�9��f�cU�I,�R�U]�n^;�<��a��ԩn�Zp̹γ(�׊�q�+�8��WH�2f�<'�NLo
u���>�����A �s��:�_���S��1���?�����T2^���T���������w�5�X����Y�{ܘ5�<շ��{�Mф��<�<�����Гw:�ΔL���4��Ww�gX�8	x,X�J� }�HQ ,����t����R�{��l�t��s"ׯ�_1zeK.,�g�U�J�|�CW�ҳV�������E��ad��p�=��ґ�Ց�	�;����m�w�
����#�`,�#۬�l��h�LO�4>�&A���@X�+�PKѨN��g��h:Ii	�����8ڛ;m��cq'F�c���]&�F�lZX/2�".����Ra��4���<s�i���hX����o1S�aǁݨ����'ư`Q/�Z��B��p+.�KU8�-��ea��U��=�T��Ձ0^�7�21��J��R��뙰9`��}�O� �4��k�(�c �}�Te%��)4��)D=�5��A\��Y"���|/�[�V� xd�.`��9�L��(=�u����$�����ܺVEu@Nk���헴�˫0z������뮓���]����O~�Ǟ}
��V�XEb�1 Ë��8�(K�7a�o�50�s��΅P��Y6{�,"(�V�
�FD����KY�8e�O�ۢ�:3ME���e�vKҝͲ��o�%���䘘��(������1-����?�{Gv���y�ф�}i��6jD;\dy��^?
��F�D��b^දބ���5t����7|^�6�u�OX����
�fR�ق��/��M��F�����w~���#�f�tU3��|�������}��ɱ�69�q�+ ��Kcf!�v&or�蔔pY�˨U,�8~�d�;%>7�e#�1Hf�iB^�@$�����m�v��Y���0�o?�aIG�:r||T��.����]Hg��+���AT��餺N�����u���KW��λ@��Ͽ�/(=]� r%��f�La:_��U��w����	p��c���J�eI�I��K�q	��݁�����ϯ~>���q��!�t�y,��J��j��H���F����\�^��i��׼>&�u��Y_�ns���KZ�����c!?G3�^�_��,����|^tm�����Uy<~k5���|�S|=u̚��c�0�c�1���5��|ԃ���_\�{�Բ�z2��~�14���S��a��z�O~��Ng�����UɢfN#�/a�F�i���F�E��`Eo0�j���0�YM�,b������E��,�@��/G𜲼��*���U���p��^ ?g����
#p?r����n��'1a������J%�΅툴6b"3-�����NЄ��C{2xL��) 0�nH�i�����d���𔝈���Wwkd���0���#3	����	t�tI�{ײn=��Q��{��?�ż�?'�Lp��SoS*�.-jx��)�h+;b��܍7��Ge�~���Ń��8б�m�e!f���A�	�0ߨ�,;(���)�[��[v�a=�Nas�!���QA��{kWǼSiêb�����¦���w�:��Ì�w��0�*�	��-
�Ӂ�]�����m�&�|���[uoB�dj���Ȅ����i�t��N������#B}*٤���& ���׀i���=_��%m�qyP��b���~�#����a*�E�QE��4�4q!빢�AV�Uh1�3Nk��"D�C�"V���L���ж�N�\oF�Gj8U)��������b�@v��#�4.:��+MJ�0���?2���.L����C���	KWG��`�4�0֪���/�J�:�^�V^@X!�B�UFSЅ;o�7|��E���?'a-��dq��'�	n��Y�)[���Z�:�|�Zlٶ7��m�U2�ܨ���ុ���/;[ ����Ii�F� �+UUe�Z�+hjh��N>�˰TU��`P�S&�ƞ����tho��2�8!��֬Y��{�a�i����
�\����k�?+r��_�§Q,e0��@�s�^х��Ϸᩧ������V)��<����3�)�nI{3*U��)K������8`�܈�-@�4���Q��c/��ObÆ�16J/�Q>L�/'���ݳ�=����k�� >|��[�*Z:Z�rY��A��VTe�քrC��J]Qm���zT=�D/fi������D���	���^��K�'�w�J���lQ	��?����n��@I��Gn��Tk��O�0}�zV���Fl�ɱ`���    IDAT��c��5�N��tV��5���:���]�;�g~��m6'�������y �[.���|�l[E!i�j���zY+��9�Q��`����35�]�_���UUv[�s��%�:8�Iy����Ԍ�2]���SU J� 
�a����v5�$|n����t��߾'l&L�#5�OG�m0C�|�i�V����@cg��0j��'F�J��:�b9��^�����U�&�����*"}�D�0م0A���0R9q�İ��U����5��8Cb)Ao���V�妐u��s[�1�\���Su`@!UHW�b
3�+U�<�o���X3��;��>���.9v��w^z�58�~a��b-M"ȟɤeѦ���0 +T��T�ؾ�K��Z���J5�Ac�W���$v�DR a[@�Oz�_�f�	��0G�����iA�&i������6c������N!�
Gm����g�(Q^{ש�}�NP�`89�fSq�HG�3�z�z�]�
x��&�h͝^x,�g���w�#U�H�;�v�T�5��8=���V��w~p{:eM����UC��`yK�4�����Zt���t��l�nj��"����(���XbH7%J�=7)��bG��*�7}~�/��ל����]�Tj �E��մL5�u�&�~T�\y-�S�� /@п��6�(T�<�fU* �cc/�b��c���%��� �y�Wp�m�"�������hn[���~�j�M ?��*��t��ak� ��{���q��?C����n��-��ƿ|���AӋ ���,	2A.D�1�0&�,l���@=����O��Ã���N�~�<��R����3O=-�1�`��5x��mx��X�d���*:;�1><�����q㍟D�Ɩ5�����~<���� �gq�����%�x걇��Ccԇj)��	��Ma![�!)j�)a�؇8�@�����w��^91 �c:�E�J�U:�-�B(Z%,[Յ��A\v�Ÿ�C�����x��mR��j�xC�MU�֟���T�����,���c�s��K�"]�������
�ۻ�\r��SnT�"3��Ԝ���ڦ�� FN=�X�G|^�"�wP���@N��H�(�7���K���88?~�\���ta�r��l���y�j�Z��p?�?x�6��o�������Y	�����YL�f&�s�����0����,�ZB�\��K���F�Jx��r�ªr�aLq��jEE��Ya+��Ц�e���G�L'e�{�ế�MQ?�BR���M!	�<ȹ����<'̧c~=��Y�0?kF&�����ӥ<<��0VG�����Na��&� L�>��>`
��+���# �0��F[#������Gjh��65"�AEd<�*L��J%G.:PJ�е�P����
��7_�3SD�%Ų���e+�Eq��Q�ܵK*�m(9j5ƄI�J�Ra>�?J\������ӑ�,�N�~b�j�� �_'���ҩ�c2��t�����2q���k-���M�LtvUp8fw�Z���]�yk(�������jN�Ŕ�t�%�f���L���Źt��M���� T��c�c���6��A�Ç��$�Je�j�3�)aNo��X{�<��pbx�^z�p ͋�a�k��Ǭ����T�%���A6�OI�x>�w422�҅^�Tu�U���B�/MWu�P�]��4?�&X���1ڷH[M������d�-���R�b��ԩb��!㘡w����'3������EM�) ��Q�Q:�S@�v�$UD?��\
ǆ��UB�[E�߁��3ؾ�yl�������5E{�b� �� ���n��a���a�(������g�r��� n���p��c,���x���A��v�_���F�L}9zXb#�[��[A4�A�Gx���r�R|d�Y�)cZvǫ۱t�b<��fD���A@�Ykο���}^|�5��t"�.b||�bA�����_#_��?�t�+�wbϞ����m~d��x��X�����)�jo��e� F�L�2�nX�K��
�0��� z���	|㶻p|pP�k&G������([~����B$�EbrW^q^|a��o��$�[[��ەq�(:&[��J5��;�A���5�>�FBֲ��Rd?GgA��-����d�q����\��?YYDHRh�ǰ����F��Oo6����V
��#V�N��������/R�A�AX�1�Xi6��=
�)Z����0
�y��~��3ߩ�����M�Q�AțÆ�m�NFs���]~.4�������S�*�j������ �^������ieApfWH��qD�U�}ӝ��deB����b1��Q�jى�3���_�a�{G�	�qCіY�`Qj>��#�1цM$UJ��Ie� �Z?
��A� ��=Sȫ�⤭�a1�'I��MXt�J�'������!5� �!�;�v"���*���V�%�d�"�ɷ|v<&�]O�B�&�eHK�X0���NՃ��^��G����L
��4b]�|��B�ۏt6���[�t�̄YT�V����1�Z?�/��TC���z�S���#��:i���^a4�E����&�L�=f�o\���jk� �ƊF��z����C]Y�cr���x�.���宓�}o�=��֛i�& ����AU��A�>0��nX�{ճ�݂��˪=~�C����	���=&����7n�\z�۱��<�e~�ȃ���Z��XCc(er(N���Z�a�(֯
 я��yS�'�@�*��7���-[���1Y(t�C�B��D�V+����z)����t$��y8��&M���p��l���x�9�x��P���\��ȳ��lVi����#��J%)�������%��r���`��^d�i>
%���1���t��)l��^͉��A�2`V\X�j-��r�*��3RuI�V�3Zq#��c���ع�n��;px���q�Շ�"��B�&ڵ�4\�����.�<��9x�E�z,�E�g�y&vt�<���2S��?�[�n�µ�~H,����X�r�[��w�~�9�L��0�>:��Չ��Vছ��i�+(��^�# ���!\t�p5\v�[����͏�U+���A4n�jQ�Y�e%r��)S�FVר"_ȁ��hĪ���1|馛q��q�n�4r�&M�''ɬ5!��d".kB ��������~�����>�H�"�\>�d�[쉴�,͜_��l&R����5��D�,��;�ްi�?S��s��j�i����Ɍ��e��5����Z�A�ތ��ÿ���Mp=h�g����|&l>��F m>`���T�0��c�F�U AX� �aJ��_�xS@}������~����.8�Y�JLÅ��jX�0#;�3���o;��4��4j�����j�nc�"��z���̛�r�t�W�|���p�l���0�jp`Z�g��b�L+�VA���Qu#���� ��[,*���g��f�a<�0VG�~���b�kj�'��YM� 	�a�0źPB�*Щ�h�OF��@� ,������l�!�ٌE�W�Dj�%���W4ހe�W6T�A�倗��e��Z���Q�+�xO�c��	�Y�����(:�[�N�P�La���>q�FO����L�^�J�1����Q�H:2X�I:�[��SR}3Y�$3�5��`����)����M�0^?����3�L��4�*E��h&� ��X,��P�.�����S��	��7]-��]�����ےiaZ�`��D�GWb*Р�Aa�w���f��AX}�O����EkR�O��^�������� ����n��&�R3�W����;���Mx~��p��Xz�j�
`�_rܤO���.bi�.S���f���z.ۍ��3)�'MMa�T$Ҋ��*����	2,0��&`������4)]A�C�bl�T�)�������O�o���{^{��x|�S�?>Oo'���5���yl�Ф)��g#��4k����t��҃���<�n���1e��
81zV%������ ��V����ҙ<9����t#W4�	k���5�c�j��B4܂B	Xе�?�_��w�X6��gu��%����)ƺl/������R`��!���L�������UW\�+/�L,n����)�}~�{���矗v<��br|B����;�z�j<�m+z/���vc�s����C��K_�W]u	�ā5SX�CG�����3y���l�#y�47ߵc+ʅDÔ��p�k�7�.�p�_���j#��5G�W��=�q�W�.��gd��\��,l���� <�F�e����Db �|F�`/mۂ��#fR	��g���2� h해�Sij�Ԍ�mJ���f�)�
�5������&�7|�.6n<[~�g�zMH(&n.����k�.h�I���R	�u_��xh������S�`���Ǟ��Mg��W�2���1�~�7�U``�����A�0����K�7�Cٶ�Gwn�ѯ����4m`:�R�A1?�x��q��S�՗��s�������Z@�QEU���5E��?��B��SB\E����ޕ�©��'s������b{Hq����@١���t�g��e��%P����k�ܞ�IU3��GY8�$�I`XX��%�����D��+֯��Ԅ��"�u�%��	c� ~G�c�F�cp<��y-��"F�_ݍ�t��(�Zл~��r��!14���D��Y�yg�x�4�(M�]�Ņ�7�)1kC{��SY�����ϙ�	�h�Qe�6Kt0�` �ی�/��|��tcb|g�� �HGG�E|ﷀ@ɀ7[��X��ȚIf�����I�A�B�7�~7�'����ɩ�q�s"F���q�'Zwp���E��� 	s´_�`Ο���H0�L'���z�a��g�q�֚/��"�¿���tlSE�yhRH ��2|�Aͭ��:I���k���>��
���:�S�W��?ٳ���`8�
T3a�����?��pŻ���.KV��d:��;^B�&��M�5��45kbM5
�,\�~��0�����gOD�#��I)_𕜙�j9�T:�'�n�Xp�����
�rO@S��Z!��9�k�Tb[[�g�[��U#h|sV$�E��
�a�ڵr�t@������	6���S �ׯL����e��=#�Q ��G�`H����I�d�+��s�����jÎ���eˋ���T}ǚp�[Ηc�Db,j0�L���d"I�x#~��_c����i��������p�|&+��Y4��"~��E�V� �+���}�_z����&L̯��6P�B�` {�챽��F�Q�Ν���#]����w�'7c��]��H>�W]�����)~,�Jw��-͙ޠ��JO'�k���8�܉ư-MX�T�%���}�eD�f��D�,��6Q��G-�b)�������_�����yn�y��x���G7�,rL6�d�XqzL�շi��G������L'��eՆ�G��1Յ�k�!f�{��H�]��W �c�s^�U���l�����TbBR��h���2��r����+:}(���Lv������2��C�i6\�e�u}��c�
DiF��b�o����N��*9����Z�V1A���p����0��cg�r��~�����2
�$`�;��F����+����8��,��*܎
,3�����^V��)�J��l;��wٹ�C#N��e�H�m��FG'�Ob]�4dц&iY��"3TM��e����9�}a�ɶBb*�D�d�(�us�X�"�Ŭ��Y�@�p�Xy���0�dDX�N� ���7����T�;w�z{�`l|~6�6-AxL"� ���:j�<.�;䞭�Le����X�q4�u� ������HM�@�=�B���n$F>��o��n�J�J��G��1-X7k�G��D�2�e���+%�U�X�fF�����4ad�q1�8�(e� [&���`*�J"i=#?�,�Z�c�T;#������`�5��J�v"g�2��#�W1Lm�Y	��8aY�M�L�s6�-��1*�i.�t�惬
����ES
�Ҭϙl
�2.d�t+eTjJ�� @�B��A�.X8������%�u��J�;����B�sy�{���j�"�M������`��5��=��[�����+c�'&�}�N���5Lͤ��֎���{��_<�j*�YSi2��K��1E ,���# � ��h�޽r^L5��U�d��>��\��T�;�Qb��pAc_S^;e=aJ�b�F�&����H���|���¹��x|-��K(!=E�7<O�C>8dS��Ƚ%��S�b#`�ŴJ#hz��O���/(n��J�Lc`|�b�q��� �a���&Ǐ݋a��B���dG�5�]Cb��d��ҿ������g�'�.'ʆ���0����ȶB���9�ۅ�t]��s�p����?~��Y��0�F[�$�9`l*)ը'L�2���æ�%���]�LL㢋.F6��믿.L%��V/C�J�_E:<����^�hT�����sxוoG[s�ozA/�y��L!��j�Sf!,�Uу��8�AL&���]���p�����[���!�J#���M�9�Ŷ�Ʉ1��ֱ�]�����{���L��w�~j��g�نƈ\�\fν��V�)CQ�͍͊[󦦒b���DP�MS���7 ?�|�^���~���e�-WT7�yJå����5a�1Q���?y���,|/Ƕ� >i������1l���كS�8=��f�>�!�z}�����j�e����W�=mS�M����C��?)&�xd��Y_��'߫�N˗-J	�90�޸���>�!��Ѭ՚��7�q^	�0p"Pw(ڮ(�7T�+i#H�*̀��z}����J1G������2slo�xV2Uwhl7������7�_$"�8����"FIA��C�D$D�V�^|��2��I��5�vTZ�r�=�h�\N
y������n�v���Uq�U2�����0-tuu���	іf�E�ǎ��ԑA��.�TI��Eȡ�l͂�
"۳���Ւ�b6/�U���(��xpYU�ۙJN�P�cj�����ejG�����5nr�m@E>��'�
�=���a�~��9fc(]���LO�L&˻Oᗥ'�f��'+ϳ>�yb��b��Qc���]�c��8�%�e����yH~W�:�T�~�N{F	��I%r��Ur������ ��g�o�H�PUm�A�\����0�nJ�1zch�������;��lF�5���FbT�֬[�֎v8�':?j����*�w�bIs�;|m�-�x��ؾ��\>x*���U��m]��"^6����}Q�Z��8�k������W`�͖_��4ȢA`�Y/�dWU�vCd� ��F�/=��	�8ι��I3���j�UZd��P�
J��y4O�B�t҂!��Hv�x��t+��4�� �b	9�&M%UJ���$EB,4�}Hgg�G�v��4B�Θ�3�0� 1n�s�V��F��¸�l������{ ��!9��/d�-W�������h���֭Z)��d�I�E��љ����;i���YF����)F�4�̐2+%ÓM3��Ex�^�O���W_��������G���t�&�m}
M1���\zNGn7Oe8~��<�l��Ma��(�xy�X���ع�����`��cH�rh������� ���na�H1������W��9\z����?��c"��4��YҀ��t>wX���|U�w�Q�.(]+���dJ�U�%㒠�׍�q<�\�W^�ND�a��
C��GU��$7�������_}z��7�z]�sz�X/��t�o����阬__��ة��ͱ���t��p��
��*���)�\x��Ɂ��^:�w�⾊���[C���p� .aQ�]�⦿�s8��#B�H�-A�b�P�Ta9�8��c�I9�s��s���?�    IDATK
�vџ�Kg;��d���go� 0
�k�c7+c
ES@�����ڥo�S����_؅���#�B��)N�{NJυ<���a�jY@���D2�ƌU����@����j��۳�;X�5��8A��9Lu:�7���*������ڌxG��䨇�T0xt�Ǉ�jE0���sV#a� Uʋ���ѩ0�p�a��D������*e�H�� !VF1e&lRUi��D�Ȕ<|ݵպ-jVc�]�Y�@[���0�#)�ݪix���u�]䈶��j���9o]0�;(���gGNTI�̫�%�¿q��E���vJS(O�F�h�w\d�XW��Ѭ����ߙ�de �0���x���1����s�^Cdr�(�QЪ�A���3aev.��l�[�9�*Y&���/�Ub8��y�q9�d��)RWD�� ��+	���K���f�,�8����0��Y�<~�ϫ6(S�6[��O`L��ׇM��@���/7$�-q=��cGO��Cg2�N�h��Kj�x�����=﷈�3ax����7ۮ�cBZ�ؽ�x�x���Q����I�����j������fhY5���b!o�Ӳ�!}aim�]%LKWL:���a4�� ���*�X�F�e�="�/�j�y��7t!�̣��"�&��bT@X�sQ�0�yQ��"70�8��wt �؈�0�@)�Gs�A�����0�� ��!�bâ8���j��\,uf��9W�pRj�^����ȗ�J� [("��BӪ��H+<��%�sA%@6��M#ͩw�ޅ�Ǐ!�J���/ߵW_܆+��6�[���������~�=Δ�VS�e���l�ǧG��aZtշ��w�`�	|�K��I�o��]�g��,���xB�;��t��]���n���c���([y��3HM�����G���Ç��N�|����&Eu��b0p��X��8�y}	��`�+���6ԤX�]�J���-Ob��tjR��y�I[��5��̓��h��7b���N��u����&����ӀQ�ou=s�?�Ճ02aR�|ǯ^:��⾲/.�H��;�4�L,m�)|����#�O5����3�9=�ǚT���G�pHI6��Jv�~}U�_�]��`k^RSS'���N1�2D�c�q`�dj`��UHN�𵻿���"f�LL!����2й��{U���a�&,fJ0�Df��*�q�I*�2B.z����;�����L>����3���tN�&ޯn{�4��������u��Ibj*��q��A���m-Xv�rLYie�0݆8�P3�3t��[��x�pQ�̇|66'pd�6i5Ķ�k�0C]���b�\g.VU���M�(Z�1����>Y $�\�ؘwv�&�VS���h�I^�n�@�fF5@�B�����cAW�Q�Z=IG҆#�l���/��@���f�4����E���@��C�M�szC���Z}U�;�V>A�q*
���a�+
��JTI�ZvjRګZ��w@�{����-��F( �k�v�zL%��P�E[��wȋ%+�#��[��Tn��E�6̌'h뾑rm����1�NP#-^�6{H�JnLx�x����#
<󘜇d?�:1�E�-�����Ӎ���Ai�B2�N�s���L	���ػw/�.Y��}�ͦ���$��ƾ�ρPHz �i��!�̒�^6�p��2tF0��>��9��C�m`�,B~�=�E*7��&V,��N��'&�s�Ĝ�Y�yBO9�Do<�6�L �4��&l&���H}������>d^X�=:9��9�_	���OX���K�� ������o���.�{�y��/�������r�j�'{w�9��Ҋ��V+֜=�L��_��wU���y��߈��c&���s�B��Arr˖t�*���F6�BE�.�(�����\�@��7�c�8����ڶ�=�	�|�p{����F[{'����|����>4kDcS�F���Kq�����#�f�j!���Xy������}�x�.��K�=��$j�֙��m�t�2_2���qQ��)�܋/�{���ê?$�n���H������ �ڌ���L�bz3��0�N���5���Z|��������/8�9�tV}�����=N��Q����&�O.��ٶ#������[�7n(TȄ%�4�hl���Ӌ�Z
��Ȼ�Ɏ�Q�D�YAt1O��f�N�<x�z�.������7C��mc<���T�ݢ��0��hGk�U�&q�(��@1�桍��J���v���lٌM�w`��Ym6�%��c3�i������:k�"+TJ�^� �aLgӘ�gD˒n+W����Բ�T���(������t�Oj�������'l]��>��s/>_@#���������܈���F��M#��V�[k�Z�1*.�YL���X�l`��-��h��@r:!���Cu7�<
�-j��(��n�ށ�dJ�<�|p�i>2<(&2����ޠ4�$0�K�)�F��Dק@�N_�{8��t�A:�Hk���L��H��~�5<��+#ެ�Z.۶����I3X��(��c�v�V�t��S�mg��Ts��ݝ���VG:=�s,�T�������B2��ZSW��#c:��%Ÿ]�~q���5c���سw�B���J��Q��g��t9[@Wc3��v!�̈3�2'����v�©l�D�E��i:��mb\*� 畵A�JC*K�S�Z�7"0�0d1\�b)v��!כ ��՚;
�y�y_4I�	5:�nd�x|�r�'������p��4���ȑ#r�M�yVM�\�,6�
�P���0,�*㞕�#�C�<�����a���ho�à]�QC�i�
���0�и1>�Eb*3_Cc�C*���KM��av
�^�iK&�م85a����+�YTAbj
RH�*N;�,i[�6�p�&��//�[�)�㵝���14:*��dl����IA˖�6���ƻSb�@�l^���<_��ga���AK���b�p����[��_�]��8~�z{�Ϯ��l�w������e��Ie�����Z:�����%�~�j��흽����+{���]b��ѵP��i���k��߼�6lټY�~���l��-��nĆ��P*�`�r���Gg�ضmz�78t�%S
}.9nY��F�(>��e��jE�T��	�&;.��ߋE==������2��[�nZ�"y\'+�ŚB��ҙ�����엮�<ѿs��c�.ұ��ԃ�7b��k�k��o��u���p��$�GK��u���}v�� �>aR�0Ǐ6|��?����P��R��R!	���Vt��UM�s���~8�\>C-�*B�xv�|���q�RM%�I "V�^�mތY6��ŕ�gM9��w{Pr0`r'/ ހ��0���a`<1%)Qw,����7�|0YEBA�YU=&)Vc�H;ɪ�p0�����a��յ�S9Wu�=ӓ�FY�E�`2!��M�L���ls�� $!#���@�Q�(L���9TwWW�U��~��S3�^��������J��y��k��6<A��<:z;�oYK�,��2ʅ2��$&���D�~D�ALNLȆ�񹱔\����1x�ni���gM�-��JҀ�����&x�n���ʆ���152��|
!�/f�ѕ-�0SH!�o��MQ�H�Ii14<���Bb1��E��������L�!�L�z��lz���LlCU)��Ʉ�~����m��m�٪hnh
�W`)VQ-V�r��S�*�4\�-�Tv���uՋ��YO�ŠiFLI��u��Z�J ����ڤLA�r�̋Js)6T���y����C�N���b�gij]/ ���5� M���i��3;��;����K�giʿ��y\�pp��1auYʾ���k�n���,�oZ���=GX0�Nx�"�s������ÉJ&��ۇ�`J����2��4��ׇf�	㼦9Y)�=�摦�f�s���5AG��ԙ���m6aLer3���2��� ��V\�5H�)F����x��9�y_*��.�0"/ܼy����c�ˁ�Rj��a�j媀
2f�JǇ�a6>���QF��@{c"!iv��	T*6�\��9��{�D(;�sEP��cl
TO��ZVlv�4t��
#N���j���G�c>[C�9�l�CU
K��g�н?O�D2��_�~��_���oGCs3FF��W�� �o���]����+��!��瞋}�������r���"x����(R�2~�����'��[�y%xc?�ŹY��_^�ΎF���K��V�u��1�(!�e�<����Ǯ��hhl�%_���t+؉���;w�AWW&'ǅ����싋��z���W�U���B.�.�"Vėr"���Ǳ}�c�UZ�lv��3�#�`��tU��ö[�\r��P>t䰴Sr���V}+z��7��`@|�t��b��N�&�Voa���eZwZ����$8����u���0���̊����0�����t�������5T��z�_��!��Zl��'�e�,7����7����!к�5u�0aa��]h�����Fj����R5X)8���w?�[�{t���ȢƅTU�(͎���2���O30�ᴀ3�e�p�j�|^�P������Kq�#$�$2Y�i=P-��JL���r��o(�9�0�(�����%��*���ndKy$r4{,���4FC�怣 ����j��>�A6���.�O��='�8)�:����-`��^q���zSӘ�����B�)��QB��K�"RբXP��.&�06���2K�imcs�D�-��R�:=]'i����xb��s/Dz`��X%���*�����l	�X
��,gN���jL�0aJL��Mв��w�U9U�~22R��k����ӈ�:eō��qq���#_�4 s`�Ľ^�2t�����`�	��zVJ�g�d���'MWO_x��Ӂ�6/�ݲ��,|�gQl��_��ժ(�
�׍�[7axt�h�]x���G<f�V[��YZY-�	#[��.E'�zv�Q��Rk�L0����n���7�-F�:m��|��JT>�`��#&�ubp�q�0��b�%ϹN��sN�Lijo�7�2^K�%3���?�A��Y6���0o��s�<�1���X���el�����X�T*�=T�H?��0��%�6�����KX��X�`hx�}��x�ٽ����a�#�Q�nQ��>��h0��l���˟:&LX:-F�L�.�Q�/`Ŧhjj���l5g��p��~��G���{����W�@wOr����i�x�;�)ߛ�<�����T����`�k1��G?�A����	V���Oa>D���3��[_�6GG������E�tZ��^�7y�ݿ�Rbl�Ca��踴�)W,�e��]��ʢ�D[��܁��ٍM��"��bhdD*�y������:�08؏����돐����yJ-���Jhi��V�������L`r:�l&��h��A��i	���妾ל���يP2�x<!)a�
�2��<��T�2�֬Y����-bO��'�_�>(��2fb�M����[1j�[�g�Xŵ�ȯ�O}:�~=�g���(��z��R 쥘0���<i���}<'��U�0�ۓ^���x9ZT�x��Ko����,��u�#��Ѩ%�p
�����#;K)�
X�b�������y O�G��;$�fD@�Z�X��+�z��1��$�y1�k���"� �]��XY'x&��C�e.�y[تVi�CA����ی��Oz�x=�	�
h_ю@؇L!��DJ�;TS�F�#���I��-oÇ?�A��=9��x�	��]�_�{&c��/BLoa�*4�͎KϽ �F��W ���G���4���kU/f�It�_��׉{X����8�{��*b�H�ݽ=hlm+.v�@GF���BIQ1���E*�r�7[X�Q��rR/���f���D�7�b<'ͻ�U�dZ�f^3�Ubr��J}Ճ��b�ꅯ�R�f۪�J�j�7t=i5��d��d�h��udz���%#��$tP��׬O��7.p⁥���zSp�7qF�h�}j������5�%q���U�<^n�r3�T(��,��G�"��H��8?��%�reK�x�k_+�6��XU9>9�l1o( @�=H-�2:�M���M���0=i"i�0��\N�Wmm-�XQ��Ҍ�-tԮq��QZ��R��@��2P&SF�:j�y�x~53&�L�^�)L����z���ɞ��);b�|�rq	�r��1�X�8߃my�Õ�Z�ui<����KgPȕ���.���8���*�)lGwk�Ꝙ��Ù�^
�ӏ�~�;�Π���N�b��#(-��ا� �&Ֆ,6R�|��gυ2[�ŵX���O���������]�=n'�.'<^'c�,�p�?����Y	�Ãؽ�twv�8��&,�H�&��������YI��⎻�g������3�����g?�.�d@�Hd��3�b����?1��/�Acs+2��	�\Y�zV� E���W�uW�?����[��9J����82����_�c-����Yj떖Ҙ�����b|^���M�tdzj\R}W_�)\��w��8��!�r㹧w�y��ݵ_��� �"PC"UPU���$��:h��4�>9q�AǔJ��P��J�q�2�rz�p�쏌I���|;#Q�3"�im�$)����L[ ;��0�+���ט�?S�F�룞�z��ڳӃ@��N&E�ԃ,�J׃'�Ω���s��sRϷ����z�S�}|�`y��v�a'{ ������?���Zo�~���M�`�:Fb��a�,!�c}���8>��+��M�Z\�ը�\2�*<�&<��>��������m����|�j�
�/��h�*BI�U�@�F2U!V��KVa�~��Ve����B�=�}j�HSK2;X�.|f�m�z��>')AX��C��nx�.�MO�j�]��-49�D��3_�;��|���lI����W��;����`��l7D��9q��3�7��+ĆǱa�*bb|+׬�������o�;@�gG���p@�b���d��Ʀ1;9-aj&Z�Z��ى|� ���ԴJ��l�	Ff��"��p�Ծ@=�]����'�y&��-�(��E�T�9�y�7 �U�jM�/��Du�K�/�8�1�0V����i'�#~�!���]5 �s�]t��=Lk����/�丙�6+u��z�����<�BAS����/�:ť=֤�M��e&�ߡ�S����H�C�$��9mE`]_2��	����%���ufڅd�a��7��R�862*��{w��_|�2Y��V|��c�cO�."0>Y"Oݤ�܀BA����3�4�0V��ƪ�&dy�uT����!��g���	�c����薬��i����r���Јh������:�p8"L�����b 2�ɤ0a��Z��&���Ȉ��8�عs�ɤ5�q�����Y�L��R���+��8:9�X|6k=�!ثi|�����F ߹�G(W�pz�(U������5;X+CF�� ��8R���8:0�٥�Ч���w�gP����
"jU4�`�����k+�WJ�_�*��r)�����jk�������E[���@Gw�P�p@2�0:4��o������5�V윳���n���1�M��w���#i�>�,2�v�=�bq�Z:=J;�O�K�a1N�k�ebbz
�	47�!�T���UV��f�:47�`�D���p�x��	-z�esI��`ǆ�}�j��}o�����|������.@8��_�*�ܴ.a��4�CR�R\�5Ϫ�Z��|��Hj�,��gf�Ã��S��l��RAZ���x���*�\/صAO��L���UR��҆
�9��7�Է S��Q�.UXfNg�4x;�9��t頒���Cɢ�ߑ�P������\�O[�����s�Y�/���_p�\{,��F�/�����o���m��e��Z�e	A_�\��u)�t    IDAT>}�끥	�*K([��#�d�w+z�y��]�90�IK����mH�H@�d�H�3�}J!( W��d=�_Q�zp�r ���ZG�+5d�%�_qNUdPRਚH�� �J��[ʹ@�Js.%V�a~$�Ya���3��0���`�a<��C��!�|^y�6��Ո��Z�1���X?�M�����Q���s�U�cuW/<���gg�?>�����#o +7�W��Y1�$H�'�e7jY��M�Qp3�/O.�������� ����(�2B�03��L+'	�5���I��~�'k��-=kQXL+�YJ!������������Ց�s�O�0�=*�Ѧ�k177W�p�qs���I��Ao�:b����@&L�j:Z�E�9.���н#���)��i{��R�`.��`��9��a�Ӓ��|a��i7�� ��J��,(+ YAx�9�H�Ş}{ѽ��?����3��	�U�.������1E�L�,�fu�fkU�߳�1*F���h�N�֧<Ȃ����EU�ڤ=-�8��dK2����bU���G@���΂ך:&jgȘQT�먽��{{�:񹚁�q1p�{�y�ʲ��W�5H���UE-�5�<���\���<s�,f�0�8�QDcЁ����/���m�z_��k8��0=l.�f�bp������*�!�49=���4>� 2@Ϳ�����4U�8��ٷ
c���R�fw��
g��)�n�J3l�H5ؒsx�?�.�LǏ��<��Y<�����������E[ml��]{�{oٲ�R��� ��@8� �<���i�:���J��XZL�oxr�|� �ia��6,��I��sfD2him���n��,,�cv~sS��؅�/�\8@Sܴt3 �~f�s���bi� !�X��IA��Ɛ����G?��?�Qdʢ�ǉ#����EC��B.����(��Z ��n�v��P`@�:�ҁ�0�嚌/�[�Oq�9�^�l�1�����mm#ȧ۾a{a�}R�g�X6K�������ꥀ����N��>�h�MK>�uF����1��V�O}@y��u���?�*�������~�e�~���Kn���n��[6�2�RI�f]B�_��N�l	|����d�/�$�9��?��	ܷ�,x�� �R���Ku!����BV&w�]]���|�~��VY1]z�� L�i|�D*�(H�Ӵ������r�צ�[�]X��eY3�|�+k&�CMX��ξ.�Q�Tln_P���2�>Џ�a��V��E�_ �a<��I�����8<9g4����m�D�X3ҫ�=҈��)1Ϭ����j86:��TFȇ^y�4�>6؏��Yz�n���PCS�4���ؿw����Q��ni\� T`V�_3��Ϥ��t���\̨WK/.���!5���ᅑ�"`�"���ס*-�B��`V��4�Z�NZT�G �d$eVĚ��ZO�}��V���q�U9��,���&iѶTݙ&��|�}�f�����v��T0���<g���5�&A�7T��Z��ȱZ���[f�4��|�;���`���΄,%)�� �hX\�Y�̟�'�f�.�vX*/��(�M���[�G��H�|A��#�Oϛ �Q%�i%*f+)��y��kB4��Q�+�#�*��a��U�OY>���sJ�EA6�!A�b�BƁU�W���	X�FLU�'�����b��GRN�l\�-����s�2���	n�|A���L��aTȰK�"�S�j�A�B,1���\�2�n�u�����%|��kpb|	7��-hk�����n?��Y�4�c��V�۲�R^ie9�V�Z�B���ՋO�:�ϣ�2�L�F���[��阀0��/犋\�Z��R�4v{���,���8���E�у�e�d�*�n=�>��h��b��@�@a�������T�H#R���F9�֯�m�G��3�$��n�d�<�FG�����m�Ȟ��XJ�e�0�j�lřgmƗ��j����������z�LM����%���F�VHQ �#�w�"������y2�G��s���_��/�o�Z�a�;qϝw�1��V��m��ܴbtX�gQ-�$Pb��=o��J�@b��UL��5C����ϴ���݀����
Ȁ�5�y�T�r��t�3�M��Y^GX�
�}�r[%s�/��K��k�Ҟ���:�~�ڬ�I������N�kV��Tϯ���g�N�|���ˠ��'v�Y���I�~���f�����t�}�+;��S�D&Lӑ]t����{��'��+qᴠ�v9� �9<��N$�>��JT�F�%�S�Z���Y��Μ,��d�A�ME��~4����(�e�rS��S�N�V����FMK��V�t�g:�2%�ᄨ CFg�8�^a]���-e0�4�Hc�T4V�e�b)L8�VW��4��Xջ��3�DB��������<6^|����l��J���,���	�K ���� r`j�J6`:���ÎM��׍�'D7��bS�͍���{�S	Ѳ;tX�e��~/<-���"�E�7n<�ДE�mk�׼>�l�.����fQe��E����<�Ky��3h6�${)���hHO��b��A���	�vt_@j�H�3�����-�<I��x|Q|��S��,]A$cάv����ǖn�����|�b=�R��s�]�e\���r��t�����>����%�0���G��=	�0z��I�T+FJX���"\�Ӌ.������0��˸=x�-�X�ыJ6;51���� ��i�o���k-$�}��F�5[�NDmԒ�c�� +cU��+�\Rd"�{:DC��#ׇ3�<[�5?��A���g�)�E9�0\,4mU�fLY�%��i����E|��n�bA�ѵ+Q���^���Y�-MIk����Âsׯŗ���z���ӂ���5b����F�~�&�b®�����������׌/��M8>2'��"�H]�VchjŚnOP:�Tp����J�[��^�ɘ��H�!)ɡ�~���}b�0��q{�� S?��-(����=�ab2��|noH�i0���<���7~����h��T�C*��)Z�h��=�n����yD9�+^q)���w��5��P\�a�P��T��臷b��_,���36����\v�er��D:t����/����	8l�48ԏ�^R����Ł�`X��MO���n����Ŭh$X  ���QF�bUaJcHxV.�9`Z.)p�f�ޓ����y|��͛7⢋.B��b2i�Ɇ��j��׊M�׻̾�o�iV�t V�r\��ԙdk��R��Th�徔��f���g�[���L�d�Jʅ��|*�S����:3�z�ty����p�e�v�j����������q���2K×氡ˇN#�O����ό"���g�UC-�E&���'��x
��N�3�� �:
�f$ApU�:p��q�Q@JEL�p��V|�/����f� ��Iu$����@��@�jG٦�I���C@�U��srӪVd[��Jݫ{O/b~)���.��5S@f6������(l��?�a��ŗJ7�u��n<��v�86oKZz�miBOO��8w�F�ş]� �pZ$�id
y��g��_���"}���
܍aT]Ņ6E��se�
�45�i'7���i 	Jׂ���(�T6����lĬc�-�����3��		�e#���@�.
��v/\e+�s)XhTK��������k2_�h`
9��L7
V)q�����M�)M�s1d���2��\�hs��5'xW�{��_��i���^N%9'�qpt�)⦠@�J�8�iqb�.Ѱ�u��y�/�	3��:Xu�T�4[?G�*α���=bqiI�0�0�aL9Kz�Z�T��I��!�C+�-[����n���8A�URqk+��:�i���Pʼ��Lah)WT'S���+��� �K� Ͷ76��f�r��X VJ�Q� �
�V�ڵ�e�CSS�lf�&���-B�h��n�l�菞8.�������M6��D�.Tki�������\V�Z��V}OZIp�(#W�`fqK�9��i�Y�����|E;p�G��H#���,�ޠ��Rɜ���y*�6+ڽ@8 bn�+�k�����iC�R�?EG�*O͡d������2<��	���k:��{؞�\�bf|S���#�L D$Ҁ�٘t�/�����s�!Υ%X-��q����>��3��o�3���אL��<@[kbqDZ0>9��z�e��\�����?�����;(j����~�:�����o����=�.������_�e�^�L>�Î��Q�	�\&�Y\s�g1>1�Í�6ʼ�7�o|�۰�ŽH-���@�����$�ż�P$,�O�k��T�\ʁM�	6�	��� +�	,�P4}�<[qq�`��H$��.SGF���/^�/ҋ����lWQ�x<w�|o�RKWy��VW}�_{z����t`�u���}�5������y�)K���dv�9= ��H̀�dj�Tϧ��G�	����ŷ�.M������[�i� �|iK�����G���k�|�$<�
��<�؅��!��cpl�
[Y�A�*�g%�lT�P\kK�2��5]&(f
��ݾF��b(HYl��"5�I�L��`bfV�'�$,!d`�����/��ܵ��Y���XrO���bu������vv�-
�=�f�i����^lZ�N�%nެP���3���w��V[�1u����k����k7������;�R.�l� Uj�߿�&i��64�H@�d�%���W
��M�BV%�0<0���9���}=BuS ��y��U�.[$@T}�Y�y�.I]2���r���������腛�ȥ���t��B�D�"`��4W	���M�τ��ϥ#�h�h�:%2Z{�q��4�J7�'���MX/�zHq!#H�sܔ	���t�<^+/;������|�s�O0�4H����P�0o��֙�<o���a�`�S9���2����<a!�;��Ɉ0kSYCag�}�: ����$rKX�֍ٱ	>�h�皖1�銭\&+�HWB�������e�{� ����x�g����9,�rS�)�8��s�O����R�/SP�z�IK�CQy>F?0�"�S��d���\�y���q,�Eê�f.�]	@���5��^��R�`�j%L͍!���Zɡ�����.������.B�N|��$V�H<n~���wf�t|0u�JLz��}���翍��Y���b�@C�V�	+[�*���P==i9�2������rF6��n;PȖQ�$���1p�T�\d�9�"g cŴ���w�w�u�����21j�9p�e���]�K���� ��pff���1���Ǟ؁[~��2>�Q$q��u�§����9�}n�����{1=������s��`1�N��[o�ƍ�q;P�e-�����g�߄���NLN�5"�HbaA1�V���:ӳ�(e
�h���cGP)�D���e	�JMZ)ҧ�GvS�WvYS8w8NR�p�YgI0p���e#r�.1����,ߟ)I��y	�8~E�h:��^է	���Ic'k�U��7�u�c�ԧ!�Ǻ��5J���:K�����#������V�ڠz�ky�3���L}ީ �j8������|Y�0�O�<q��o��M6_�F��Jy�����=At9����oGeq{��"��8�r>����Oh|F�Tɢn��F!�ya�L�~%P�*̛���z���t�[	�5t���Vgf�����a$��BŦ���C\��4{F��� ��U�	M�tA��5+�/e129���vѳU
e����sX@X���u��UlY��'0?C)O��~��;��s�xr�<�=����nmÙk6�ڿ��@G�P#��뮻����T)��K�8XB^X"؂^4����&�GQNe1;1%ƫ�����m��-iY2z�|Vz�QD`G?�����sI�z�v8�J�p����{�Z���4�n������a�VD網�B*���N�i�|T��4azQQ�5�v��9�	�8.�i*(mKPoHH���E��i���"@��Ǎ����qS&��f�|S\4�!�
S3]Zv�������u:��H�N.����S��EJ�e� ��aqI�0����qQ���R��N�d��-����Jۢ/چ9/C��e�r��`ŝ�ƙZ̈́�E��4�O
�7�{�V��D���҈x|QLb�l�q��5�Wd�����8a1��6������ӏ�b>/U�Sdɚ�ZeP�����������M�+�8�yM	�G�G��&5�Ǳ�52r�_gU|�saڊ�VE�Z����Rq�P@�߁�=�x��^��}훈W��|�CҤ{�������vz��Zb��O�V,� ˗K�������c5>��o�D�4\~���PSZW��td�`��6?���E�QpNᴔ�)��_�!?��0�� i�٩q�}��8P����Ĳ� ��q��d�����o!��_���������o���Q��&�M#��G�!�Z�&}l�F'�k��x���x쉧�b��T$^r�6|��W�VcqUN
�f��������A,-�02<��?�l>�������.��/�z��
>��k1?��
�rŊbpI�,,��uo���#Ȥf�u��������A.��j^1���qGv��T��d�Z&�Y78.�eQ�J 08 ��s8�9�Ȍ	Ke��G�qΜ����5�sK�I��׳Wˠ�P��:�̔6�>Li�����[:�����LY��� L4��k]�Z8�z�ӑ|��\�b�΂�c8��|Ω �R���v���0����eeQa�ٓ'.���z�3ص���)�y��l\B���O_�Ndf��9Q̧P���_�!t�pB|f�e�es17����-�oV���D˃�N�e�Y�\(��YP�EdM0���W�2v�x�y�yX�b�l�R1�R�"�W4'�Џ�L,h�
B� |A�T���^������66��4%��4�v��Љ�z�覸��/[8?���W�Ўg�e�;���@sc�n��7��w���E�\D�Q)c׮]��_�lD���ǉ�[����d�e:���"��C��:=N4�6��(�*\���ȕ���sx��q�������@2`�Z^�l�t�LN��i�\p hq�+�#W��P���:�ѓ[[E���#)����f:�T�4A]]�xӓ������Z-.�\�d0EŅ@�q+��r+�`W�f��`���5������|^�
E�{�̹hr�!`���2)��s�M_�ɔ,{U�T�Gel��T���Ӧ�SS/�#���Zj�99~D��� ��?I�rr������r�A�P�����b˦ͨf����3p�2RJ��b�p����a�9�է�C�Ԣ�ttII)q�����	ٰxL�N�hH�<VI�7Ӌ|��ˉĒ����)F^��tZ�>�I��Ѵ�����k�cbU��Ĩ0�= k�M�cE�5���S۞�I�s��d�4�dҔ�s�B���oS�[J8w�*\���'�ݎ���oy;¡�w�"��!��AXFZ�P�984���"�mX���IXlڻ�����;8r|L*[�­-h_ه�������+�����z/��~��4\��˟ �^������@sS6�[-�Aj����Aw��-�٤{hx��<+UJb����,�d��X�C���뗴}����C��]���\#ɀX�(!>�"���#}l|���<��N$�r�FsKʕ<�}�����M`�(���d~l���11C(܊�i�B�Θ���
�G�8�0�A*1�-����t��E1fe��jP`f`�j�%�W[���_�LX0�mW�`^���ҀKg^�Sfd�]I��"im�ڳXp�b۶mr.�O�Q5���S��L�a���A:yX��#�{&6'~c�I?A��d7�>�!}_�W��x���|��D@��s�z޷�&�a��F���    IDAT,��3�kX�s��+��,3�|��C�-�����s�W&��$���<��;���-�5����ґƷ��q���w��k�O�Q�/�i$��m�-���f>�7 =5������\"��Ua�_I.��I�k6ӥ�4�T�aj
���[l1�p��*���NTX���?����f���J��|Ɋ�Ã�� �]�H���bZ�!��)f��|Q�5%(	=���=���B�jM*F�ӓ����H�%�����6`S�j���oK����Ex��U��,n��ϱc�>�>r5��HS:�:�K���K^����gQ)d�v�Ϩ(b�G�{
���OIZ��fΐ�p ����~4�4�vct`D�a^�6��kW�%Ao_/�f������|\5نM��( e�����%�ө� �\"�|*#�z�[��N㯯���q�ztZ#��ʤ`6�[1U�P�q"q��S7.4x�����z�K��I=1}B��EoϞ=�|"�%����>w��ƅ�&A4=��N����%+�M����o��8Q��4����-@5�o�tO6��e+([ma�J�iL�u�o�n(͔�II%��dZ�,Wc)}d��x�y����6$��tM`������[��D�FIQF:�Ͽ �׮���K�[��`��+.�Ç���s����T�&D/+Ӏ�s���J_?89����cI>Y�BQ1���<'������V<.nhZ{G�>��7n�(��ĉS�?/�#�.����i��e�ߏㄟM�G�J�����|�K�#��}�xbʛ-��)�B��]u�(�J*�k��g_���n��Z���p��ߌL.�{~
V���mB[{7ވ���&Z>�$�7>6���drIi}ı�J�����_�tZ�rg�����L�T��������U�pV8,U����G�O����?���Ʊ����ރh8 פ��/}�����q2��[�ē�cl<��9���"��z�F�s�-�e�H�c�.h�����i�F>���xw�y?<��k7��/�������� ��=�p�m�������(bs	�cQ�0����7��gelV��]xd�v��w��	��&�X*�����pJ����p��cbz��l���$�EL���e�K�:��4T,%4��8�֦F�#�k���U��tB:9P_(�ٱ�����m�b��p{D�Y�8dU2��p3�#���W�Z��=���Yh���On�G�{�#�Z@���xbI����}��#I���j���0��R`c���t6#������,��L}1�7D%�J7ZM1 �Ք��Uv_��}��k�dZD
�}�2~�3ҥ�k� g��˦��yd�i�
�aw�Y�v��^�H���B��b����Ǉ�j5���v^��_<|}�}�F�ˇ��	XJ1�D�X�tF�ؕ���쀳RFviN��Ak e0gs8hէ�4e*��ƄU^:',�i�h͑M9JC����LG݌Й�)H{[���͋����xl`
���J9�e��N8-6�XĤ�!��$�-��#��A�L-�H�S"����c��8�Z�l�;_�:Qw��9���$�}�����ǐ,�ii�B��p�<�|�D~1�Y1�h��}���o^'��5�+{�U�?�L�8xG���[�I�b�jL/�о��֯��il������_��W��75D��	��� }69��>x@��j�$&��guZ�����HW���(��@����4"��2D5#�����+�ŀF���h�dA��<�Z�U� o>���Ӳqp��̈��Y�q\��5܄�(jDk�tJ���U�C�^���8�5��Iv��#��RU@ S�ʳ�a��U:T��1��*0�E����S�6-�{3��l��-W3S��0��hSR���Q,U��)a�İ�O<ޭ[�b`h��3��bw�[vq�]�A6���ԝ,{����q�t��q��v�ycp!�T2�,��"e#a�p��`[�7U��UkW�q��O�������bA]?�1�s>��_�y�.���I���?]�A$A5�a2e�*J�̮kM~�@���Ӱafz
�\�v�]V��&���o�}�jǡ�C���I�P�I�O��V�.��#�� n���`���.g����cp|N6AF�pm����Tibw
�5���-�i��A�E9�B|�ZW��v�Yxz��͌c�;�M%Q���L`���:#;i����e��D�(��Y.8���Utw6���/���_<��w>��������԰�y��I��;$�J=\lvg��U@XK[���p�m8|�h���cx��¨�"���| [���j��bC�{~+>k?��o�gQM�=�/�t�w����E�K��lV�oC.����Q��.8$��}�s/0�\����1l=���یV,�=���Y�AWg��!�),Qc[N6�]�cf�~Sdq9�|�� �6�U�)A=W�3&�:Uݵ�c����] T �]�xԅLڬZ{�q��=\��8��0���ȹA�/�.����iQ>����DR`�v��%/qHl�]-�s����D��*h���uC��dP�ӻ����l=�k�����]:�G���w����H�f�B�͌��3{�� >�Fa_�̇`ϧ�f�)�E6� �����]��T��Bӣ"p!�jd��5��e���ǋ�Z3U�#1g	=Ū��J������e�����x�������C&�X9/e��]@+�$��j3��� �°��JE�n�rI�/%$�шpt���Xj���n|�k߀Q�¨YP�e��g��y��ȣ��=�.��u6���[��UlC%��ۮ��X������ZV�"���f�5,�/ _BljF�*1�t��	�v�4�4��`az
����LK�0�v��(�j������|?҅�169�l*�ǅ�׏��6x^>�������H�D)�����IG}Ō��)&L�#��_�/�0�\bD�IJ�G���2�0'>�a�L����y)�_\\� K�&sF��Z[S��.�\ 86��R)D�̅B|��'���{J�>�Z��=Ƿr�Vƹ'��ja�|/2������A�0Qf8F]�D�ZSa�
�p��a��Q���i%Fʌ^���^a}�	f8,l�b:	_8��ج�Л��l퀫XCz>�遶̄�����-4�㲲R.�����hX ���0���r.j*��E� ^��Yb����&�Ug�b�Y�'$�I��A�2i-/����5Тan�7��L_w]���n@bI�+�e�x�t���T���3=�*�X������#��:��q�Y���׼m��'�x��p�P��!ܼ�,��tH%0q�"p:�;�t:��E	�L3s|�_���T���_�A@���j��a
`������k3S(������u}�3H'���M���*��Z���zq�w��v�<X�g
w`q)K�?��~Y���5�|\�+[�%�p�yga||���َ��%<�سp�iEҀT�թ�����?ۆ�xt���Vvu����=�;(���s&֭_��~�ALLNcrb3�	�<z���\��t�d0;�{�eb��N̡V�F63AƬ�!���$#�`� �*�1jH..���4�%�~���M°��q<r�g���x���֘п�O=��HL�������h	�@Y?�t?���s����`IK,h��1͛r����c�s�s������D�*V��1��Y�-�|o,�P���a�4:/(�[~mq�c��y�A�+��/�֙�<i==� ��i���|��Uk�6?���^V �'�'����[?��K5�f_���Ch[�v�Aw~c��h.:c�L��2H�ϠZȈ6��4]�ij.���^YjЋ�[{�,WJ�e������z��hK���3��+_���dﵼX&X��v$lN�t���=�B*��r^D�n�X���4�AX�R�?��턥Z���+$�@��X|I�F�a��c���\!\��|�+_��XC9_�ֶ�fL�O�o~;v�3����<�Y����+�=z5���Uų�=��ȓ�K�5����mE�̪�E$��-%a�d�]6M������+����R�1x�D��ZI�/����lp�����,� ��� 2NRF,�W����C���QC�a�ؚ-#30'�(���p*�V��Lm	��}_�& �,߮OGj�s2+l�+Q"S,�R�5k��j!�����O:�Fg���X�Z��W�u��{��!?W��	�KJ?^^8�"E[]贚�aF���(�Ǣ���&�S���H��|I�Ś���Ƭ��=���T�1RKĶE��	C��H*����_��|���|��E~t����Ғ�+������&T����+�ul"T'�fjXD�cV?��mP��PP��aa�a�u�)F�Y�Je)m3����s��3��w!����:�PU�d�Vȴ�M+��k�k�t��o]��͞yܺʖcK����*ퟌ�BY6UUQ���*�d�T��S��H�ej����E�R@0���7�ǋƆv��a�����M#R\�0U>�er2xu18-��~L���ٌ���z�e��At�^���)IEZ����m:��9�l�]���g|A�aMaV����^������a��=��֭g`dlT$#�S3r=���/�3}Kc&�`��1:>�/$� ���/�[��F,�N�m�gw��s������X+ع{�rH�r���G2�Eg{�-�X��o|��ؾ�Ai��,���@�(jU�lI�g��ή���x�'�N�i���E|1�'��T��C�ٹ����9��ӨUsh��P�-ajlX���!��B	㙆e�ǱJF8���"�"��c��Ur<d�X�A�#�0�h��BH WVF�����/�K���6�Z.A�Ǥf�4�K��F�e+�q^��:�3�q^3J ���^�$ĕ����6!<�v�s�$�N3�5�Ǡ�6>�s���@�,�*�i�4��������lg��'χ�Ģӭ�~-.���/��T������ho�<���u;*�X,/�t$/�Ϟ�������Bmaw"�N�nKc��T�p`aw�oތu�=�ii�Ǡi`^�52���!�a�ݢ�/�&���m�h�,w���͜���b�YT�&{F�q��Q���T��\U',�i�7��wx�G�	̳��G�*L�������~v��Th�H�$jĺWv0�K-a!�T���əy,N������\����
 _FS��'��j��o����P�A��q�������ro��Up��4�U�rT������a��ͨ�������0�ͫJF����wl�4���b�%!�K�ȁ1p�0��4�X��K&�Y[�F<���wEl���d�Hꓞ6Ѧ(^��W�xs�� R��'�9N�]�x�5��yЮ����f�� �ד l�	���? az2jf�������ˁ\Nyz��LRb|�^�(a7�P.n��C~��2$p��u��fZ� h�L�VXf�4H�8�3���+�0)Pk�1Siӆ�5�˓�BU
��3��S4�K3a�̗�SU��K�b�S���Q���O�D���n��ĶmJľj�jˢ�������b��6���[�31q��7"3�̩��e�U��\�t$�S
!�-}��]�n������,|�+u5ܔvh����v���]=¨�1F�<'lbvJpk6��}�0΍�%?G/��n�>Cw�Ћ>?_ k�(��0�����[���Uٴ���>}�l7�9��v�-2{Y)��>O#�F�S���zHf�vJ+X�E.OP��?�vҥ"\� V��( �Hy���5�ղ�%b���\DzvZd"�?�ڛpޙ�'�uSC�5.���#b�+?s.P{�G07��t��������QY�3\�(�dp��ލ��_@&�Bc$,�DW�씞����ţ۟�,S�¨t��.}Ņ�GG{��鲙2��>�d�s.(�c˖MG|��Tm�5�n���T�@(��ŎB�ͷ�-��Wdך52γ�E�mi��THczr>�M�襧@�a�m�VQ�+]%�	��3��" �\Q`���M:08�xR�XI�K[�DZ@�s�=��g������
&r�ƨ Mk	�}�_�S�z�#����s�+����L�k?H>�A�����<��ù¹��:th9��g���;v����3�@��}V�?M�g����@5`�Nz��Lg41#��j�ڵ��=K,�a���6������m�_Vf��Z�����.���n��-Ҿ1]�s����ڌZy�ۋ($�����RM��%x�.[R�2=3#��F��:K�|1}�\�	�d!_ֆ�ǩX`4n���ǆ�hV�J��jGG[�d�L�R	�2�s�Hٽ��O�ā�<���1W+�a�Q�{ٔc�T=�a6[���+�[ѵ�K��科-V$����R��E�#�s�lƧ>�4�(g�
x|������-?B�f�B&��\V��W�Z��χu�=��k��QT�B)���a<��y�|�-8��s�o�`j��)$�I����f��b����[��5��8�����CX�������t��փ3��%fO?�*�>?FFEG�z�Z���t�\u�U��������¤V]�Vtaa¬e�CF�@�ա� L7�V�䟾�΄Ճ0�Ʉ�����A�D.�d�$�-�$}&��4�鞯� 2a��Gc��15F�uZ�����BQ|��1*��b���q�f-Ǡ-U�T��ᲊ�D1o�
��D�&�ǍF�NMG����d}l��\N���gg���>����e=V���Cr엽�X�~=��wf(�g�nѰ"�т�[����fc�Y�h�$ɠ��A3��F[��ﯯ�n���s���$�~gr$�P:'��"
^>���K���Q!a8	���t�ò�(@JW�D�<�����d떏�b���3%�c��q�P�����6lb?�������`�"�[E	b��)����ҿ��͜:ֲ���P+&��D�nؼ(	HC����j�B���'iX	�屘�U���ѻv=�&�A�e�U`��uM4®Q�$�E{Sn�E��G�㶋6�}�R ���7�|�_@�P��\՚�x�_��LLM���+�:q��.\s����~N4�Ԙ��W���F*�(curr7��1��~4B�^�M(������}}+d����V�~��E��v�d�[�F ����m;�}ݫqL�}{��/q"�6i�NFQ�-m��4�*S�jVK	�^��Ec9�,d�����,�o��lJҧdtV��z�h�8�)uX�v��P�-�:�J,)�7'3�f�?����c�c��H� �w]�����Wix<re���N�� A"�I+��g�}V|̴�Bi�U�9AǺN�s��kt�^W�30|�ނ\|?��%�<~�]����{s��%�	p���5Ov������]^�>�3ֽ� �n��/��v���@��W/L���o��lݸDʿZ@���a�6���l�xJ�N'��Vԃ)ϟ�L ��2h
E�A���]��(�`��"��0��׸�bA ^C$�Z1k6��6�ŧ?�a$&`)��fN?o���G��7n������"b�f��V�)fH;۲y����inD����n���S��f�R��*�͍r"���":<Q�����/a}�jу�������G�~��P���c�Ζ6��a3��җ��hkj��\<�]���׿�+V�!�\���(9m`iS��B4����Mv/n���x�G059)�۟��MX�f%v�ٍZ9���@&��7��D�T'k�Å�O=��|�h�:W�����)����ځ��a�N�x�n��[�p���tOf�nMK�M��H=ş�i �ǘ0.�d�T�R�.����R�F�!��b!�*��VF��!ǟ��ͱ��lߋ�ץ�R~nU"Sbv+�h*`�B��T�i�hy.[R��6FvLC��L�����C3}��Ε�J�Z*.Ԍ���!�'7�0��ȱ'NAv    IDATê�NM���5/y��	��f���C�#"�'�2�8G8���N�ۺ�t
��2�E4���������>�$ȔE���Rh���#����Bf�O�s��=s3 �@0ě6���4����	���F�Țz���?G��Q,A'o����#*��A�b6r�Ap3���bͲR"�b�����	�*�~Q�;Ƨ�D7Y�`����T���:"�q�|���u�n�\v	Cf�9P��p���7bf��,5�]NUq��V�+W�bR4aLG�y��Q%��LXF���������.{o~�kp������O�5��.I���ǰf�Z|�����#�yb!�ɩEl�|>&&cXJ���׍ޞ6�ݳ�~�[1p�������o���x��ߌ��A446��� ��/�T���aqȹnl�Vp߻�x�����l�w����ݛ�J���k����8��~|��_����>�ox=~���p�������a�]���sU�&g値�(���,Y�� c�6��2`�Fa,�J�(^e	�J��&��ιr�U�������=���Cţ���������{��� 2!�B���V��ʮ��_�U���%��EU%llM���$*:�J�x�E���$��Lj6���iiNa�	(�B<��_U�R�8�Ľ�����6!�V{��9J_0%��W�2���z��Z�.�Ka|O�9��t�k .@ѿ�s���j�����{~]��"�/Lnʥ��S!�;g������gt�deX����W�j�B�2�e�Z�|_�����%�WI�(�e�D�k:��̍?����ao��H��:v­���;��z��C��E�J�o0��v��(��.$"���	�f8�g�`%�d4���d+Q�3���E�T̞���j�|��8�E�oGI۪�cX��h��,"`Vq�[N�W_�bjaO��t�+3ւ/~�>l�a�Ls���mZ�S���*�*Ua����Z�X."��	s�}H2Һ����z�{��e͝�T�8a�:!4�!�ٹ��(�y�i�L�a�nb�R@��A�DK;ښXݿ�ЇaR�2aR��k�;߿����+����3:���n�;�p��S��
�6�ek���ţ?��,���λ���y�޷G�DZ��6��2,�-� N>m#2��y����.���1JsXum�����F��ݎx��|ᜅ`ن�/K�U5�e/��9�@�¦���(�����F[_�t�$!�;k�PSp2���-��U뉇�KT���\t >���c�b0ҥv}�3�P\��A��rM�ϡ��e]�>�j��9A���j�G������ �T��&-<������0�������:9=!m���Z.�R�c���BQ<�����G�&D8U.�C����\6 v�DrtMD�
�tE�`���芟L�9�0E�Uc�b��!����M��Y��y)��)AA3�˼'�[�F�0��#����6�p���@�w�ὕH�+�2A�,מ�c[�Y��s(�U����'��������s�1�~��T��B��pa�}R	�D���[�E�nA���:4!mT�/&��j�%��j�:v5������}J��^��P�}}80>5����$."G�0/�����c�����W¬�g�|�s���]��g$%0�7�fgq�I'��_�fg�0,O�0�t���+d
��q�%��k��m���pt?���G�@���)�y�f���?G6�*#4����04tP@ص�^�ɉ	������E���A�����!�ڇ·�����2��ͣ���x��ٟ�[�3暥(<�	����J�A�Z���n��192�x4ҫV����?V�T���ō��NY<��
�y������^������L�`P
C�����#���'m���'<��D`�?�ͧ�N\tʯ�aZ~������ӭM]��^ԕ4� V�I�g�����	�%ܛz��?�{C�m���)��[���7��g��1@s��k%>�mM$i���S_��
�V������l��r<O�ϧ�����Q$*�۶�ч�o��O5g�ה-y۬����A���/���
%U"�|�/d�1X��yP��sE:h��T�~�M�ʯU둜0��3�~	�A�[������L�+%\z�F��ꋑ�A����N �B �/|�~<��ҁ�mSl?�%a�9D
���:���q
�U�t9G������E�\A!�G�/_�B3|�	5#;1����7����Dq~bd��8&�"��ߍ��	�BA45����#�,��߶�N���C"����)�d����H����޶�LI҅�m�p�����	�+Q�Majd��ø�m"�O��Ɓ�;���lw��B���[�؄L>��}w��G����;�I�
ư
�Fz[нl >^�L��9x
U��T�f��v�=t�@Q�F�	���}ۇU�Ň.�-��3���^�@kp%_��)�4�������ԀC8�diw^�m.�ɱ��?klG��M��əiߊW�)*5�Ç�!U�կ�ϭ��V�J�d�� ^n��$g�P߬�M��7Ǣx��W#/��٩i|�[wbێWh���{�2,?vF)�aA$*2#�r�N�]��y!�$����e��T 9�ʠ�۾:x�-���uu��/L>Ee`�֓`ښ� ��p1�s�xx�{Ԛ� L�y9����r�
�tZ����"!9�*墬_�Di_��
]��lrN�4}ݝJ��\ҍ�0��1��!kC0��;�g���Ʈ�L�����E����(�gE,z~�vPqT�T��Dك�����ڰwd-��ț�k�b>+�u�	r�:�3(e��77�H ��<��}��v��M����+�׭�l�6'�b�&L��cv:�X�%���:��P*��[���tv��*��$n��flذ�̼��B��?��p��f(!�k�v�j�����W��N8�rY\�����'?�H$!�d�G��Sa�c�[�r��(�+r�}�I��-���.�2�ϡ��\�����\:�X$�V�B������R����&zu~%����Pk��a<���M���x��[r��(�h��p�A �A���Me\�{E����Ndb���8�ר��1al�i��HMQk ���+n��r��Ɗ�j�*��~}�X���x���(�����1�w�E���!ܫ:Icȕ����>������P(���������{���ჿ��Rͷ���B�b�I�.#�R�IT�)��������kJ%�2-5�'��z�JgЊ�%Ƴ�B�,F��5is3Q!�� :f]mM�uD��<�,����Cnv�zA�N��?�b(�[�{?��9�)ۃW9��5�vPBb��ũ#�G6z�9�����0�b�d�a��v�{	;�5�":�Q\yօ���V��_���N��:�wҳ��ݸu� ^=��lF���@��,Cw�	���cV�Ʈ�_��2�Ju�\��X3��axf�kW��G^7������߂+ϼ ���C{�I;��k��\f3�ڋ����i�M F��Yg�/#�O<�k|�k_���n��oUE��ӠY���/�(�I2QIqɱ,e>1�fJ��r���!�|&T��n΅C����5���Ց �A#
�,<����*�(y�'�x��XGڍ�t���_��#5��ʢm��&��^�E���*�-
M��v$���
��Vn�geQ�X��]�b�S���ɖ��ފW���+.����G�I*���Ǽ�K_�/~U�97пn�lX���Q�����0O�B��J�� L'U�5K�q�;ν��} �{�,��?ݮ���z� Y�ZE��y�)®�jr��rV��>t�?�d��"��g�uП������w8��܄v�d*ˁI;4^�����L��ZgvfR��Z#~k����11;�������)*庨�v;_?��I���l�,�(�{�n�<i�����,�f����b|��������F�7Iu�F��rt=${!Ė��ƁW��g���̧��C9��}�� �>�K\�'נp<� {�qY����!�����m��be(�d&�ZH4S�����y��>�X���nαXHZ��^&'��!j�E�E�v2�3�K����va����i�almm���{Eg���գ�0�bK�uxh^?�{9��/�N�E ����ܬТ��X�UF*9l�A����5�X  ��n"���'*�"��3D~�㑵�yQ\_|=&��U����O�}.t���k�=V�ͫ�I��y�5�SF`-vY�ɗn�2��\1�4`��L'�����a���+�m���%�*��W'V�5���������*���hהF�G:	�s�j�����U �7�b��?�?���/�]ѕa4R��,����`x�IC_.H�n�JXZ�?���N�f�	+qU�
�z����f��I�2e�,N�Q3���"�da��K�:�_~!��q����z���Y9����+���(����*�^�OJ�lY�)pHi/�q���̓�1>3�m���M����L��
ք �/Y��>}�=���œ�>��/o��O���۰u��
yQp��CK<��W�����׶n��Ԅ�S�k��U�f���V̕r��vb�	Ă�X-I��!��	��^�+κ����}0�;b���_�h,���a�L�#g%�����̴+8}�YBh�=�'?�)9��Nd�a��%p<�䷱��S0SH!�L#@�=Y��d!`��Z�.�H�~�����ͫ����5V��-����e�����4����AG�������b Z���?�Si⹬چj���$�����K��D\E�%'�PA�������I���Q�X�0���?����U�ScB��q���o�}�����#�� �s3*�����/}=�(ܱҰ��uX���c��.��~�g�Ƀ�7�#�J�c�D���:��+�o��u0�P���J�.�?���u�W(K�y��9������ziK=u��䵋��V�lc�0��1��mM<B(@��~g̽c�i���e5�0O��R!��CG$�ӏ_���
�.��&����g?����;;�`b|�bf��{7�5���c5�E2��l�X�p4I�7I��{�h�@���LGrj�)��{�|,�)AX��V�÷��e�|�R�VL�M��W_������O��[�\Nb��ߎ�+�K5����ػ���T�U��UQ��V���}�~7��v�����i��b��vU�x��YY�X\�`��I1Z'Ǐk������L���
m��G�"PE���)�L~��	U8EZ���K/7�W^ۅL��T:+S��uXU��3hk���S���"��C�I���Y2l�}˟s ���+W-�u�s�N�ZH%ͭ ��B����I� +8f�\��r��%gEY_&��d����±��v���|�Z�����u��2��:��O��� L����?� ��A#����k�����Ñ�z�8���-��E@�_o����A��IZ��/�����n��b�o*�"��|���?~�/Ժ�\�._	]}� �����FNiݬ�N�Y.�b`RK�VA� �ΰ�����(XsZ�lW������"���e�X��m�b���Ӧ�K�:�^~!����|�Z�*$h&����܏W��x}6���@�˅�|�8eh��#>uU�8��D1?�;��+��dUP0��Xш���:<����	ة����A�6�g�v*�{�w\���w�C�܂Cc#���^$
�ˋ\2�+/�_��atb�����ߋ/��뮻N��_��vT�^[��;n-̺��ڷ{�4�D������'��nl۲c#���p캵��������r4�\��NQ�|�x�Q�_�:��;����K$s���0<1���A֜u2f�i�e��c��k5�⸩8a����)Gӊ���Ig�:8頡۔o���4Ҝ���]lq��
	םnG6����t�K��a�)�X�bZGKs�t��&N��#a5yD&�1ǘ���>��Zi��Ƥ��$) ��I��?����qx�0b�����D#��/���_�f�$v&|�h �{| �޼Y�+A��]��U+09;#.lC��)��T�(B��>p��a����y8�G�%�I�c�p���;-F�f�����X�'�y�|c��k�C�|�����}��K��5X֟U�0��:�׭I}@���
��\�������.jVQ�%���ჰ->�h�ڸpө������������ϻ�//KV	?�V������c���~)��L��}���lizL�K�fE�]K1�LKL2����6,�)�0��o)����;�'`U��K��m��y�xӻ��}O�o��"�E#���߂�ͮ�Y�4ô�P8�\>���ۈ�n�����hD�s�GI���B�=�:q��*���I�r��B� �&�{*�A�bQy�R US���U�En�[�`�T/m��e011��ν ��~���H�(U���b���C!����;����Q�$��lD�����hk�UU�C�9�߯��|�s��g>�<��j�é�kuz�,G����Z^�x���GF��O����I+tP���N��F"?+�l�2����J����)��t�+e���V_����YM�`K�a�3�/=Q�����_�tN�uA����'ɥS������x���~���?��a�o������\��Q���S@{���f.�9�2�S������*u���R��q͢��EYtUmH�g/�lGe��R	��v�S�9x������.\H�����M��܍���X�NrU]ȑ�Ԥ@؞���M!p	# $h `�)9Z����	�/�2%W) �K	���A<��G��9<�&�f2���n�x�	��⋅��R~��Ů]{05:)Ʈ�|�a��iv>���K��o=1��Z�k7����_�*^~q����Z�w�j�%ɰ�Ȏ����Kڻq��c����$��`���!$�q(V2��t��B\�k@8�r9	ۑP�YAO_/�9�x��3x�G���iŒ��#[-��+a��$<9A7m�aښJu����:�՛r!��Pߡ�p@:�ȅ��� #U�V�<����qJ��Qo,�7�!;��mAzC�/�"�A�a\��<�s������H�0��c�/���k���� E�X��e�ADC�.Y�@����qq<�aaU����@�X�e_��.{���).��?��{~��_���noF��Uh]2�d6/��O��p�����5�?���d�N	�AB>�>D�4���!��[|V.4 ��٪���V�^�?�e(H�fk�0�V��
��v�n�� ����X1h�X8@��eIؼ^�X��k�,���phh��$��.�p��x�9g
��W�l�G>�i.]�l��D��P�D�xJ%�t՚�j��|%E����ڎ�ַ�|�*���m!�֊��>��UbXa�0F%Qa#H!gWVz��~t6Q���{�~��W���7'��Y���dۜ��m�@(&���[v.���j��3N?����pß^�b6���I��RzVt� `��-_���e��%�u��Yte��.��QU��j�Pu{����Ƥ�l����) �ˣ�o]t	^߳�_zY��m�WP�:�E���hU�n[���I�����|�)�^����i�~������a��O����I�N@�*oG(W���~�{�-듃T���SmD]�R�h�6P��e~���%ū]^���%�4�\W�5�s�P����"�k�9�4��H�p���������1���J%PW�uE�i�5&�:���hz��|�W</+a��t �����?y�K�x��i�s�nT+s��c�ۃ�9�BjM~?�1�����i�[Q�,3�p�^hCj��a���@,�i�@�?Ï�N8��v�*�Ex��c��*�Poo����#�H��(r��IϽ�20[�p¨J�BZ��    IDATNDeC�\�JH���Y	x�`�����IdFg�h�Pũ��V��:�Ŗ�/��/����j�ٜ���D�!X��0�2�$λ�\sܱ�����!9=k3��qa�-W
8�{/2SSh
E�����+:a_z����z�qQ�n�Ą�J_HNؐ�a7�q��X��p����$KͶd���X�ϣ�<b�>�m�\�RM*aiGzU����0`0�r�A�5k�<y�0�U��d��b#@z#,�a�e���)��T5�p2�����Ѽ��2���жA�kY=�(��o�.�A���ENn�`�lͬ��
�Li�r�xu������*��@�>�.`&�D*����Y����x�l��]8���Q.�Кh��%т��#����Q��jkB��H�v#GQ\�+���j��n�E59����7V�+MGW,���l�,9�y��o>gA�\N�:Y��l�'cUU+V�g�|3pNf�(�荧<�p���mܲ.Lȏh+7�k�-R��ɹ�:6k���ڴ�	166,&�.J �������/�;�yο�l8�4����\��F�	W]H��@��"�&�`6�1��W���/�ƿ��]��T�(�7u�#�ف�B&\�r=h��,��၀��˂��ý߿���o�m���ӏ��Q��Rԛ�g�.��R��m�"I�SO?�ã���n4�v��+a������x���U��������#�`�_K��t���')��8¥��@�A]������(���I�f�����vX*�9�+qkZuX�*�;f���He�T�+ި3�ki�#7�+��T��c�e���ؿ���?��#G�e֞�CN�ց`Hilq�i�����.�w29�(۫�j&\
�)P&�qN�B�6�FP�����4��k\O+/ $G7Os�t�k����	������ L߻�ϰP�:"N�v�&�/����*d���N�D8W�77�痿���X>1�F,�Y�A��ζ��0;#xۦ3�Ӕ@�$hr�`��&���v���`��qY��QM̯��%��	¨���)��z�&"��ZF��Y��*Ԯ �rE�]��w���	�Ǧ��8T����C����LG�Y�b����4�j�	LAe:�EJMW�Eu����x�RC�dML"����c>���e��	s�U�vt`~r������!PM7?�xl7��8�mMX�
%�B���1�|:� O�_ݍ�+Vb�102:�C�F��� �N�j�L���<a�׬!@�(eERI9�Hȧ}�Lj���:ٰZ��
ª0&�jp��ʠ"9����HV���M��4I�Z`��}�y��t���|fʍ�$��Ɗ'�X9z#�����4[x��J�z�R��U���ć����x�.S"E��T	�e����V	�:l3]@�*a65'|�ׅ�|a�[��?����g����	D�a���u�����]w�y �+z��D:ۑ-Ď���#Ru!D�WV����q�,�������n+H����l󈹶�TOS\j���o$�hq}��!�p�`�=�db����?'�#��ʢp_�RIi�^.��E �x��� 0��U%�@�S�|]��z�ԯ�137-	O��F�[�Oş\z!�{�-����w@��Y����%Dm�Q�B��WQ([b�cx��h`A�����?j�O*aL�:�zH�1M.��KWq�JAX���e�8=�g{Ma7�r��<���c��%Ri��g�V���C4�&Jy-)��Lep���v���DgO?����q�g��.@s<�|�U(��I�:&_��ۓt^���(@�`]��R��ao��<��?K).�R�$��G� ��+B�uQ���b�`ú�����������k&���cr�����"Uv;|�����e|��������^�z�-r�=#ʸ��V�(��5�ʘZêmO~�\Gk�g�p�v^����B�w�;z�I_c�4�Q�M�9����pʿQ?_1�A�q�}�I�$F�TxcKT�Y��k��������0��?��2i۶�����m>��k��eÓ�hI��R��"�O#��u�l��v���^̡����]C8�I�#������Q�\h�!�:$u��ة��Q.�F*��#��}��.�՚l�?��aW-����w�Ů�
v��"p#k�2�"Si,�3��3��gD��&؎4�t�r��,f3�2��GK�sSp��hŐ��~3ʖ�v͊h0mݺ]�}jB�n�Z
�1`�S��8n�Z���*{8���\�W_�>������&x�q��Y�UG���R� -�Z��D$�X$.��f����8<2����8RS3B���=׻x�Qݞ�c�@h8������*����Aϒ>�EE[�\��,<��5>��v<�!����A�,��Y� c��r}���m�`|�C;+H#��J֊�Ց���R�'_T��_Q�v�w
"�ha*�.~n	&��4Tq���R]��Ƚ�ε芨H�3-v���g�G��`��u�-p�,N21������]Ll�h��e}Τ�U�152�~��˸��Kq�i��*��hoG&�y���g���-V�g`��� �тt.�j��j��'��:z���s��d|H�oP�C(����n��<�5�(}B�����"'�I�!TiU-�^�Cڐ>��������	��|z�RY�{M�S�=�Ŕn�;��u�ϯ\|�V纑�ť�+�f������x`Q� &�'0;=&��+�;q�E�ayw;>��۰qәx��>(�Vk(s���xQ��H��"0:����aݱ+�
�mُo�A�E�`��g߲��F#���	M�.�+�A�C��&�an����ho�������O=&v;m-m"�&g.�
���o&_�G?�iC.o�`������+/����]x��®U�+��ֶ �A�]�W>(M��`�Y#�K���v�A�PE���$�R��Y=V�%��'��!���75#9�D0S:�,y8W����n�I�R�<oN�*r;$���2������=���sv���xF����I����Uu�@(�$N%���]�l	.��B��}䢍��#a""N�Ӟ���nI:��%ɁS!S�w\:����;��)�Eָ749_��I�v� |��������}��u0��)������H����n����a���?�~���/{�o5��e?���<�[l��$NZՊ�>HM"�vUQ)fQ��E���Qr�RL׋�����h.�X��Y�t�	��܍���Ϭ��grZj����L��H��=x|a��P߂���8\a�T9�&�B
R��]-&�K
�Ʃ�P4$0+1[I�4j�2�E�079-􉬚&�{�P�Օ�7}e,�-�k&Ab�F�t#��yv��ɡ1�
<��}X�a��~�i��;�D�-=}�[�T*ri3�
`G��1�O���� �l]�yx�d��E�j�Rm����zM�qb��\�&ދ�F~L�3�B~d����`���h�C9S�Q�����,�J�て�F�Jqa�\��%)��:�����`�!p�Pd�.�i����${�w˖)<;
�F�##����CiV��$� (&:��Io�S|[�3Ԑֆ��/J�ti�8��u�jR��0���SIqH�.�������C^ly]����=$�E�GM`�t\8���:�K�5{�%��=��nn�U�E�\Tk�,�bN�����p���b|tM-�x�}|�_�g�=���<B}�Xs�q"<1=#��f�o�B����*�7�{��-_�=+��jV��"�M�\�<��ZZ�d]�0A`"�����Eتr�T E	ߪ��/ۅJI��F�����u(��"V�ydH������p��ѵ�W�F��Z�Z�ݑ	=r{,Uis�
��Lp�%�����;H۷����8">���.E�c���.N=�<\z�5"I�5��罏DB����dZ�Ӭ�p����b`p�yzn��; �R].i���۰l�Z���K5�:[f~�R�E�0�!������A{GTl��^���S�� R�����ǚu�17���ب|���Fp�]�""�!�W���N:�x|�k_ƻo�S�K9X��$�`8O`�x��&�'��h r˴�����@�⣿j ���:Q���8�ʩ
� /l��I-�t�Ol���f$6q?�>IW@e�H��/��1��T\08ްzR���|p�)K��Ylo�FO�2���'P\�l	���
���O�ߦǫx����Y�3�����I�:��^w��P�l��LG�.��J��v���9�]�E�td%\�-�|���+ZG���}�9	^#�֩�������o �ˆa��@ؿ��ԕ>���5#�L���yx��|�{2ظ�W���I4�i��A1;/=� �}��R�j5�)uŃRO�� hݔPVW �Sf|(�2��H�IP'��^�f�0�ʡ��G&��{~�����2e�*��+v�j�8�)}��D$��rap���g �K�J�R�V�}��^�{��` a&�R8�ۢ�ǆ�J%�����`�����&.y���Ξn���G�.�W�!7�D,q�%�U[4]ɣ�#Ϯ*�⪂`�d�E�ǫ紽�͉M/m<��LyU���QuK�u���k��,+!4�e�	�'��Ɩm/�*v�p����ݨ����B{��w����hqڭ��O�!}|/��i�!��?��/�{���.������l���ۇ��'���jYڣ�~�8wE��=A?
�
,��H�@�\^�Oy]�Zl���� ���tr�m@�/W܊%K1;6-�'�Jb����u�D@U�D3��=���q~��J�R����>`��)��y��n���X�=�@�/�d�E��BѨ�hXH�s�O�G'�oEe*�������'�����Vn&�ǟ|�q���� ��V"�ъ�tZ�ﬢ	#]�MUo0ٺG\a����\�f�M�[-��.���y�hUBy�LNxNԻ"��v/���s33�G���U��@�˭<:���Qe����dd}��I����%gS�;e�r���]O�Qn����1!�㵧81}TYqڀ�d����H��	#�xH��97=����^����f5���GW_��������l2%�0��LHX�?8<"m�kWc.��JJ,������_��g	�[�PK{��km�a
Vj�x��L�)C(���Л��41����m�4I!�RC��؆��^�߳��@ww���d����.s��8}��­��C�&��H��1��w���8�������7��V)�Q@�\">/�2e�ն�Z|تZ���ev���������]��K)��"��
��ȩ��9����
Je�&�q_y��p����SO?.UY^?vnD�K�g��lv9H�6i5�����f�Na~���&�ݱ�qD#MX2�ZT�&g5l�ڵ��+P��(3��T¼�ǩ�{�9�*kJM_�+��;�Ts�t[��w$q`���|�L�: L�6+܋;,,�.��osěu,;�J�PIs<u�,���}Q�U��Grpm��-��x^2�ذx�`���U	��˽O^��c[����2N�lsk�����⭧��Y',��Gw�W5�Z�by5^�~9���,����h�X���9c L:aMY�H��ĝ�m4�W���B�PF�w7��_���=��6 Q��y=��5S{��#Aa��e�<��zz�����Q�&�d�;�H�F:���D ��#���&�e.?ۭ�́1߿��B�0�z�1����Z�/��������D*�2W��Qn7+4l�Zl5x���$C7)�]�!Ƭ?_D�@s�	��9����03BHML��-�(WQ�U���a��+�ig�˨ar�0�Di>��Cc8v���A��J$I����P{Gff�ؽk��UNNq0�/]�B>�o_|A�1�+ll-pʓb۶m� ����D $��UV,�.!�s���I_�	��2L!������/(��Q�y��U�����+�Ė-[��󿕑���1��Cr�h)��]�)*1�&�uA��6��kn�TTؚ�*�>x]hc��)��'��fttwȐ���y	�<����2��2�(�5��j�07=��p�\�7���k�E���*g)���k�w���܁����Z�V���9�$�U�]�[�&�?�IKi��m��eب��0�%ªy�q'a��>��ڻw?�[[��E��X��XK#�"�*qg�b�A^��O�XL��8�/���[*�yVM!���br��#�0�V�:Z�_�>[�$D�=�qQ�A4yL.��:C�C�ḺX��]A>�*F{,�&�W_|>N\����]��*�?���,]]="���`:�AKG��;�@$����������?�c����?���'D���X��]���ئ�Vi�z�j�r�ݵ�p>�!��@%�;��6,[ֆB�D4����82�y:�������-Jpl:��۷����/�)�!�X@FS�fg��܄������{E(�,��2Ma_��g�����Δ�t����Sq��sgG�[Ƴζ;��Tv\jz/_4�����|��G��-�Q\uť��G�Ça�ޝ��/~�l6�R!'�+��n� e��.T��n�Iu���a\{]�=��OL���>oX@���`�������ᕩKJ�T���8$T����ͤKO��MsjU[q�?M���H�Oz�AO36�6���k��,5���4fC �S� ��6�#�qG̉ú3&���8(G�0 a7��o*6dہ���?~l��
F|	�n;�zeǬhF��睈SVv \� ��<�[�R>���
�K���V�h��*A��jc)&���#����".Hf�l#����x	tH`�aۢRC�Y>�bk6J5�P���;-�[�u7����(U̅VZ%�e�ג*��a�3X>����2I��ʘ4EK�<n|��F+����?g�)�PSH��(�J��n��O�aO��6�r����6<6��tR|.�*��j��i�a�}���S�9�HГ���)�31L��(��h�ı���cc�y"�`�^�"73���c�{BÇ'�l[���nDb!<��\��#�avd�hBl���	��S����DB��(eB@�w�p@�a4���GSK3֯_�����>��u�d�o���T�D���8{$�z�-T��S5�DOkN;�4��}p?~��YcQ����-��ݥ����΀�f�Zlܸ�s�8p`������Y�:a`��ސ��
\j��_�b� |�o�*��:$�*+
窀�j%+�o�M��҆d�'gg���f@P861&� �?4ڥJ;9B��2��]EmnRY��Z�v�i�����5@Q�bzb�d����׷���(���F�U��yݯ���w��=�$Ĕ���T�V�����Ҋ��a�߻_*`R-�f\�+�2�x�ч�ͲqxtD*2aX*���!
�\Jwg���=A15����$^��`K� ���G�lX�]��*���R�v��"��b1��`�Ф�:A���C��7�	��AKk+���I�F�]͂נ����|]�EzY�ݝH�Lc�kۑ�{��q�o?�>tP�}h/���m=��U�Q2}:VA�3y��m]]h��B(�͖�ۋ'{w�� �ވ�:8�Ű��s121)z~l_vv��g�F�?�`( �,�<����o���S�%4ǃ����ʗo���8�.]&+&3�!���ˤ�����;�FKs�p��e����/�3.��\w�U��X)R�۔�+��VU�g���Ρ���t��� l1iq*.7K�%Kxm���Q����(B�U��l�3�q0�{ԧ��E���M��g?-ٴ�{�'p��~���z�Z#��ms~6N�KUU󭜩[m�M�mF��%=k}^�NL���
�E���X�W�ĵ�^�x���9�j*�{^�#uҨ@5Դ�L����-HZ8P/�v�n��=Z���Ўt*\�1���@Ob�    IDAT�0�,1�[���.�6�0%4�~�Q*aa?��������]̓$�z(VkN��U��U��������Z�+�!H�dY��@,�*-�85���D�MyJjХʜ
q�aF�����i}$U�`+��I��
�w�ys�������V����ᑗ�a�lc�T�eU))�#��deQ�`h�� �xv�;r*=)�,��:s��J�2\Dl1(�>�\�"��|�\Q�
z���L��)�BToM�a����V4��v�t�R�jy�����`'�r2����I��Yz�pb��*_)�*d�X�U�b��ϦQ.�����3�S2�C [)�h�5��-b������Xٳ��+	���N�t&Ʀ�1<��#$���b(dMD�a���R�dRbl�hn��l
�㓢H��(<���R�=��Ԍ�.��|CCC�g٬�T)J�U�9=>��!�a��������썛䀛J&Q��sh��Y���DP�*�qVH�#��=r8��M8����H�U0�42��I�䷰�)EG��ؐ���6�9TC�[��5[�H��S��,�zq*SU��^�2[�cWWV�Z!������̟/�Bak��Jӥ���H��u���c]�R|}7b�:[[�Q�f��҆��<��_�g���C�9XA� [W�wă:'�8�P��S��e9<Aj`� ��WV�8�eM�m����\Œ���go�F�EK�4l'(���I���6E5ɹY�� (@׿q"�����r�)l�e,�Y��;�#��XU9f�3�C��5�/bݺu�2��c�Y���A<���x����{$9�d3[�?�ȁ���b��E��)��F"Ajz��q��h�]��3�܂K��O�\v����&�m7"�f�]>���q�bMR}ljnE�r1�(�S����
�����V݈&�r��g2�x�&�^<0<$�[�P�V<iQE�^V�sS�e����@&ǧ��ӁC`ߞ�xm�+X�fN>�d��޳O�kY͡����8��gؽ�T���{�D�_��q����ށR��.�z�T�ru�hȵt:U1��ؗ���)(4=�'�͘�JXP� �R?x6��**e��>(iĸ�`���%�ߨ�M��_�W<���x���b�ݘ��=O �$��V"qr�	ܠ�.->Gӎ�א ��J%, o�ӽ��Ue�]w��������aq7a��B�
�9"��T.�z�{�/�
z�Es��`��@{�ʰ���-V�[4��rڡ�8�AlU�y'�)Qꤶ�C�آ|#2����ߋ�l��m3���Fm;��>}�O��򙂫���ǨSuǮJ���{�:'.o��8��a�c[�(�e�ځ��9�ju͊x�X0����.⦞����|���1
��%�EOɖ�)�����Ŋ��<�y�����-�0�/b�v!os�{e���_���abB�3$�&i� }Ɋ%H�fE*�X��!��"��"�����
����L��(�yǰ�,��Ȳ�azL��9��T�E��#� ���oY/�1���mڨ�k8���<؅�rs����s��%i=3���ǥ�W��D�Sw�jU@L,F!�U�� ���U^n�yٟ��.C-_������m<�<�ԣxu�Kp{���ҋ��VʑG�W�(с��KB,G(D�����	�e�@�6%���XX�''�D;���=�kʠɀ���o	�=�/Aݍ��ZZ���6���,<���}>M� ֔�`f�l��`�����3X�g��(�<X�v.��mصw�h �'��I'��D�"��ԡ㽗�]x���rbQ'r�T�N|V��z/ٴ��p"W�����?���TjEtw*��5s���a��ۅ���	�-Y�!Oi�P�$��8����<��3r_N8��ś`T��hj���Q�:�T��g���|�1��"�~L_�z�as��SVC�I;O���r��i��r����E�Pۡ���.��m/o 6rX�I�<�5S 8�6�f�3#��3�gպj��s�-��mUQ3ͅ	9}4v8H�f��?ЋP8���^C�,�㏓)�CTN�0�t ��@�Z��c՝}"�ޫ#eC�X�}����Gy>�0��P�r*.�t� ͊Y�o6?/�K�}H%8��Ӱ|��]���r�	�Yc|����C�zw|���1����x�Q�1kH�4czj�����\r1~�󟋫�Y{S��1��g?F4��k�J-G�"I'�V��
F���I��|���/n���C�X"C,���\s�e���!��C��5Ð�۸��@�vDYt��o�f�� ,y�a�C���\?V��K��ii�SS���eFT�mY&������������8~�_wcxxXT���ZwZRC(�Z����1�PH*撔3����sֱ��"�F[H:A=�]����E"�N�xH��6���A~�9������I"+\��J�q&'��'�)�
u�5�A?Gl�"�`��$��O lA�bQ�`l�~��7��^yS��	�������ӧ��CM}T���ix�Y�2+s�z�_�
;3��m�mY���D0���kw~W̧��\��d���ʄ��� �N�x�ɦT�B�s{$Kd[��a¸�hu���R�?���L�����c*�C��EŭY	�c=�ƉE�.b;HMz�;NnAS����*$��Q.�-◪՝}"Q���h�"�
+�'�V�t*^���e�止X-�f/�f�f�����	=��H��b6=����E ��a`�,_�
��_�$M��Of�&g����Qs4.&�H�Y��2�ժ����<1Xo0�&��%Xy����߾�������UL(����c���Vb�������G.ˤ��E$S�BXP#�³�#�̫��b�ű|ʓ1 sp# �7 d��h�"���J�LX�! �٥��*������T��<��o ���L����.�u��x��e��m��F���c�-j��t��I'��뮿/���:����g�t��ƩK-5pB�U5p��SL,Tێ�0	�ҊW��Җ$�p������	�xK���t��a��e"r��Aѝ����FД�g��Gn��\�J��V���ذd��s�V�\!�ˊ����%8v=~��)�-kCSc�������4d��Ynx(ʪ+��l�8r"��#p"w�F�l����ZD��9�%o��dO?�z�����D��k�dy����m^Wːֿ$i,F��US�ͅj'|>�>��9��o�@{k��螾n���M�bjnZ����8�����*ԃ|� f<����1⹺h0�*$N0�̌M =9�& K[:�7w{�N&k	�Xr[S�����`���IJ�~ETݢ��=�)l��)����h�[��yr���e���E����wH��^����p2��w�qH���M�]w|U�ZE��R@�ͤ�.�n� y9�\��*%eʒ��=��䵦&�����-1N�s���?��}��!Ϗk���`��
��q����b���PG�~-@0G��	�Z4�g>�8u��( LIV�	²r�D"Ơʼ�ZЕ��w��7�+��%ڏ��v�?�Q��k1i�q���m*��]�-Hm�߬@�L�U3&�zS���	A����1�ߋ��;�K�J͂�c*a��DmG�}́ݶ� �`J(�J���i��AX�t��#M�V#7�R���O[ bGW�+��}�y����l�R����h	
�)k|ncU���`�w3�%c�����#	����������~�`'z�
]-L�eM��M�s�����6#7yq�!ܤRل'ǁ�	|���C���g����Ǒ�(��K�\�^�u-"�E���<�V�.�ټL�P� *R�h�Z%�h*��prŒLU�!)�.[j�S�G��xG�� �ш(>�IV��/�c�Q.V����-N�q�pb����ORm��2��9�!"f�@�Lc:9%���N�<Y@�DOO�����-�1=���ĴT���>nz�� F~��DWD�Z,c��\��5\X�l�|�Ww�@.����/��3ss�#\�Oc����]��G>�w]y��LD�n���+[�ò彘MN��&��{��/'E[��R;3S�|���hi�#�/brja�|>0�$ɗ�D�Pd��4�ja����<9>!�zj�����0|���xn�K�dM�v��{p	j�-=�8�����O��2F禥ZutA�Ζ5!��Šv'�.���163%����Tl<�K�0�c��&�A�J��VrD��� Xۢ��¶���.�ZU1o�ArgW�\�@(�=��addD�Cvub��5�W�Hr2������-`d�~tŚ�a�r���O>���U�kr�n~�	\|�0}��ͯ�eY�x'kE��E=%�]��V��\A�2�lT(�B">���F��k:P��ka;��7�O�d:�*VQ�K���O�Yg��R��{�>a��\��eKh�ݻW�y9lhI�(y	�>����G�a�g!:;U����R��T�z�
@`<=;�=�v��{�G@�trF@�$�.hV��5Iz��"�쐧]�^w ��$�F���p��a�sx�ʈ��(�L�]},����i��F8ԌH �'�X�	�\^�{)��j�l2�@���-_SyJ���DbC IE�� �oGg�V�N^�O��!t�5�,P�D���K�28�pR�؏�%�r��T��aDcM���EWG��g�Ie����p���۾�m�^�����Ȫ����]Z
���ab`-�FM�q7�{�D��cr��jL`��(�n��,�&�泎�6+a�����2٦�J�s��_�	/<��򡟡�ϊ;�c��RAr&c5��A��# d^�T�JJ<���"Tʊ�W�H�ӕ�W�-o9�}=�mCV���@U��Ry<pز���٩A��l�'��T��XF����bi�EB���rڟ�ĩǢ�}c��h��H�_�*��5��J�Sq��v���X�{# �^P�0�o*6e������w=�������}l	��Sȥ�a�I��n�j#NX�O)����+5�������/�H/���HuD/$=m�M��.�b�UU�j�X����HK����n��#�U�b�EM+�nHDf5�C��O��#σ��b	��4�=E��]��dHz�u�u ]�%��Z��k�w"��G��/���#za�p}=�Ԓs�B0onn@�qx�E�c ���R�y�YD�aD}Q9`����v��OՂd��^ۥ ,Myit���?\���_t!(]��+�������K�ijG{�V��%K��{bzR�*D�)9��l���_�������.�&�p�9�������UxY�)��7����O�-O��He���7��rI��v�3��K��d��R�_s.�A��̢�O�(g�z�%��@�}w��H�#�jJQ��������.�?��'x�͸�7b���163#��G�~�_|FЏC��21I �ɴ�}}r�ħ�0��@�#A H~��h��u�+ز}�V���&�u��S���5%�v��L�j�k&Br�W��Ctv�X�$㗀���ъ�e�2�Jk�L��{z�d�r��e�EXn
����B)����a��A��x��뤒vƹgb���h���SOcx|�H��������a��u��suW�&gf�AeT�$EEeDĀ�����b�u�uw�WY#(P2��<��<�s��]9���{�ٽ����?����{����y����wB����f�F&�A�4�$���[����V��k;Q0�P4��&�g�Ȣ���P�HY�Yk�될5K�Z7 Y��kp�EcfrZ~�xbY��\� R�v��G�_��0(�I�sYB�-W}�:!����*~����"��*����hfq��(��'��_�6�]bO����o��*�4EBO%s�ɳ�3,�1��(P��fqbvj�8,��Z�X2�p��VA�ՙ���׆��	d�%�}-��20[C1�N)�X�jE~Q 3xR,�U���?N�
���X������eGR��K�A'�\�u���Q���zY/��F����W�?��K�eȬq�5�Q1�"X�u���v���A&Gx��CQ������'��(���AN����U��fw�R�c)���R�Ź�p�T)�\@@��g���^{A�:���f�My8����8���&<IG*+��]Y�T.���&E����
K-lV��X<.��4�}dD!.���V���IQ�4�(�}��B�L[']6��A��`ԅ
�NI'��Q��z@�@�-�Cj-��x*����0���1�g)���f��V�pH��(ʟ��/E�u����<�̮;a
�E+P���4�-k=�d�p�gcS��J
�zI�"�0�ŉ�|�wC�a0YD��$Q��\�1(vm�āF���b.�%��bJ�{����Q�A ���#3崢�ie\"z��Z�4�����B�jl����n Af�����!� ��> ��3��8ٴ�4��E
DË���\е�T�������P7kQ���ce��:�1jk6�Eߺ^�F0:6�|��D<!�+�pyS-F�<�P��ُ`{+��	�9]����َ�p'�v��y*�Kx��GD�E���
�Z��Z��k6`bd�\��J|��kd�`ҙ�KD��?���Ż/>_��=�]�bv#]�Dn�:�_:V�ň�\��Y�����I�k#1%��]t
�5id�����BW��j3"W̋�<�L�O>���غ��˿ߍ�p�s�025-��ÃGqx�����2��PXN��J�億�zc�D?�*(�AO_� [��]N\��+�k�^I��Cd~��\�X��K׈���5�f^��+"5̒�LO�na��)$S:�j�҇��NX�ѨM����Cao��>,�3�5B�X�
��2Ƨ`���\EWG'BMM���m�m~ad
��4t0(�i���cȍX9��0h�Ф���G:A,_��G�wl�E��nh��p|Y�Y�����R�^�"f��a���:z��p��g��2;?���q8��
��&:'��e�Fȭ0)�Y#���H��T#?��3��R>���n��ט�bB*��`\�/��σJ�L��RN�?�[�etEEu1)h�U�,64{��YF���cnz��Ӱ��pLȧ2�S�4�$�֤�C���܎�B�ndR�m��RӢT�)����i�l'�Ĕ<2pį��x�r'�'�a�T������+���K�l(er�٭�U���/_N��*^�Sو��q�8E�FuZ����Gx���倔ɦ�r����E���*���`�q��}�0^��j|�	%�Z�v�d���t{�>��x(g.�$�s�PW��7�L�l�t�2��i3%oΠ���`���&��O�a3!�I��uUiD���{�����>� `'�y�z�`vR@y�:��$c_z�%�tr�P$�9��HM$���ک+9�4�jz��:��.���V��W� `|.�%�_����T�'�����Y��5�4����}0��a�����7o/i=-B��#��sX�a�67��\�0a��2�u�֙%6��1bt.�o���05���|�:�.�櫞��t��F������Div�	���H��J"�	�ŀK^h��n�N�>-�tBi��4����$E[�.7>Ybt5;V�N�-!ĲI�TɄ�=���	���m�h�@kskz{��ֆ�o���Ѐ,�d7��4�	R��?1� 8W�Cg�H5�����L��D[��{��XN������#��<�Q����O�f��j	����n�q8z� �Z"��m=w~�6�-�:��&p������`��84ԏD)�U�עw�jD���5�q������ې�(��C.��'���2�8�T�pÇ�&��D`6+cf�ز3N6O����
h戢x��PT�?YF.�'ۦYd̤y� �y�<W�ZO���7�b)��%�^����0�����b|Y�.c�%�y�0v܃��qa��sZl��jkH�G    IDATG�!�e%�Hr��9�N�F��ǄM=��3q�ygal|�3SXN$���14Y��ɊIE��\`X�%�u�Q��L�"V�cC�D���>^���9�`.ݑ=}ݰ8�������,V�Z��l
q�ժ
SZ�H�5��X�α:]���>��E	����tf���Dx]t;f�Td�����8����A~y	E�#�$~��d�dØWǡ��>�X_�l�&��%���E:�F!��^c@[�UF�̣�����{)�T6fAs%	�%c� `���6��H�U����uy�t]܂v�C^���.ɘ�-a�F��'S�4�FjF˒����F��p�Vry�n ����3�4a|t\�?�B^?r��D��=�����Q��z��B���(B�.�rz����o�~��� A�#����P'�{bU6d��O��<���%�&l?�4���ì,���ce��!^�4��J�K#]]��hV��E@@�a~�� �I�T*����Gػw��W�tB�cXȈrf��l��*�T�-#�E�)�x�Afq٪�%+d��dʽ�p�rT��J\���[�\:� �l��م,Vf���8Qy�����^�� �S�
5�$�_aT�����X�x'�014�T��f�+e�G�a�9�p�����.��&��/q���Q!��[�� �����}RU����0��'�R�&���O0]��wA�|����^� d3�lШ"T�[Y9��`vF���4��G4+[��&�����������j�pV2��hj��+A���G�<��0���h+"��&f�9|���j�S��jR�{䢤������h9u�Oh�v�����1���0@U
��RdmO��J�E�5/�I���2JFGJ��+�\ӯ\l�a�¬V�	s{]u���Tdt�^\±����]��+�_�O�p���:�&&075-���U}�57�I�)�{v�.��ZE/"�R)�I+���`�Nc��`��m� �� ��( ���~���rb��U��������\<��I���k��ہ��Gp�� �[Z�I�p��p��>�h��rY=|�Z�E�xsҵzV�DG'S�#0Wu��ŖQ��a1X��O�Ⱦ�����M���{D@�՘��\@*�.N%��܁X�Igˉ�/�2�T��?��J9*�2Z��6LF|��0e���f#��4f��Q��1�?�+7��݇06���K����N�G'����ݘY�����26v�T>��k0?5���	�H�u��`��a���p�<8���Q�E�����w���ǎ ��$�����cqX4a@��F6����):4����xE�X�ץ8�Z2�:H�
��`K]=�0�M�닏�J&lUb餀�T^	��㧗���ҝ���gG�^�������蔔�[u:��F��넶َ��ɠsQ�W�cK(����T/�����4^:xY�Y2�&֡(��
�4l�`��YU�O�GG�0=[�.��S�mś�JFG�ܘ�X�M�N�,���;)��bԑn�	�Qc.'�F�-Ʉ��anf��  ��[6Ke���\Z�npL�$��S�X�8ޣd����d�ɉ�T�����!�H�^. �qIy��a���F.�1�U�JM��rã3(��p{C(VX�mF��J-*<��i�,�Y�Ѣ1�w���:�W6�1 ��&a�e�<v��Z�r��ز~-�v+�:���UJ�2e �$�P�se��&@(Ք\;�ɵe���J� �Ê;��9ė"��T��4Q��P��EJ���vsS��j4e+l^N��{�\�#�M���;l}C��|^�4��d�5-"�$#K0�Kc�``-��:���W�y��4#pcd�b�9��2	IS���Q�,���&������6����H�|C�>'y,>;LEY����T����+.+=E�"�\���3���Py<U���S1j��	0��"NK�==э���NM��Ө	�����KD�::U0��1�5a�&�����9�sz�~��l�$`8��hN�|���_�}��g?�̫���u��Rr	.[_AGV4a�]~��0].�Y�B.#�9�݋�D���?A���(	�T:�Ș�9H�0'�r��)���޸cU��̲ ��Yq���'�$L /�.WPd~/@�Q7M����
�8����b5
������B����wF����$������������q��!\�u8e�)A�	��*|�ײ1�`�T
��K)W)B�"�Ga�M7݄pk#�Zv���=��7O9�l޼�6n�m�A"Ȁ�Wt���f��$��*��]~5kqx�~t��H=�R<*L��j���!LD�ѷv5֮ۀ��1�&��>���y)lZ��^�lc�/���.�{ޙ�(T$	ۊd�"l[e��;� +���%đ$�^�-���dn�u���=ɪHX��*`�qB4یR��8с����03>��N�o�x5�C�0�@�F�h����Q���_�n7c)��`Dtf��o������vb~zFm�����߃ǟ��^7����&�s��U��K���r3�dzjJq��H������c!u��,ɀS�jc��'��	]ɭ#�P:��������F�T������"�������\J��nҧH�?�y���T�(ZG�Q���@�����NZ(l&��jQ6T���3����M�F@�1]AH�ǹ+�`�T1�Lcx>�x����5:������$�Q��eT��Y1��.bvr�lQ��q�����aza.�Wj�8�q�H��yE�l�)�7�=��/��M��	60���L�	1f�e�t�q�/K��y�',��̴��x|n�2i�*;��T����T��c&jCE�Li����Yq��7�����=���UW���~�5+�|������Ԃ�=�,V���0I�~�"�f�6*1;��R랼n�q�F���$:bU�Yed#��G�4�*hy�]���L���>��v���@6����0�z�Y8�X-ND�q	=%�I��;-����>fs����V�N�caq�@FFF�J爛�V�=o�!a�^9J�?����K� jV��L2!c;�ˉHt����5y�d�Q@C#�Қ+2��
���8U90J�n�m��*��5 �Y���!r	�.[*L��Y����X��NN�N��S�h
 &�J%�O@ICSE���̦�֕W^)��7��%�'��X��@#S	zV&H*I��e\G�����Ca�Na��o>�=uB/}�#V~����q�� b�nM��9���i|ݸ>��bP����I�}����]i�������o�R5x�X���f�EGНң����`K��tnS�fvz�������N���y8.��ZUĖ�F�+���?Y��D��r#��vu5���H����.�>z�8���:2�
�Z=2���A;¤��q�p��D( �lab�	.���V��ia��S��>6�{�d׿烸�]a���H�㘙��>�~����Hy���}�!����6���f�N;���j:�K|��/ ��ǋ�?#�����{�EhM:��s�x�%�?���c��g+Vl^/�d���
��u�F̏L�P�ê�cdx˱(
�"
�*�^�&ѽj�hq��&1~h�}�3�����3�H����1<��/q��Β�'O¥���#JE������T#y�d}�~�k�h�ԑ
+����L+��q�S��D�q���G���ժ������%2"��o�x�]�A�}�;Q�k�!U��P0��ů�#����`	�]gD��G����9��"��( �)���6�9��G_��&0����u�&~��g����Q���� 15ٝ�I^�L解I�/`�V]@�u��N��"�ę�".��j�
<>�-͒���[X�ߗ���@3m-�d�H�0;l*���rC�h('�Ze��I�׻�(���]b؄ѦCA��B&�����(�t0뭰�u0frpT3�� `2!=��2�4P(��+�P�L�w\��ˀ=[G)��z+�&u����rI�)����XTذ���n\64�5��ue�-�YCv���ߗ�c�X�s�9�����]����2��l ]�		�,�m�ʺč�ϝ�G��/���& 1�0҆����a��݁{var��M�Z����^*u��݌���=��Q����~��ǡ3X�B�QF��a{,�N���+<�(�y�n�:��h�]a��x R�N�C�uZ�b���/�-]`�4��C����_FM��EBe��ې��'@�jԙ���;�@��������\�h�����c�a�ƍ���07���w�_��ļ�р��s��~\p�ŎW_�^Xj��n�HG�}^X�FI������#�Px����ݸ��;���pzQ��-�ϑ�r���G#��tw��^�bzzT@����<<�3Q�}#�(U�ZR�_<X��/5s|<�䣲�¢QH�p(�c�nJe*@���W_)k5tJ��_C�t<����Fƚ2�$3��7N�!���xZ=�����q�� �NUX���ԟ�};yl��{u=����Q�'F �Z�㗬�5�:�R���z$�56��F��d��!�Fsr����E@X�^w|�����=����"�El�؆��:Cu�S���gc� �,4���<r��'�V"�,�f#���fI^������О�.�0�BՈQ[���T�W�
�����\Q��F��8~��h�'��9L�/ �ͣ����Q���	�N�
�,�0a��0�f�,?M��,�]��Y5���	��x�7�c�I���] ��D:!���<���a��P!5�QY0tFm>,D����>�P��#C�<���z��X�i#V�_�{~u?fcԭF��%��a��g�H��)?5u-rKI>���/ǁ��逧-�H��w%�*����4������k��&ca�Q�5����^�z�)�v:����G>�C���F����s3i�B��fB�W�㚀��St>�\cM�0��=E�O�
�aB��Ts�L	�G�cv|v�w��?�2n��V�^�Y��.�X}6�O���M��܄T$��p"S3h�4a�ˋQ�ډ�c���1P4���f�����),W����4qMnش	C#�X�� ssb�%uO��J��F+�	�s~P[�L��u4�Ȕj2>��`���nFK[P�!�RA4M�{�d��y�>�B[L'�`�@��|�`��S�9�V��S�Rm��R7®WX�R����
[���&�����J��^g3���%�U1D�M�א�+6(���^՞9�����6Er(,$�05'Q*�V���"VWq�-d�J�7
F>Љ��W~�
C*���=)�4��k}�&�_�ܶ��X�z5v��!u:��Pjc��A2͌OX�b��40s��>����XL�
�'�Hս��E�1(2��%�ke􅃰V����|�^7�q�m_��B�T�Sr��N/R�<t:+�7����P���������<�禯P�L��i�1=P���qډ.S%���xSq��8������E��1Y�������5|��_@:d�x�M�R�(,���Ȍ�����z�E���OEGG+�����\~	�9���'?�
����4�������go�[Y#0��|�Pn��*�gj3��!��6�8��h`8�DjL�w�#n��F��98�V�|c.��
amN�E�50Y�"e�����a��0�GG{�L\@�Ť��Έ]E������U�fJ��N��mb�w�uc%��TV��"}��تNƫ4�{ww���}�<�t:)����f�l[1�9�Q��ϟ�y��/qo	j=Y�2a'�dK���za��	@vr�ncO�_Ƈ�H�{���0ѐ �_S���Z12����~���͡��6�d6�o0�W���u��~灿y���`4��"8���ڋU�&Tâ	�� ať,��e�w:�Z�i_4(�g٘"|U#��d
T��k�g5vd1nP�t�Ŗ�â`ެV��}��RN蓑8v����1Y�H$���'\j����5ad��
�H��	#�#�x2}�
�хz������n�A��<����Z���_$ ���\##x��ߣ�烞,B� +I;��E�M�[\�D���Omm��
�Ǹ�~<���HT��}х����{��c�p����@KG�Q�9X�&�V|��[P���s8�8;���Q���+ر�u�l�<u3�^e7x�w��M��y�%��E�Ke�)$q��V��ƹ�	�ۃjو��"
[��ĩdd)�����WޔF�Q9!����e4�ӡXTX�b+��fE4l�a�ڔ�&m	v�SC�����ڝ�Z�'�AIk�9�_��N'z�Pg+n���X�,a!������+�}�
c��J*��� ��8p� �q��0W�Z�z��v���<<���eӦΏ�s�=W6��R�����l:�d4��bL�Ȝ�Ҕ��!�w�,�P��Z�ȑAF}����r�?��@�T�ܴ�@3�ZÈ��H�R7�J��Ⴜb�J��+k���у��X��ՙ���ds�9����غ}��<r���4&3�� Le��-:��2��"4<�S�""���~��I���� +%�Z�fti��;4���Ia�<V������)��U�)镔��R�rU"N謃��E���G�o�l�dL���⺏������G$��	S����P�~������ǌ��"q�&��2�B���2N�0]�L!��\YGU,�i��k�c]Kw��y��y|�k����%��]�����R�q�vw�azf�E�F���0�J+�D_ޱ��˨Ȋ�Ğp����K��6H�<S�El�_[\6�d����/|���J�w� ����O�_��?���ss��v��*���,��C�M�0�vbl�:;\NFFY��͟���~�������n��4����s��+��5	ye�G
��|��V������67|�e�����R��/ގk�y��4�͎��xǗa�:������@˼H�*�D��r)�����W �^����ʥ�D�Y��qв�O+�>�,��h�v�cX2���P�E�]�$$lH�%�x.V���̆ ���alY�Zb0,�2Z<h��hF��L�`��cP��R�L�ǘn2R����L��ȓ����;O����0%���񧺗���4\�V�.U���4Fq4���x,�����)���<w�=A���*6ϵ~���~��`������#�ǰzE"�ob��fd�ֿ���xt%�RKД
�f$���A��,Br��Z++ԥr�c�6�xQ�)�t�)�o�*k�h+t�ԥۍN:�H�(��d�U��L,%�g_ĳoA
NLǒ������*:��2&�A.b�S�$�Tx���u�5�I�0��;���p�U���m*U��Q\z�Ű�JJ���C��ҫ���t�օnIe9���0o�`d�b	���gE��y~v^ʭY���̭�Gd>����^����A-�;�:�d�218���k���S��n�,J�҉����|���_���Gլ�!�Ŋ-��o�^���ٝ���p���o��"����]8��0̰Y���N�Z&�oTF�:��N�e�%w+�Q���J��0����ĕ�U�j��6:�x�(Z�F|	�XZ����a�sY[Z���/�^��)��	�Te\��$r`bb\Ƣ��[;��iF�����U<z�p@��=�ڳ�\L���ٰ
=�`22�х)L��hC�*l?�혙���䄔+s�&���ǖ�5����$�/K�%�X���B�\���Z�!,��!�I��~��<v�z�#H�����h�Oe	��*���r�<)��arrMM������߹����Qa���8�'��8�#7�s
[h���O]����t����z\�L	,��v6t1�5VYE�� I�����1Yn�Ԥ9j:��FL�=���c��:����'�v�*1P�M-�D��c(3�)��4F���    IDAT6��h���n�ĚU�����5����.�tJ2��i8<n8\Nlڰ�\=ڃa���K������F��1[��1<>&��)g�9،V������ݗ�m]�y,,��l����i�$o��ᷙ�������~����]|�+����ݍ<=:�h6	p�f�������/P�aWn D*Ý_�*��4�ADfsZ�'����EtK�Q��2NU��B���4�L������&m�r^��x-��w� �xc7��z�;��丝�ig���|ccSh	���ã�<�J5����?q��R?�y>�d!x$���^ډWw�^GÓ�3��Z��*���K�rئ#P��8P���Y�uz�v�q�=?ĚU��������9���$v�> �֌`��d�DF�`�o��b�a�T������F<ƐVF�V�����5h���/ċ/����477!�� ]����ܻ|��Z<pX�\�St��_X�W�;�]�{�9���*
�!u���R����ew
Xc%�[��N�N����Jt�ހ����l~xp�,VG�\c%[��V��%汚ҥ�2X* ��Nֶ�˕��L]��w��|�W�.[�	�jp��y�D"�@�MvO��Rb�ػ�C��I��+6��9atG��h��s�?�����~X�
��g&��TQ�N��� �.����a١��4Pȣ\�IP��f�ά�y~U2]�Ӂ��Eg�8"MF�2eT`25�q�6��� 4@˿�!I���aR���=�,$�ПuaQ�O�UVk����ۗva*��D4������Q��� L�Xt5a�A@XsWf
IѲ!Y�&Q��Y?�
����h��p��ģQ�Y��}W���3SSpX�ػ�<���V�Y�b��M젤��n1+|ꓟ����B�}ni�����~�u[7J����,>s�������D�iD���h[Ճ�G�b�P?z��]8}�)��7!����3O�=�8����P1�8�{��C�B��~I��p�D0r���d���=8�u��m���1?�B�j�
`�kJ�oD��*�Ԏp���U\WuE\�ѝ��#(N>�,'n^�'�����@�����; ������3/���v��r�f2JTFU[������ �X�n�����=�\�Q/��+�y��5~�嗰��A$�9��Ft�[�pw�cs( `��G%������8�3057��XL)�����������0�L�x饗���/c��Ű�Q;�;$�w~v�~61h�'��˸��1u_�����ʗ�����݌��)$Ri�_�~�{sS�YtQ�61��/,`���alr#�/#��	}T��(��Fٔt(����Ӫď4F�|�	�(�'�1��@YɆJd�Z�`����C���M�G�<��@X����;�.�S��>)��}<��(����'�B�?��O�����˘���k[[���<��H�K3��Q�ʵ�#�m�Nõ���;_ށ\2���1�^�V�������VS\m�Z�\^}>D�\^F�������tS�̎chjJj��A�YW��5=�����ￆ_�����]���C4�,E�/��<zV���䑈�ւ����&LN��}�f�*l9u��[x��!F�
`�(R4a�bR���<� J����,��J�y6�S���rV ��^'�[.2�p�����?�Ç�btd>��Ȃ���O�MF����RF`v֙�#�\���>�+��o�Y����!�͠���H�ǆ1::�X4)ڷl�9_ē�u`9��F��Tl2�%O�^��b��������>طk��J�?�i��Y֝ɕ�q��ڋ�@+v��#:M�l�
��;05=),X:��u�:��Q�F��*��r���h2g)�E[����z��e�EK�����@PqU��i����eY�	>yN�Zm���
9�/x�ȐE�>.�\��h
��w��#\�O� ��!3L6��h~?��Z�E}*��.�A@�C��Y;�1=M+bv���R+��W�Lj�?�]u���T�)�172�*ӧ2�$x8�8�=���R-��LIȪ��Ҟ|^~~x}M���`!L 5�"�aÃM�Oy�b���W�v,�����>��kVS����|�z[�!��]tֵ�`�.á� �
ԎPlo5�hk�Z%�U�CC�øfs�q�����L%_���2e3`�s�%��k�vwjo��G�����tc`��I�{>��D㱔�DO��F�i�FO�[A�Pg���R�3A|l��0J�����8}�Va�F���»��a3��
�193�_=p?�^��pԚ�Qx*)�Z�J}��n6c~1*�������O�@{~�B�u���G?��g��hoFSW<�f�:�gڜM�	v���\�Ɂakt|�Q�k�k����_B�u�ⷣs�Z�,��!��m�ʉK2�*����em�>c�,,.sX@j6E*����ť�Ut�R�5Q`N�"c��i�7��6[��M��F�K�Ol���V�0?* �^� �چ�=�^8py�i�h������Py49܍�z��l�9h�4�CW�:��iijx^z������*�r�s�J�CM�LK�uEW�edh��7�y�F)�N
X��%�/Њ��p3�QT��]���z���tV�f�m;n���S����������-�Cby.���mD|�	I�#��l�$	�&��t	=]+���08<�\���{w�\�֨�p��]ݸ�������~�ԝd-ut��
�:2aea<,�K�a�/V�h8�kFȟ(�U2���"���si9�v�Gw�A%W��j�ٛO�./^�Ë8��X�4�����V*Y,���blfF�s�^�b!�ˍo}����O������+c�&��^�����҅����xw��q�;ލu�+�ㅗ09:	�ծ���&a������r��2�lר��>�b:���a���T8L.�xX)���O�@�!ąm�Q�ݮ��f�ע�O�������ى���/���߆��r�j	�]�hn
���!�ESs+ҙ�$V�[�����߾�;�P��^#{��2�kh䎳jc�i%"E55�P-f�[^�m�����Z�̌�Rtq�C#x�wO���a�����L���RVX�xlc�3hnj�AoFw�J<����tt��g����.ގo�[��8.���k�/���YP(�N�<ަ���
����cn~:�82�N��ݘ��$@��dE"5���I\|�v��e#ҙe���K�T��-�E(؁@�]F�d�����+U�}^�N���3�f��|�J�B�Q��ǡ>Yy}��4ܐ�s�"	�����#��V�I�s�x�حv訛�#�\��Z�E�͝Lb����R}��O6���1'����\���'__ey�3�`���[�&�TR\�Z�<�9�L�R���#�J˸]��������:�ol������硂6F�`�$B��bQ���f�=0��5���$@��??�����$�N٬��g�Dv0�N����5'
3��JF��o~��r�bq21�������00U����?����nq�{�Ȣ$����Tq��f��x�i�p�e����^�X�\e�������b����Kjh�W��j>�V.N��2��F�(N%O\���=�:�ՐӔ�di��+�2��π�d&�X��Ə��P^��8{	�2����4��6~�:8��	�le�!�h�t�E�KbqN��1~�ݾd��ٛ?��\s��v>�_#]�e�]��kנZ*�n���(�y�i��^	ݓQ�VI�gOO������r����t���ď��)Z{;�h��.�W_���y'f1,����6�<.���`��v/��X�ڋ[��8��Fa��=-4&^۷�����U�Z��Ug�w�'L���0P�Ek��'��:�Fl^݁�N�  �n`fj�:O獞2��LӦp;�P�dztZ�����XN��EC?�;J��Q��ݔ�Z�Rl�6�@�+X�L`t�P�"�։���K��D��GI���bD� �uy8�FY���
z��kn���N����${�ı9Q�������
s�Ѻv�-~L'�i�J���<s�Z���E���s��H�F�m�Z����+V`�Xa����������?-�q��9��m��7�x-��؝����|M�Չ\
��)�ު^�"h��ӄz� �݉�hTF��|�7Ҋ`0sD�3�٧�%�2s�~��/Q�$�k�jĐG�V@Q_�Q� `���9V�L'��Eh�((o�[ۄ9�g�8r�l�n��0uhH@�Ck�y[��E�?��O�E]X���8��+5S�����Xx��u���ÀڎN���Ɓ=��K%e��v�K@�q�v`�1�@ �fn��f4�<x��020�&�O/j���&8�n��I�Z�c�ZH�!��cزjj�<\f;�	1_8����3LE���O�Ľ��T`3��p��w}�����؇�?u�V��+���u��H>� [�V���|	�h}+נo�*,Dcشi*�"y�i<��a�j����H���]e#3J��qt�2��&"gLI���S�ο܅��ފ��!�,���3��~��>����##�Jb��;0����+V#��"������~lذI2�`�I\u�eX��?�鏅e�v�{��}���C�H,��T�7XQ,(�i����"4ڊ$�� ���	~O��att5#_L`|d ��|\��w{���q��Q�)	�w�h&��P��f�+f,ɒ+��֌ޮ0�g���B��;���|n�C�䙹na�ʵ�^<tjj��N���,{�f@$�Zت�DU8�nm*�VN�)�0�.s�	[j5,'��Y:C	�Xr9�,�[��{l��H���0�* ��k*A�"a�L���|�f�2f�;�e���^��]�9��5�����5�`�ω�#�R���ߪV����7���b��A�E&�q�ٌ��(�	7K��-����E>�����w�C7[��A�&���#�����s�f2���{�c�?���@3����<��:6�����A_�7\s����-��I!�MI��J����ٴ�l���a*ݩn��*�\�t:}��\��5U��:,�2ja�F9���ș̙�`@�n�b�������0O�օ �N1E���lX�ž¨	�H����bVjHFgѿ� V��PIq���ť^�7v�!�+��\H��D�2�g8����� )�rAR������J�3ض���$iL�����è�(P��ނO�|�Z��u�Z��нa��'0�rfp���&�l���n��c��LȤSH�x�������FĥGۆUp��Io�jިL�z<p�S<�M}m8�2���1;��Jf�ܼ���c2K��g�y?]]\@��^���M��������'g"�jB��}�%ˬ7m��$F���^H�9܂��0�����pX�%�mРbb%����#X�_�MkA��	��ڀ[��	#c���N�3s���?~�t����遣+�E���!l��F�uDƧ��-Iiz�9��+Wc��UH��`.j�w�4����Epl�_�z\��GmO�^�)+�b�ΗP�򔮈�5�G�ɈiD���X��P;i7ۊ����]�����L��h2�7�3��	��&a�.�KFw4 ��W?CN[C�cBǖՈ�3�	+5�6�~�v����Q\S�yP5Y��A{_w��8�#���B��I�xm�f��a��0®&���ԷN�׽��h	���?��/��\6�P��hp��`��~�Z�\NL����ӋFldtM����\��#C�{\
ˮՠ5Ԋ=+��b��=����PU�幜09lX�y=�����Ò9`lU�����ͧ¦5"[B2��Mf`x �y��?����%�G�1ข��a|����̣������ddƮ�P��<��M�x��w��mơ�ǐ͕����߇��a͌���/��=��h�I���{ACS�`���!�D�-���Ț#v�-Flz-���W����=s3\V
̋�d�صg�K	@gg'��r��������	�5��ҩƐ˖E`n	@��`�u���~���aj�<�l���/~���aLO�#�#2��g-����TE�&�������	�5���p���3Ȅ��mf��p�֍x���uv�������g�-T09���R�	etF��j�ybz�d��KX���>'R�&Ƈ�|���+�(eﴻ`����,C�� lͪ��}��q����!�Dώ���5�Q�+��C��}��g�z�h�j�K^�`�YI�@�,�c/Ƣ�u�����\<q����z��K�Ep��#��A����dF�@��.�}�9�nk4������ĵ�{�?�Ϗ�ɿ�9_M�q�n��S�E�/7�|�4g�ת�h�׎�P|�%5+a��U9���lҭ�r�j���]���CLSUL���x��z��oݔ�8�:s��p;�pز��cX���uW_�&�,!�s�d�����ШFI�ڀ���|��LInV [���-�K��!S/�es �[���Z6�6<BU�0<��*���?�`͈�xB�B�yM��j�d#�l8IM��I��0R�.�Ka�,��"�s9<�6����:��"�r�&��L�՗_�o�Q/�h�~��D����j����1�!Y�w��-���BC@�+,71O��pXN�L�_,$�z�&����ciz~�!���{���oFd|����YLxm�����5�<V�8}#B]�@TS9�I?��ܖd�s��ga���ӂs�ޤ�3���KC��KɸضiI6٠�34��^4�8��E󥜐ؘ����ο�Oa��SW�vj_DA��"����!�ri4�[q��O㕣�(����I�[Q��P�c^�ѢW���$r���~����ҳ����052�J�"�s�����p���-
�醽+���	�}��=�穩Ԑ�-cin�BYFe��:�����܁�|�~�z��.T+93���:���+lG6n��������V�ۉ٩!�'��V(�Z7A�85�j��ȧ�%lܴ�P���py��'���/aǮ�qx������nݶ�֬�Ų)����[��ֳX��Ӱ��(��g$��8�AH�y�j����Ըe%X�Rm�ք�2p�F�C#�C���}GPJ�m�F��X��}�~ƹfө"Ѩ8�����w�)��j���2��l۸-� Vu��;�����(F&&141�|�*���Bn����hq������RK�05:�v�����[�F�����ގwm7~��#hom���<j�
�4�����c����@�aj5ɤ���a���p�q�Ǯ���y�whk[�/$�.�#���l��P��i�V���"�x��g�?�ji���?���n7�z��~���q�{�13@�dH�Q2`�0�%��[5���]��<>�����-Ls��:t�P/���'twwc���0?3+l��LMP�`xh.g2�,�{���8p���������w����8\u�{�`p�?�˯�j���O��|��Z��!P�-C�TP�u�8������N���-p�Lx���ƺU�0��t�v������c�2����Z"q1J�D>���&�H���R1�hdf�I�^�eRA��T�mA9�PrB������?���j4�.���h�3�H�	��k�LB ��~@ 7:1.�$G�lq SD�?�cs���H,�C^ Є�A��-��ľ}{���'z+�_	in����E�+��V7��6�ٹi%\U��Mp{��2^���tN����8ep����[�Qms��ɉiia���m1���b��U��]��jpn	"]R:y	��Z��~,Fd��V� 3���t0s���i��a���:������Y�F��s���q��]�z��/�v`��%�����jm	G.g	��ZV]��q�&4��I���*%C?�=��i���C!忍>,~�QǓ��:��N����n�20ԁS7���e��t���PnC���b�����~T��&FW9��    IDAT�$��歀B�hTFF�j�զtG�e�
��b|pT�X(�b%�T����t�)2�EriI@X(�$�?7��`8,�dR��8�Å7��ܼP�|��Y H����)��t"���^��'�`o�6�֬D�=��#���ScD��W������旖%^Ho1�&��J�X�h_ۇS�=KD��TFn�R�,�}�ˁw���c����y�l��T�
��9�Q���`4��IW)d�I-�+2���	_��,|tX*l��-��
 �xXz�����G+��x|B�0�	km�ݿx;�F�kCk��g���Z(��ˈdr|R ���l�[��n�ッб���3����, ��Fpm7̝��3��/�G�X��vj
ez}�8c18�&l�z.ֵu�k����?]]��T��5k����/G8�����f�V@��W_D">M�yIe1H��tNY�" ����[��\v�EFF'E�l��`�����������&�J��+��	��D��������z)�0�$iFI��qW������_ V�d0J?"�Q�V� [��
��.ḹH#���-!�i���5����	VV���57adtD@�/� =&`�.I2.���:�8k멸��K�2�?�ls&����8~��3����h�
[ɱ1��^�������rcrt]�������o�+�<rH6&�]ر+�s֭Y�7^݁-7���m�D��������x�w8:Џ2#6��պ��îCgȁ���qL� ���r����E�2˲9�]��$\�B�^|63Z#��I��Yg����><��3x���a5{�L�u��)5���o� F�;M6�Z��u�3��A��s��Z&	]���Oۄ/|�X�+"�JbϞ=��sy�p�<�NH@0��h�`v!��f�QZ�6��)^W]})���A�\�x��f���7����d����æ�0�ј�t��E,-����"R�͠`��� :�Z��D������_q!͞�5Z�cw�?�ӷ1���h<�/(�:D��U���%�=�,+ˬ�OΡ©�B�tC#ݠ���$TPd@Eg��q�A��HP�%#��Ρ:UN�N���ٟ��gw�˼���g�a]W_U}���	�~�u�{�k�t�0P� �I�.L��I'D$Ϙ:�?V�6E�gZr`��:�B
�� Z��_�+�5�.����g6��0�>�,[��a�C!a��v!�5���8�d���1������y�ɐ�Ig�R�*��]ssfffź��R��@�m�(���a�ۤʟ��J&l-mT�2a��=X�r�0������f���I�LLL
0���P�cjj--��*�gwD�~�~���۹�Z���,��/�������������l�|��-��	�9����a��3a�)��Y�Wa/�9���'�~}���+�/�Jvg���(��0+)XLet�6`fr�tR66�J���rl��ʊ0_�Յ�<X���{IQ'#��bcԪ&1�t)+���I�}:����5�A_��Z����:K���"���0�Zq0�@X�*���D_QafU���p��,�����F����#�%�2��7��=a`�O�vjƆG	�DgE����m9R����L�!K"�4�\Q*���^�B�R���x>>
��?H'3���(rCA�+��)Ќ��1DF��+:�v�
����#ƪ���r��z{+^z�%�7e,5��b�r�8��,"G+������Q��mé��	�M6;�����y8�EѰ�#��KC���pB�ۥMt�mGĈ��!�=�kdԦFu�>׍0a�_��"����PJ�v��{?�O��׿N
�q`g<S�XC0��M(B%Y�Җ��]* lv|R�dz������_�}��M6�v"����v��"��!�lZ�TT��39�yw�f<F'z}�X�ҍ��,�v� �MH����{�Bs�߼��Z���	ڏ����&<��}0��R��� P3�<9ML�����ȕ{e��\
�Ɂ={"_V�d�rL���3OaxbD�U�"$�"f'�kmkâe��w� ^x���h\ҍp%�'#mF1�?*j��,��D��&|�La�����"��t˔-}�h�k+)0Щ�hE��6�,�������d*.�Ћ�����G����T�n4x�h�x�n�*���4a�\�q�Y�H��m�b���� ���Ղ��6����W��-_�R6/�l�������7����w��T��������|�b�vv!�Є�@@��kU�����I�C�`B*�s���It\x�_ah�D�8�Ԋ{��|J�#:�[��J��6��o�qkV��� �ap�
�"Y���w❭�t5H���<��|� �ӦM�0���ð��u��
�˦��b������k��6���}�*�4�aT+�N	p�hi��3�j��XD�ՙ��k�����wݏ��8|�LR�E��/�'.�^x�9��ℓ������/���M�w�btlR�qs�U�
'�6��X[�[�Nl ^y�u(U���hmkD{�fsW\~	NٴN��R��t&�����x��o!�*#69�����v5��.������cA�e�TH#�M�P�lhv��>���^�L�٢�d֦�:;�e�v��# #�"�"-Y#�狘+��Y6�ONm�S�?>9!@�]���q��3	�&8�~hm�"��?�7kS��b���&��U���+�}�g��n�K~�ω`��{Y7>~ݦ��O�m���<�������K`Ž�����?��������xx��N���k�⩤�/|����s2��D�N�444���	�L��O:�j��r�o*;r,�}ǯ��^�>|����ͫ�1Ԕ7A1��(���2��� V�]O}g��,�8�QN�%e�J���-�u(p5i�u\t��X�PW欳,v�I�_�n��
tz�S5+q@�T	eՂHIſ�y7�aá���h�$�Hw��%��,�G�-���&H�2��(Ѩ�h9j7��M?,2U|NṐ�kg���(�R(IΜ��BQ�dg�ӑ�����!e��݃�P���|c�:8e�i1�f5�T�^�����`S'�y8�|�����(�P03=��XO>���������bߑ�tS��b*�
�h3#ch�,V47�3���E=�Be���0�Rc��UaF�2Vàb�����@S����h~O�.9J^`�� ��&!�L�Fz#I���*ߍlz�Rv�w=��>4cs�N/*�e���	�e���%���Ñ�CH���v6�#���i�6":D,��jM_���M7ӱ0�+N;�+�+a��.k��6N�VaF��2��sH����lĉ�V�s'�Z�R!�x,"�lV��h\�L:���F�����Z�}ػ�]DB�0��6l&U{	�N�{�HeK�5�`��uh�����<2�����1<��3�gR���݅�/-�ѱ1��4y�xn�k��D�P�(��
�&U3Yu�%N��N��ЖTuir���,���������\GF`��(�R$%-E�Ӌ�=�o�FxrNtVn�S������cr6��%Y��~�&,@"8��^qV��J�5���nr���_���ppl�|4��x��'X-��SWJ�#C��:&;͂���ޏ#���iP�ˡ1j��Y���n�f���m��͜P- M���C���6�q�����)-�CC��t�4�#)��#����6�[�[�2_]/Y	�I�ş�"��E"N/4�S k$�C�"���QTPC,�ƪ�k�9:=)��&��^#(�"�.��kף�'�r!��1$b1iS%S)i��H�N�z1��@Q����y��� I�2����	�ŀ��9����j�����n��̴��vK��z�*������r��>�y��}N�>w�6#�{}Xw�2���sh�ɬ�bD8���}�?��ҹ��x[��'��7�N=�$8]��1rh?�ĢA:��ؼ����55d�!��f��� ��܃���kĽ�{:ocK��7
��^���,C2��C�V�<�D".?#���VDP��w�d���R���s��LJ}�����x�3�5�V������$n�|��hZIݥ��]�w!���|����3��N��P�K��n�!��*�UO���N��g�z�9� ��\�§LLOa��U��&�5f�w)
3���?�*L�ޙh��>���v_Q6�|�Z�j0��dy��,%�(�S�T��F���/fh���H��Uq�ט��=j�Fࡻ���＀���2���v���z�&X̀�R�נ��k�D���Jw���5�TP6�0��ট߃ɚ���(PWc���aZ,/V8:�4 Ü0��L*���R ��30ڢ,�u��t�E&Z�a�L>/��������d)�����]2�O��X�<���l/p����E���������$���(&wDC;��p������F)���U��*@��c���d�%Dk9�!-�����7ۇ�	и/����n�y��YկE0rdW#�Ʈ�E���d�4l�mYwHց�~Q��������S��xy᳚b+6_7T0:����|~�ȓx��(�v/*����y��`�ٱt�j^�����}@ذ3��$ �\)
}�����}��!D8ۚ0p�d}fD*��1٬¢�q��!���)f���"i��=�O+���W?{�-Y���C⽴oߐ�0�B�Ї>$�f8���xxM~v��:R�9C/��$uW2Il4Rv�ӃT����A����P��09B:_���B:_��O>!~<��{`3p��砣�[, v��V-�G�\>��H�-����lv�>�!�Z�����8��_R�4@.W`��@UEtf��qV�i���ߤ��,.�k&�x�y�u�f���occ�ϋ�����K�}�^8<���*�,NX��j�~&�\�XB�C���km���>��М$H�����a�qǡ���g/�D�7)���V�����>��HB�Ί�]4�a�ڤ R���
Vy��a69��GM�9��#����MN4��r#�a�E��b��)<��r�{���{;�t5!�+��Y�J*q����Ccx��71�	�74�op@ 1�OӉNشI�4#�G���3xM��@1��Ȥ�xQ/�N������	�{q�e���	�t{wnl20�u$:(���ڵS�D��p۷���v���[hl����.8�_q�$��%k������^x��R �GI.�H'l\�_��6�𞚊���	O<�&������BKSN���lE/�xͧP��`�g~·cع{?��L�Ά%���	�7�;ؼe����(*9r/��G����N�$0�]�ײ�f�� EzZ��rMZ��>�,Q~L��F������ͅt2Y44�$~��vb��%�p҉�:������1�5'��u��~�&�@������h�7�E,o׿/~�f��.����٦�2V�������[&�k��1N�L]������[R�ߗ�XUk�MI„o�~�~�ݟ�˹����#���Yl�`"puy=�`�]g�}�ߔ0o4�u�/������Tܭ�|��R5�R�Ԕ$T�g^�����Y��5m+N+����i���s4Z�AUӃ���A7d�!<��
Ԫp�0V
�T|��+����f`�d�H��WQ6�1�)��?��5;���ĚB��`>�fQA]�D��W�M����Z�n�"V�J�0v��S"zl�7�p������%4+/�\6}ԆA�'��?,y�E�_lG_���D7�^bdu��&����TsdCa��@�͋NW �{�S?�b"���� Ff��u�6�9�f���0�ۥ=�B2�S6�$U[(8'~Lj9���`��8u��ה���M���#_�^�;�&�ue��i���Y�h-H���+?��T;���4�#��o�Z�6���ؔ=�$fa*rsk��/�����071�6
Z6L�Bh[�'����R�q4)Nl\|.���0sD<CSK3����CO��t5���Fxw"^�iE�ՂZ�<�Ϗ�-�b��T�y�#`�"`q㫟�|�)�ߥ��wr�DD��{.�:;�I&��D����cǛ���r!!��l�P@-�3Ó���s#S���}N:�4$�%��Ő/0��!�ʣO<.Y�lE���NCK[�LJ9��L��	�S�|��� oЬ!Ȅj��x/�]���e��`L�@>�\Iڏƒ�b*�ٱ	��|Mtwvk���2\�^Պu=K����1=<�h]J%b���^֏���_S3jj	��	�����߈�}�\dBQT�Ea1�ʯ�m����፝�нd �v̈́"QXk*>z��q�E�F�ZL�٢E��,��w���$J���\CeR�eҙI�0м� �J��tPl�_J"��4�`&�؛BFCI&)���p9��s���n�6}��<�2l'�lv�Iz@����&�o2Sl�����B�6�/�߸A���Q#f���`jl�T�Z-�~�4yp�G�����f�a>8��_{c�G�=Y�a�Ȩ8�wvv�ɩ�XT�g�j��I�Xb���wmلxt���	W_}�|b|��6��=�
~�˻111.�� ��'���mp;�'K�-����~���p�����M-f\���>,�@��1;�X�w������46:%�����߹�[��G7�f�V��\Sw��S<���p9�}�����+1�<��ܔ
�x�5�C�XҀ��]���e��^Zd��m�p��w}�k�V&˗-�)�7���R[��(:L!�5�	om �zT������M7,�	��M �LIf���%;���n���9�i��"�~�E�sGK��	�~niϜ��l�h	���K�h`�2��4���=Vc����$@���
�Bv���h2ٶ)l��>�*Lء\��;�����_�hY�@�Q�q~߀@�A!P��$LX�@s��V�V������ڛ�Ө�_U���m4.զ'꓄�,jE��0Kd�����h���~m.#,�P���vIŀ�ɉ�h���o2802��@#
�cLY&�>���ȉ��
_c�	�Ƞ$�)d+%y\R��r��d�R���j���Z��r-[O�񡸐�L�"_o��0[H�j L{]�u�E,��I�*4�2��ߥ��XmT���]��@|x=�f4t���]-�)d{
d�2&�s���Fe̗�p4��Vo���*+����}'��L<�|:�݌��#���dq���LOF����X���"ƘlQh#��h1���t0�}�`R׻��]�+"��S�az;Z��g�w�����Q����T�����5Vo� V�ۈу�1b|v�aK]�ppߐ��-+7�����߆���f�O��ua,8���,��rV���G�gC���ם�v2A��j��c�j@~.��L��Mf���8���$� 
፭o��74ZT�45�vprtn�n�	/��4�(ʿZ�����!�**�U6'A�	VWV�>+ƦfQ,�rXS���O�$���6ɹ\�?�ǅɹY���b��~�/Y��e�84;�-`f��A��U��$��5,�a���,�0(5���M��C6�	,]�M�Mg�sxச�]�H���%��fF���sI$�Y�i�&#
l��Y�;P�^���\C�,:����E6�?�Gf'ѵd1V,����v�Fز|>}�ň����B����Σ��ɭH�hdl���@�f��+�u[)�n5j^Gl#�����0Z͢�Ke9�����\N#J�\v+��կa5q��"���=�jū�lE�f�0o�Ã|���/Aݥb��u�j0�����O�Zȋ�M�c��8�E☜����	����0�!�JHv&Ewk ->4{]���@�ύG���^v�%\"��?<�� �+>�)�رs�	�ca�Aďk>����Ũ�������'�������V��{�Y���#F�-#���L�}�Ǣ�^����     IDAT�*�4~��[�͔�r�Q.�b��� _�ʵ��i�����[���˯�����v'�gB���2s��g���m���ڑ�s F�ݿ�9}�w�99=������d��	ВM4=���&�Y]�J��.��?�{��y͉)�������j����B�-[N&lakQ��E�g2O��i[�������B��,Z=QA�&g���CFt���R��ϡ��%���I�4�ެ�w�a*�6ޯ�媟��٣	Mv��NO�`S�,0,`R��]���M&�VEQ�V�s��˳����[���o�\�h�	B�k~}���0(I�T+i�9�*%�j�e�"��2J�f�@C�>���=Y�u�7hf�������4��t��.�!������x�U�K0�r0 /h�jF�`ǁ`���=H��	�XФ�0��|��g$f���^��� SE[G;��Sax����Ş.޼�2�)-.�Z8M�
@\��>�h��yx���˥��]��E���.���(�#;� �ڠR}���pH���D��Ќ�l��1t������]p���ۜp�
�m��V�Z�`<���y��F��Lf���P5���|���D_�Z)��ѽH$'�je�'al���YT8l��_O"V�␯j���EǜO��D�օ��>�Sg	�t��T�2�؎���PgW��}o�XKØOX{�O�a�9�{��$2X�ݏ�� y�q�{�0cHb�둈�PM�p��5�E��p5��R�(��|%SM|��n+�.#
>��|qҪ&��u�[ ,@ӿ��
md�c��L#`���ׂ�\s=>��6����h����b>��S��@�a�ۋ��n����I�\I4�-��$�'yML��e������'���;�@�T���u��SO��CN��wjŪ����ep�?~�� �#֮�D|����)m<a�j�x(�	��)V��ѯW2fN��j/���i���Kp��X��/I	Ó����,��w)L�<����Ɍ�sT�RŌd}2����]Bԛ;;�xq?�3�0�h�8p��Ӑ��KT��	��~������p45��-� 'c]�p|�|����׆��9a��?������
*`w��JM*&��Y��D�YE�V�2T� �3YZ��}r�5x=v�Cc�g3ِJD���H���
Z=������s:=�&sr��{�h�_���b�}��) �|�t9%#���5s�S�bE@Q6��(�mR)i���\���qؑIE�[��������	�V��7���o�o��v�܍K/�ǭY����o8�Cg஻~�p(-���������Y��b>��>s9.��B�{�`<����#8C�j�l0,E���.�tcaAN�t��#�h��jG,6�+����Z�S����*f	�~챧q�w��L� E��(�/3���ƦMk�o7�+M�������O��������T�r�sE�h�������a��և�tk&����&M�i[�i] �<�0>F�[�F�61�0�֤����@��Rg�t��ض@+T�����3V�������� ���45-�T4�<?eB�Z�xi��~��>�WF�&d����1ɍp�n	s�E��N�ݵ��d���(J�
i���Gc������Ƌ�F�*Z�I(�(���@-#�RˢZ̋��WVǩDN�CX�7hգ�B:
�Y�Ԥ�|-�ƒ��O��V*�ڪ�ࢩ�݊|&�E͍�����V����.�ł������8槜~G4&�H�k>a� �vju ����V��ID��������%��T�hkmaZ�vH֫�Be,�år��#1G5�z�k�-<Y�u�Po�iL�"S[����O�z�]N9,�j����$ײ���%�]���~TsE�۶]Ĥ{G#Y��>�g_{;F���,�ц5���W��ω��^XÇ�	V���y�M|jh�ԑY�
��Tx ѝ[��]VA�V`F�]ٴ��6/��6-}c����k�����8*ꠊ��s�\Ů��e�2MO��/x��j����|2��D�l~����u�OX�ݏ5��q��5h�������;�	0A�b7 ����c��0�f'�vY�d��L_��&V˕�59P�d0`�����_���)"�."_ȉ�.��9նf�qػg��$M^�Xy����6JXU�>k�׎�L=�Y�\�����u6:��k�
e�=8��FCPN~q���	'hɄ�v��}��[�y�Ak��>DKI8��p��"�'�%�	2`P��hm��E�g���j����P��Ⱦ!a^�����yc�6�I,>���Ɓ8�u;
�4Rd�VQ�pp���Jő!xP8�-ذ�8L>�\(�3O�S�I��$̢�PQ���>�8�
Y,Z���-����4�#>��11z.�C(&^s�\���>�%3�ep�%��b�-��BV�����a��:��)0c��r2����aa1�U/�aW�tؐ�k����&$�`nA!���j���5iR���Vъ��7(����f��&8]8�nDc����|3�&#e�\��K��3G��T�����3���ea�|.3�&>����%.��s>,�)?��-H���ĥ���.Ł������t��!Ɏt9}��R+E-�o���~��$�_�o�����'��l�הL�}�Ѳ�4;��˺���*�s��cN���@�����C`F0�_�V�F�EZ!�e:rlbK����]������M�S�_�?��(+��?�{�G��+li����ϫR`��á(<�4L;��>��_;��,��_Z҄&a��]v�NXnٲE��a����^c��]�J��̖ު����uF�2ޮ�0�)��ݣ i������{�1l�IϘ\x�P������0m�������Q���D�[��U�n��EQ�<�Wa����?}��/��|e�3��0z�0��0W#0�h��aQihX��l��D�,|.��P��/Tׅ�NC_Z5�}��}YH*}��4w�~�6&җ�/��l<N|�g�;��A��\��� �08�}t7��}�:��{/�J���/{�\\]0;,��L��
֮Y�����H�XsC#b�0�L݀���l`t��mh�ꄉ%'�ZQ�)�&�RM���f�����`�K肋e��lR�'�~^�֬�	k�ᑻ�Cj&$��6���?��{X>�[�x�p#cØ�k6��v*�<vF,�K�Ł�V��/\��P_�B!�#����w�r�p����B�X	�D^�,B!���,ؚ�ۨ�0��@��7
�B��c��3�y�+�$�o��T��/?	��
�Mkw>����t�GйdFg永�/��*~��SH˨t9hTeLǖ'���a/)���a��]H�H��X{�zlڋM��.$�%ĭ�L��9���($y�FMF/mTb9$F��7 5�ׯ�9�lay��f�dS�ѷ�}'ctdD"x�n;�ٔ���fL
�j��?�JPe�j̀"�q�&��p2��D*W!k&��������Q������7���E=x��?���=$I	&��j�|�-��]�%SҺ��������\Z��<>o=bE,�Q��X�-��8�g?��,ڛ[1��O�`���!��._Zlnt��D�_��d�0����wI2���ɸ����nN�|

�$:�M��W�^*�"���j������Kp~u*:/��+׭��uk�������'?v�����f	�rC����O�DCG7�f��`�6 �V�Y��zX�?�t$�l�:,�H�"�8-82zH��LZ�.RI���V����{gw7�8�X�L�>O;���"�Լ�h���r�����,F�lv��������԰:]���q`I�����ɀ�R�!�4U��֨�3��%��H�D6�*ّ�^q�7�Eima�JiG�gO�e/Kf�سg�dGnw�����ڎ ���	���D��G�A!_�E�{�5_ī�����.q�g���@2��LA��e�ה�0#N����;ȯɪMOOJ�l����п�L�����F��UX�.�Nчr�F��2���� x�������!�w��#E�Z@�FMJ!�ݚVJ
Q���
��cҹ�'}�^��Pf2H}oӴ[ڇ����5������������D���#���19�&d�@�"�7Gs�焨NX�����C`�^��^ =�����&����2$P���M����1�LЋn��_�g���αǨi��f�^Հoa���Ω]���=�:4��X����H'V�0�Q��æ�a�EaA}�p[X�*<v��x�^5���KB�ʢ\�8	�XI��ZA���-�����vzQdL.R���-��X>�E�4�2EhPU�;�g��w?�y�ô�0Q�O�0�����0>D�0V%�ݝ0��Ȫ%$�I��)Tk��n���p������U��ܹRE�qo�۱-��T�!"fa�
���8��Փ,\݆���h L&��ރv끪��~<7>�R4����E�O��+_��M�ؽm�\�ss�V��'ho�;Ј��<�m8�n/j���{q�E����t7�$�������r�:���e���mG<��Q�ʚf����G�p�[iSR��鴶<�1�����i�uzƙ)��,�F&x�>8�*nV�V��г���նs�������kx���ڝP�&DB��`M�b��_nF?M#g��s`/���3"���+��7�3��%��4�1��Gz5L�5ۑ�GېJ&�f��z;��0%Y�?}�k����K��jC4��3:J��3�kxj#s�x��{��H�&��Zˢ���`'���Ս��y	��t�ftu�Iv����m����ˌ�ի�â�>�^��lO��|�'?���B`Q�-�����-���L��&?	S��L����Y�R��8�N�"`$9X�b��d�ɖ����N�6�>��x��m�ih��,����N��'d��"���;*��a�ܸ��d�@o{;>p��pݧ�Fz.�\Jc�8+fq��@q����]��6>3�F#�/�՗^��CC����6��{n�f��G�ar8�t�`2*h���|� >xʩ0V���c(U<݀�P5W�«ϋ^������b�M����_���
���<F�C��9�p�sY�OLk�}2�3B��0���\P����b��"�/�@t�!��oQ�H+��%ӟS'��0^c�s+6��jj�Uʧ��qล}(�bPK9����ɏ������s"�·���)���ݗ�`v��!	�m���-_�;n�f�&��_�
��f%���iժ�hmi��F��7W=��J�����ʾ��ي�pH�;�{���������IY/��*Lfj�
d��+�n��FÒ���@,B<6����8֯Y�?����wbtlX3I�}Hv y?$�Ǩ��+,έv�Jښ��<;�̴BR:u�C����M1�P�t1��Z��p����/�b^�Kޯ�b�ڌ�8E���^ۗu}�nu��U�R�>�0��g��B��:[Ȗ�@Hכ-l'��pE�3ZҰ��5U�z�i�B�M�ۜ��up��ihLKP�p�N���'���8���oay�o
�M�Ԏ��r�Mo����l��keؐ��m��ciO.����)y��FJ���SwN��5�Q��1*�/|}*�=�A�BC�Z�ВdȈU��e%��ec'�6������8Uņ}�'q��ż�C1a����X�+�S�����l��#�T��J��|^������V�ȢO��807K�)�.2x�H���s�&#���Y�R�\�v_	�7L��|>t�WD�Cf��M�4�.j�hU���3��ΠN��ჩ����+���~K6V��ИiVh�#�fL��Ԇ���p������^iǐڿ��|]�~lX�\*���`�#�B>)ZN���J�Z�Da9-ʲ����T�z��t�Z�5&\�3��8�A�&���齈�fMcղ����!Z�l��Xs�I�%����;nAHMC�Z���s�;�mj��7��u����.@<�ko���#�qxj{�5�gw+~��٤0�<ȸn��&$�zP�g%�;6:��J���N����H������A�-�.���,�ǧ�}dd��jB"�ݮ�j�kA�Y�uh������{�6l@*�G�N�6�8�������4��6b��}�{O� F��l/��
���MXP��#��T9/�x�?iq�kE�;͠�*m�*׬���Ѧ�gK?pX�&hfض��������_)�@�?����8<�n`8��#����O�P��	���"���RX�f5�z��7|�r^��ۉ�i<���������~ѡ1����T,��8������ �G��14��];��+/`$8+�;۟�/d�X�|%���U8���0s��`g|Z_�8��m{��|S6�v�VcJ>��\�qX�'V3���5�<�4�93M!��D$7�����?��dM�.���W�p�y,����El1�;���0%\�4�&����\�wQ7��Z�\9���q��Y8�&�9�^�aӺUx�H��1?5����񹫯A?5<��mj
���/�dzxl��]��:����;��FP��'?�?��'X�|lv����V��_����ذv-����v��I�f5!�M��ۭ�������s�:`��p���t�`vF+��#I❷w�bu�)��|�l}�{�7 �������ǯ�/q+��*���b,{ph��M���J�P��d9�^�	@c����V���hۨi�LӉir�BQ#|�������@��z�)�aPɈg�t�_<��&ή����`�i�( �k>��I��u�zk�lO�����d8"�m���L�{[���h��'I�����"ʹ<��{[�<�u�?��¿�_��i�����F��ٿ)Mؘ��~z���ց�+��ե���ŦU0f�p��K�e��3�0�0Ԓ0�dҠJ����J��g�M;���_qA�u�Lc�P��f�MxlԖ.�5(VN���-Ȕ*0X�H���O��~�yO+���#
����5�ٌ�i(A?h���@��yP����QV�2]d�T�*Vp���xߺ�"�<03��_{QT��a��a7�5=T���bo����ɚ�L	���۶�@���!�?^�#��\��X��r�e�)D�搝O��郩�.�6�ah�!�3 m&T�x�� ��r���-]p�����q�g��CE	{�l��O=��������y���U�D�B���*U0Oj�(�j���r�9w|��D���.��B���G�և敦od<��P(L/�1��E,Dxf��V���۱r�)ذ��j�����Eغsn���h^��߉�����%�|-?Z�^�]s���D�Qa����77��ׅƞ#!��i�l�p켾
Q)���j�Z(!6���|f;�l�ƪ���A��N��E�l�Z|?f�C�y\�������N���7��#�p��/@*�đ}G03�bw����H����2�?=�l,�Ӎ���ݱ[�}�leK�4��<�����y`t[ѽ��J�rN�X�*���z�h�VE�'�[��`ƕA�3#��O� ���5+WI$��omE)��[q`��hq6b��׮G_/b��0�o��&^x�LL�ʵ�wv��W�D[c3�6Z�D@K�A���������^�D��QmO����x��uG�k��];�-pjf�C�Ʉ��4ր��V/]�Em�"柏%�,�qhr[�����1T,U��C�ώF��J	�-h���n�"����o��68B!8]-�Y�FV�&̸�kA����l��R��)�M�(k��`�;d���0GF� %8�T��& cۊ l6��U+���.��ĕ��6�?<N:���3����[�{�;���}O�(X�7��$��`h�0n��gȗ+h���7#êKE�ߏ��V���mM8��U��g?��脖Bb�`��~�#G��ڙ�יd'a�%����    IDAT��.xpp� �Ca+=n���������pz[�{h�
ԗy�=�|����[ob��!����~�Y��V)�?�C��?�=]�H$"�����s��	6�Mlj%�_��p���"y	�1����:j2]ɳ�����l����H���=�� �:�Q(R�_C��������9�"���%
:�g��M�<�)1n�a���~ԉ���Z�Y�9�Pk�ЗSo���i��{�k�M��\���~f��z��٬Ό-{�~/;�_��b��~�-���)&lBU�����w���<k���fSK�ilY�Cv��	�>�\Â�JV�fM@/�Ƀ�ca�;/�&RG��&��bXz�u-Ҿ��夅ֳ{�0̚�M�$�Át���Ɂ}�Fq����l�"쟋H��>ORA�0�Ӫ����Fd���5A���A��GA)b>�R+ï��q����<SSh���Co������R|^dwG�ȅ�S��/�s7D� 1M�����iˑ��>��*�l[|�F�aG�Q�PE6�����ƪ"-a#L�� �A�6�w�����"1�\�fj�.9�c��%�	�C6dfr�=�$�vN8�8�������R%- �z	���H�\��:9�u��ѩ&Dը|3_wz��i}�6�mi��(QwA,n����̅&��ՃT,����X��T�s�%p���8���뿄w�ǲM���h����x*Q�E_���N,]2�H"�D*��Q1�$Ȱ7��$K��$a�|;�E�7���Fmr� ;̪�H�#�b�`��A��G�h����4��������~�/�l�Ǒ�G����I5�y�i_����œţ%�4�q�)���>�[�vb�zD��<����"٠�.��V����>'Vo<^�X9N��UaH	��xq���EU�i�Z�@o�9���bnjV�oV��xk׮E����n����X�h1��8TڛX�t	.�����ؾg^z�e�����d�;�b�h3���W��@G/saY�l�pr��s�ǉ���#�|��1x}>y�==�>�e����!�K����4F��x}����Bg[;��0����2����#�$f�a��n�;�������*�j�4�#.9�lXs%���}�̤s8q˙Ȧy��q��f����j�`:4�݄|�L�S�W&[��ьH4��P\r4Y�=��	�/p��٤
E5��V[w'6l:	�J	o����(�H'B����༳>�Zƻo���[�b��m�� �G$I�y��Ó�s�����pyq��#�J�=8;�������;?��C�þ����sϠ�ч������%qw6sf=�Xƛ�����
�6��Ũ�h��֠ +�~�U�����f'�pzp�ŗI���_��O݂D*%CTM>)&�}�?���K��x�/���_|S�e�lh�?4����v��	��/iE{E�:ۧn�G
�d�X%a�8qk���c;����V�X���;G�OJ���`f<�6�]�c �`��\�;�=����^�I׆	���N�i���P��^�J�R��)�k�y���L@�g8��k��;�e�e�`0�d4���a#y�������&.��Z)�d+)��1�u�r�B�p����A�5k-��^�u��X�-Zݐ�D#:mY�����5�i3	���WP+k�w���-��[s�"��v�|����r��r{��qۃ�b�ֈ�D��ԝ� �oK&�43T}���V4B��]fc����C@�W����Ͽ�6*no���Į�i��ew�������P���Daw}�L.
=D\�����C_A���2!%�f5��#�F=���3�Z�*̋���S>� ��G�G����V�(;>����54��ӟ���~�B��c��\h�u���$b�y	�X���:�"����m^�]xp���g�(�gݸ���U[
u�E��ր
�8�Wʪ�]��iq��3T���^yyz��aé�Ƒ�S� ����낷+��%�0
"�����$�S��B^4{�]�kB+����j�ӧ��S̿ύ�z(��d�6���O�P��`3��0��UA���Eߩ��W�A��aG.�#�f�f;V,^��˖Kk����;Էp���֢�E���V��+�2�g�1��.���T�M6u΋z{�q�՞�T���S�t��촢jRQ14���Q�|�B���� ��㹐�f��/4��$��i��p�����0j�hl��؂+/�\�6���#���gppx��y�*U���ZFwg��ɸ�s�-�	�
l��Jy���C(T�;x 6�C��MV�ℕ�����p�XL��L� ��[�w`,8-�%\��/CGs�����7�7ۄ��'X��*^�<���P��e)!�L��Eͭ����:8�??�,~��s��+p�9�noD����*ZZ;%(��`>:�� �{� lEҬ48�5�ި��������! � +R��3y>��Dv��AA8�@ss#�*'�`]�y<p�/���m3��=x��'��s�I�û7n܈g�}?�������o|�=���j�F�d{Mtj�H7n��:���v�W�/��&��Ї095�o}�[b�pҦ�������^�U��/=��l^M~r�8k8�Y�t��:�0�AI��X���ǝ�h����&�þ���F��t:\�����=�֮^irO�{�����o�Oo�8&�r)�s�A<��"IĢ�g'4��H`����Ә'�L��+�:g=��RՌY�e�EU���"&�l?Rv�~�J�w����8��D#��(�_A�!�������\|�ĿQN�H��][p! �W����#��l�We�� l!+����� ����BQ��w�F����@XL�宇�����ˊ�{���V	��(N?e9�3����ρ�����MM�Xc�{�NTaGUqK�f�s?��eAʬ0���R��d��w� qC��"��E$�n����r�bx�[��$�����?���A�݆(�˚��΀Q�S=���[�vȂ&�����H�
���0V˰拰fs��X�? �a;��?��I�?V�]�ž�Q3�m�k�W���ާ�5�Q�*F��G�&�#�d��L�|$���,��#FGr���[V3���I{P��̪9�Ś���JR����ľt�X�ڃ����o��ك�HH�8��.��Z���؈�~�6������4��d{���X�(�v1}�R7�mע?�u��@TF��˦��4��	45�M�x��y�ۺp�nMaA�~��N:��7�H[+��cbv_���aj� ^+:��!U*�b$�0��$VF�0a��Ȝ�٪"����,�U�bNک�%�(#�F���f�Ń��/�E�ZVŖ��e2z.�C[�>�h�ha��$��C&�&�cwわ^�uk����^�h���Ŏ�|X3���I�8=�P���N�H5Mb��.2M��A���)f�� �;\�F�$-V��,LA���n#_o�-Eל(d$��'�'�P�S��Qv�&'vN'�h^���/��v����9,F��sa���g��ſC6��H��)$Xߵo/�:���i$24ȅ�2p���O㒏������ho��\�B�&?~x��84>�
'���[��فsN� �t���9 ��6(:�ѫ�f�d$���n�W���fǊ�%���6c�� 6�Z���Y�j*bq�i�[xg�n���Z�\E��c�WM�>�Gq׏n���A|��B�s�EN<�p��$�����KO������Cs��.�6��׊������X�
�IL���H� ��m@Km/
b��ڡ%"A������e(�,��7�`Ͳ<t�OP+րR㣇q�}�a�����O��| ;�mǇ?|�.K��/� ��"���{C��d�
�ٿ_���\�+?}9���.ff�p�ڵض��aڷo�[����Bg[ �}�p�U<���x�&(�<؛��e�,S!h��X%��k�hs!�,c�ʍ���06���>��#c��tyQ,T�%��; n���I@b!�jre�u�X��_�X8�l:���x���*�'��XԆ�8�I�X,.'�ƙ����X]cy辰=��d�n:F��+�2�`�J�$[�'�_���.Sa�0�0�j�L��(E�M����#�PX�_�����s��"���}��-M�,:
����m�>}��Sr�{���x� ��S�	����9��ȟ������s����p�m�v�O�aݲ#����_O%s&��,^]�ȕ�0pZ�d���EMah6�;8]�eTi���,+-����	8�i�Y�(�7j>b��F�TVI�D�H�����d��CG��G��{�0;�rk|�����'�23ɤ�@�HQAAT@��i�����P8�HS:��P��л�F��dz/��^>��Ύ#���]������̞�g���gݫ���9��|^iu�r�Ȇ45�D���*LF4�7@� �J#��"I�|)�F�J,K���&��d����3=�P�\+��%�T3Е��2ޠX�`�7�b�ɽr�q�,��2�J�u�[���]a8�pA+YA�TFl���a��)�7 �Qy:��Ak�h�ҁ8t�
jt�r|N<���Qй�R['"�B����>X�z��I�d��m�kK/�O��0��zdy(�,�އ�� ?���+��NҒRM@\]x�p[�X��2s&����� �����w߃���@�8jg��>5��9m(��x�pߚG��sW.���^R�)~&��JޙNt��tR���4�Ѧ! &��[�)�1<������F��R�Ĺg�%���v��rRf�YN���}V"L�U��R�� �	@a�wCC�m�&��f�C��mv� �|)/�V�E�4*�7�T���uBt����-���Ҫ������rbl �*+���SSsԻȢ;�8�$���pL2�,Ofs�9����"��o'�]ði�rb'ðd�\�`���A����m���l߳�� R�"tf�(�3��g�'��9�M�O#�����G��!�����x���0%r{>*����+��N�[7ȶY�b0h�݂��q<��Kx|�S`��ь֙?��u4f�֡��0M�[g?�Z�'�Z�<�����$��Q�����q����-X��L��+.���G��{*��t��:�x�b���`tlH�l��LN�`2:a�y�d�
���+�;G�mtG�J��p�㹖Ё��cl|RJ���^��hV��B�.;��������}�¢���|���ᅗ���*�����ї���S�ŷ~�����ϡ}nv�?(ND��C�Z[��]���;D/��@C��$�d<!f��wcNK3.��h��ۯ?�Z�	6��TV��|Ved�ȮeX�6�)��[0�Ob�' S�bˮC��5��rR\��He��4##�t���+�T�Hg&�����c�F$ �:�c)��?����E�ļ��zmMⱬ�S�*!��� тM��1�q�:pRϖ��O#R�,��L�cg��ph�*�>j9�]}4�F�*��'Ъ�0%�VY3yؖ��)�Su^V5^����IU��ʘU��L�j;	�7�}:�8��{e�������'}�tr��c�*��ք	�8���(&�;]iz��Wn���C��V�֢E�4���z��3H:q�%߆>��u@�2�p$�3��=����`�D��9�RFmJ��IM뾒蕩h�57S3y��P�\"�ᩉ�B.�aH�q	[w���?��-ۑ����%��p�C��/LS3k&R�"�0�J43�u��L��E�W�O���cg�WZ�H���=jL��-5J���z8~1��А�(C�+��CiyQ+�7=j�Hc�m�[��O�B<�jw�E�&C9����ۑ�1�p:r2���M��(I=�
S'9Y(tf�c`��)�TZ�sKE�V4C�R�Lz��x*u���fjòHg��:<bbX�l1������X(�\(�(V���T�� ���\!�S ����-E�|Y"/���/@:���("��zz19���Xg-|u�4��pZ$�v�`?�^�,jg����1��lB&�T�0�I޷<���̹�!M���"��J�GTd	Y���MD��{�����"�=YC
{��+:�H�bv
SჼP+E���M#�;{���{�&f͜���^�3������RX:�W��^�"���	5՘�`9�J����>�d�t"�MH �^D~Ȉ��兼�d�H JvJ�ELI�.U�ĩ���������.�\�fY%S��R�
0��J:>C/�,嶣��MF���>
1]���s�n�=���g�S�!UEa�:�jl��+�t~混c��=ص�C|��ϣ��{:`��=�����h������/H~!������=�Sr-�a���'��&��BK,Ē�q����{���$��ށA̞?�.Ɵ�^���nhM�B�56aEG�8�;xs�Xs�}��k.��c�C��+���t�ڡ~-��J��d���Hũn�#����;����H	��t��y�4���v���ID2I�Y����r.���^�b)���P�P�s�_{��CHf�R��˃�c�v한7Z8�ok_�P,�X"#�:k�����3[�I&M
��C��ի�d�lݼ�]�X<�W_�}��{���Q_ð�
��r��Tt$Sf6�d��ġ��Ak�b<���#N��9�l؁��� 2�2&AMt���~	}=��@Mm���$�kl��s/<���9��
����d`H�5�'�n/B���MZ�6TT�im�t)�T��U�+��#���BF�F���S$T����*{�1p�,�I0�?Qe�SNFE\��
�
V��Vݿ������#B�U ��� �k�t)��A���i�gU����'�_կ�j��?�
�?�%����2��Ŕ&�?'1(Ui���Wn���C_��<�T!�p� �|��Ж�ރ�/�&�!?�,tO��I���'pߚ'0��V���!3{�V&�3o�Rt��!(�7 !E�[J����L���FH0�"[=;�DF�II�\sY9��j�1�)��3�j����>���jފPS�H	�#��t�E��,��bDZ��� ��#�� �U�A8��
���bO@Ś�d
�l	�� ґ���صfgd�Ȉȅύ��7!R�1�̀��㕘�#TZ5jjk�J'��fh7n����S���u�֥�1��u6E���:��at��H���Atl62.��<��橵+��*3��0�V-��e�B�/�E�G�nۼ6���2b2Wt0ȩ�h
��R��V�|�4:�u�B%�Z��4M���X�k�#����'.O�y5\��f9�Q�����$u�왒t�D`��$���h�;㘐���JK�l�lQ�w�����2_����8 <^7Lz��j�y���;"O�0f��|BR�Siz��^�LdQ)�aҚ��k�����ĤT�n!���׿�u�vuuKP*]��TJ�#-vb����5��P��r���ק��?G5�F/�?�L�wq����z���\�¦�Yh_��v��,�{_�爙'f�ٌH4���!S(��Nb|pXw�Lr�N�Ǽ�64�Պv��`���t�X7��XB0-1a1���A�Y�	�����1�T�29�ik����:��n������#�z=�,[�9�ڱ�͒�m燢��p�k21{F<v'Ar*�Ø7���㢷*�����T�"�c#hq���~K��'�y ���	��޹hi�+���G�\�GC����*hOe
�԰���=k���F��#�S�蜫檣��d��x"%���^Av,Y���Ft����H�Y"G�Â|8�/�p,~q��0�x ���.�&aqX�>��[2�V�����Q�7k���C��Ȥ0NC�h�5�͍���K�z��D4�s�='��UG��Q��M�0�ׇ�m�p��.�V_ě/=���q    IDATZ�v��t��~�>S�H�B� h�*d�)	��*�=w��9���!�z���#{jw8Of�b�j��}��q��Zx�>i��f�0Z����e�U����ܳ�pp�hu*��9�3�Sr�|SR���po�r�S�,S �
Z$ύk1�~Z����l6��f�)�8��O
�s4lE�f��g����/#�5��2aՑdu�Xa|�.�K�C�L�cAN�W5aU�4�	�lH��M��P�Ӟ�tpV}�*S��H�0_"*��GET�*�|������:;]�X\>J�q�u�q��Ap`.<�L��AhI�"0��N�a���6��^Ō�EH��(��"ZEثTU]�JN�"F��d�V6-.A�d*�{
��p�0(�SL@I6
�n���M�-�asz$ހr5
���$�ec�B�xq���'�%H�P���Y�Z%#I����Tz��CO�J2U�nNҼE�*��u�"8<&�mZߍ%�t:z� k�3�H&M:"e�W

�	�F&���zd0�\ˑ�c����� �,K�ĵH=�?T�X�l@:#g�*L�"���d�(d��J���g�M6�l<��'����W�3�K�`s�01�/�F��se=�qnX6'��s8�؁\.�UFw&�����(ymRh^�
C0�Q�����f2�a�*�,�F#�ل��((�x�R� s؜r��m���mw#�� T.!�� ��Am�H�o2�o�w�a�0�NC�t��bϡ�d,��:�rS�lZ�Y�29>�^+j�Qv�v���<,V�0��}�����P��d 6@ɿ�J�l.�E2��� ����d�1�Υ�/��+.��J)�0��B���^�I֒�sd sp���p8l(T�e[PP�2�i��EF�>#�̛�!�d��6�gJfM��:�*v+�d���&�09���
{z�ǒ��`m^����;�4���~�x�X6��;��}��NU�o��#
u5�tN��d�F涷bv�,	�L��Z�=�tt,�|B�.u�s��%2�s����5��0��+�>
F�	���cuL2އJ��d5.��_�瘳F��c_ޗ�|Zh&����h���W_x�{�E���kXp�
�P��᰻��e�l%1]����Ǆ?��y��GS�,8>�x�ؾo��Nƽ�s����7�Ί�/�Be4��ko��iC��^+��=Ff	ayG+���2JNF���b�X�R@��v�O�����(g�����_����f@�C��f��c�u�\���b� �D���5�����Տ���u�q�_V�s�vd3��9qHrv@ى8�*tCs��ʚ7���?��Q�:e������e�!1�P{��oM#���i��.���f�\�p/�l>7�ӟ���u��%��qc��0��ὨR2B�cKIE��	d�^Ȓ��d���Gޛ�xO���=���橕u��ĉ'~+���-�3�U�B����?z!yo�:��x^Xu�X]ӵa�>E�h<͙��U���k:k% �cگ��)��2���*#W��������ΪU?_�ه<�+FT�D�ѿ�U��ڢ�}�>��y����F��8����|o���#=��g�Gj|6�C�yx�N�T�ƾ�>���;�zj�7z�W+�'��Z9MTk��⸚�Q}#���-)��+iU�$�������r�����)������*�X���e��|�a�ՠ��I��H����"�J�xYOZN٤�"[L�-Q����+�;؃��.�X0�7
C�䭅YF)X�&���Tt���R^Ɗ�r�\F:/����t�+��ac,��$�X�K�T&-'9��F-J���p��;L�E�j�������=��kF&���و�l��D8P��
"�.�|��'��"v�(
���F��(i�84<*�C�I�%���`s���С=r�Z;��1�LY��Z2ӡ�l)�h:-"�lQ�<���Z�>"3��e�ԗPa	�Ռh<��A�S�X1��T�K���L���N�������t>#��M���P��T�|5I�v���E#V"C��u�0����'�0;]SU!ʩ3��IbFc���J�RI��3g�9���E����1��Ȩ��CL�f�O1S@1�E9��Ek��.�^�[6$�� �0���ec�g�(Ӊ�ߑV�O����t�2�j�x
(d�b�������&A�X%���C�(�����1*k��B�Y�U��I����HdA���e]��&�M�ύL��h�VgA�BP��:�pȑ�����b���<�e��U����E���=S�E+.I�ܽ�ܫdfkj�h�Bx�^a���FG�$��b�I?lF+j<52#XǮF-�N:�派�G�Z%�m��;vH�9ǒơV����c��-�ޤF�RF� TUg#C���,j���׎������눅#�}���-GcC����A���尦�$��<�xZ�m6�=��1��?����*���M�]��'��V�s�G��4?�h�k`S�Z/��`q[��fX�@!���=;�A.��0٭hniA�����N��cR^�ē���Ftv����x���u���C4��nƖE��l!:)Ujܿu	��|<|3�����B�-@�!������!���A�Tf0��M.c<�ƧN8Ѥ
�mځ5O='��#W�Ċ���<��� �FC��f`r"
�ь�/��݆�^t��������f�I���dT4>%�zo����T���zE	"�mx_+��S| �/���K��:Ǥ�l	u��B(�Ivٲ%����P�gEVI�Пꐜ���*x�FOTG}������$蟾�Np��R�7j�?��M�����~_5�L	_�߀����@�H#*�n�Z�c�F��J�J�H��ǿ�;�'Q�y���nٴ}��Q�8�k�w�s&���a����n;���B߾=0� Β���ӊw?؂����i��M�RtO
��G�'6-���@���ݐ��%񻇁[���^tbd,�ǊF[OK����7�o.�l2 Ԅ574ʩ��޽2�\�x���	r$v��ꕘ�j�L&�p�u{�`�<t����;%پ��z�~�����k���W�	�y�Jp�T.�r�c�xꙵ�8m�S��?����K.B>�@�ۃ����[\�>
$l��c��W��\U��F���o�7g>��{l�Y�d1V/^���{a���r8�L�M&a��7/	�srb,���C0������c�h1j��P�Q�d( ��,�ۻw��fu!�͈р ��VؾP"!���׀�Q?ٲ��N�>��R
�A��As ��&/r��Y��^kD�:B��\N���Y��!,ik����<�tF�#q�����I�9�T~�Q!�Mb2��W�݉��I���bX�v¬S�n�"��#3�Q].W�M�df��C����z}(@��J�X�`9#Ya&���;=�����wRr���8�n'���lRj�A@&��Ia��kk`ՔQLFa����h��\/Z,4t��9VAg2���SA����D�q�a�a3�F�c�UA��Xl��}�)��S�+4�i09�$�J�OU+�c��"�Q���e�je`3�p�gN��lŦ��������#�b�!���!�k!���q1�t,\�e+�������`t`�w�B��F�2at�q�(;%k�
9�J{C�"�f�Gq�8t�SD-e,��S<�ı7��`�	��0Hz�	�DV�Ff��X8sn��/1�y@��C	��C0�YR竓1�^c�kE�1���!��Q��z6�|Wp�-��P�_�a�o�}�j!�+!0'��=̊!f�I֛��X*���R�bɐ�Z��}�KM�M��804 �잁~Y�7RWS�pЏ���6Ob�1�m�E5�{�$�~tl ���K�{Ι0��Ȥc�����.���s��X�p.�.FG{P.$a2�,Q����rs��.�k*C*[B��A{��X�x�o��_��U�����m;�㭷��y���0�](T��4hThn���?����x�/���G����V���R�my�T��ͬK���R���D(�\"��Jʯ��`�}r<H1_�قP<�3gɚ<<8��N;K-Fׯ�Y��WK6�ce��W%2ܻ���UGy����r����΀U�A��G�U����R94���0�5řT����/@7�[���>���8+6�	�TT�*��j�F�J�RtC���OV�����6n���֖:��N9��n���0�K(�#H��c�K����İu�&|���������Q.�8�2\��>���:�"�,}t�J��b!�+��Oʱ�*�C_
gR�ΫP�ǔ G3{Ŕ�U�;+@��Y5"�!'^�RD�Y�"�X�?w��K� uM�����ϟE�7��cCR�k�O�'@�Ն����M������C�̓R"��1NX�)���&b��D��a��^�|6+�#n�F�K��.��%0�B��>Ԡ�ق��y��a��m�Ȧ�2�jkkC2�MM9GI�l�^z�]<��k(���= V��^�\���[_���0���:�	�l&�G�<u::�Ȥ�غ��vϽ�4��@ *!�,nk��w�>�d]��ʠκ&��xܵ�ڊ���,&��q���kx�o���L��-hdSl�𝯞�|h�\���}M�h��i��d�PӒQ"0̡�W�͛�����S̬��l�`��+:���N�&�A>�����!��6�ז�,��h8���D���bY�)f~�N���X�xc(�R0����\��M��"	?B�,���F,WD,�C"���d�M����B�ωx8�ӆD2&6x���F :���+�*0�mHf
��H�5�&�5l7�xX���8r���8��:�2�<^6_��1F:pl�2�el?Ꟑ���v���e�K ?��1��:�}K����ᨢ�!�1ۥ�/G)S��d��H�Y�T<�B>%�P�>�q���r����oa˶�r_ۨw ���� ��O�̡Va��Y8�K_���ɱI�Xפ7c����:SHOו�����N������=�/��V#� �0�㟪h��d�q�O�s�.�*�b�G-��$��2�\0}�(�bk��w1<2����%�3��c�"haD!ϗj�No���E�,�Qɛ~�[�)$R9�R)��}�װ�@�\�r=̲�-�X��u���\$8�3���kg2�����˟��c��б�9T�OL`��M"� ��H�����?w	:��-;�b�j��IQ��mC,���|7����C���ԊPF���a�d5�Tr�B����i�F �5�H�ɊH8�Z���1ح6��vd
��hQ,i�m�Ȑ�������}��G��߅C]��]�����:�uޗa4i���~/<�#~�����D�?(�n��JE���b:��	
��,��B)�d�`�I/:e!��{Z�P���V�qF���0���_�",X�Z�x�������Iu�H&I�f�<��,���՘�*H���52q*�|:#5����Or�>�?=�4&��I���"��p��B�T�����Il�<�0a��Pi~��j׫T*΋���6��s����[ϻ�����,�I�V`��͘�A�'V��p^���N6mو'^xf��ڙ88<��݆�J�)�/�.K����)����˓'a���[@��>�\$n�'E�(�
�p<e�	��"k5�����lUV��c�>�* ���3GJL�������!^��2�У�/���^2���21R�B�RA�B�^�C=���F4�k�59�Dp�w/ç�9��q���F��\�F�XydUX��;>�݂^wj�0�����lA�׋�u*4.D�8��������$`��R�Ѷ`.���T�ڗ��7�ޏ���B7S�ː�������6�Pg� ���j���$1Лd��g�k>�tr�� ��}�����a2��/㦫.Fbb(���k��S�D<�lV)�5YLpչOE�E�?�/��:j�[��?"��7ήq�?�4� &Ry&7���P[mF��	d�!%��~�ǟ{O���^7�&#�k��ݠ��R��W^���aNC3l6'l�u"�ey�z�Yd
DsI<��3ؼk�DqʈQ��b�����e� � eRk�s���Ԋ���T�r!aɲ
�=�����c9vT����i��pˍ?E�(�2��L�#E D����&&��?���!�{���ꁾ�^����E,�5߿�|L��H)�*��pC��Ș:�H�j�!��K�����#O>��ׯW";2)�z�	�g���^��İw�Sy�j�e����^�"�KI*7�d��g^xѤ���Ē�B&��桩փ��:��㎇N��N��{���mb���x�w�1�X�dBI%/�p�b\��`а��N��(��ڃ�#�˱�Q�����_=���h��~�5rm����;7\{��Y7j�x/���,����SP	�����=2��r0"3T�sHr�͠B)���gΛ'�=�~&���D�q�j��gܮ:h�FI�כl�h��cR����ob���8�o���O��F��<�g�	��`,��f�l�U�Wc��-X�����"��a���ww���ƙ����>},4jJ�޾m��&�����K.���}> �#�QU�߿�l��~7�v���N+&��p�l����y�u 
J]�Q�DPc����@�lӋ�JGE���1��^t�nv��P�=�$�f��������s�<c&^{�-�jk����c/X�!L���G c����"�H+`%_@cS��)ޏ��<��kע��&�+�J�*���*6���+���(���TΤD��K�Z���}���H�%^_���<p�	[�p�aVRd���$=J��V��cU�V�D|�|���:��>r�ph\9�؜ꡬ�;e�:@U_c�I�������_;��� U��x]�ǅ����Y<^gj�fW�+�Z�f�J����?�- �@�R���zw���,n�w�2�z���`�d@c:�lC����FO_7�t�h�ݎ����Ko�����`ث�Y�C�s�
e�>��Ƌ��E���i�����7�r�O�ǈ��sr:/�&�)�V�x*)u �
��):�2%��:�Rx��,o|E���`�*x�O����<�: �Mh�^ڱH��J*� �"pe65M�N�%t�?��6��h���sp��'�vLo2�R&ݮT�P�L��D�B� �E�m�v��^���3109*��/�\�=f�A#=�^��h���X4o�O3�0T&`�?�_�v��9ŬP��kU������퀺�G��p: �I�N���0�&���v������B�D�lf��N~w��0�ߍ�xG.=!Pt�,
z�ͭ-H�0ڍx��o�����!؜u�ia�7��#�3Q���*f��Y
���\v�zC	(&�X�5���o�
[s#zF'�w;f3*��3����0�}��kd�<�t����=R.���!]����݉MnAM]#����=�6c������h��u
�VR���2n�.:f�2���ǰq�^��NL��&�p��hon�e����������]�&��p�K�e�!��Ťߏ�<��۾����bR��-�pD�\|�yغ�}�mmÒ��EKTH���ؑ�D�ߎ�W�\�Rx�>lض�:	J-1K�l����W?</?�.���C]M��o:nK���=*l^{�M�E,�G,��C�^E�_��u֙h�zQHE%��"nn2�[mnؼ5ML��Co��7ވcȪ4�f����i���ļ3:0�ьD8�ۅ��1,]�X�m�
MV�#.���J��5��j�&�8��U��w����Yc��ج�<FbJՓ0�4i ��w��B�� ��!��Ak�k/C�-�4�|[��f�	�����b�g�����[��Y�-�0f��>��P�@����f�>zV�h��j���0:��� 5:a~��X�&q�s��l�L�%�xh*�1���ŵB    IDAT�X@"Gogzz����o`�GbѢEصg'6oق��~\��Kq����߸�P]��h�7W�+�&���������5�A�ԑ5҈X�f�KTJ"�����8V�Ǔ1��i9�pM������Ƭ�mbPb�1L�_z�2̛׮�456�8�TR�T�h�H���2<�����"��
��$�{v-�>�FG�^�@��\|�ša���N�#+���A�T�%�D�p/�B�Ä����Ugg(��x�I�W�����?A�Z�H]��E�Ueq������lY���Su�S՘	�!--�p~�i��0��8�斜¦3g�EU0UՄMEN׃�ߴa�{M�fk�j��*�J�	�����4<�ֆ+�ڰ��G&���9aN��J�5q�j� �
#AG!ٚDCã��Q<����$j�O���(���>����T��BJ�	�SR3�(@���I�<O��3'��n�n�bZ�W>C*[#r���s��%�]�$S��s��0�ȸ�s� ���&�$�P�ζD4�ņx,"7����Gv�#18؏ޮ^y��;�҆�D�\���$�%S�c�K^X%�ł9�p�c�x�bšVJt@,�S�٠�K�6�x�i�y��h]؁�hX
����D��ϝ��>}�V��H-12�/�#���ՈTƏ��X��<��0�����"�ϦƯ���6+~q���7.@Sm�6���sS�`c�N��l��w�r�p65!^6���K����Z\��3��ip�7�Kg���KWb|t���"�;Lpz,���hlm�ko����>��,���hK�7�Ǘ]��x?.��R\�ݫp�	_�Z	�xN7��LZ��rl׾�"���.\͍��
Hr3M�P�Q1��/�֏���>,[�
ǜ�Y�ci�U:�]^8�6���d*i���=<��Yh���`��B;���[p�x��Gq����
����(hd�1x�ȥ#��xb݋x�oo��#�^EW̡��?��՘��C�<��Ym�ַ/��j�e�ʴ��E�\
�Y��7�����D.�֏��>�	��y����7�Сq�2�19�1�;��J�H��4�y�l��C�W;��#.]��+����l�FFP�+�Q�.�%�G�7i�e�kM-~z�o1� U� �CWLC_�㼳����=�|�P ��pf�̒��ŉB��迦N�w<� ���	Xm�T������՟�u߿N׵��"��n?:<���Z٨�A?��z�l����WJ_$G��+p�8f�J����b��b�"k�jaq��~�jȣ,���{��_�:��b��tOR�&&�rNک�dr`N[�Z���l�	,k_�\$�7��p���K4����$�ivX`�8�ƺ5kP_K)�򑩔�̤a3[E�Fph3ꑈ�亴ZM��蒦/�<f�	�\w%흁�	��M����{_ƺti�%���.��m;>�����	������,��@ .�N����X~D��^s"B&�n�y|Q#%��8���ۭr0d�A�#c�����{�m�.����.U�U!���Kg~�<�	>����\�y=�̈F#p2f'���$�]VT��p8m�=F�y�������P��0sY��5�TFi��"�I�^[
X�F��X@�h#K�u����
8a�wXMG����K�.`ɽ�����v?J��z���}Q��v:-��ǵXUB�
�(`ȬL���ǯ��(�__#V����UinQ>������)��'�Y��a-�t�l�c|p��Z�R�ח+��t��*�T��;��?��?x�o�/������.\��s1���*�U�d8�X$�ٍd��Q�����?4�Ɩ�
�!�����|/r�()H�.�j$�����M�9T�0��ݽ�H$���V�`0(7?�N�dq$;��`�/.*!�ӎl>#����O�FxΜ9S����R�mZ���b	k� �}�4@�$�i⁾~{����C�+��y+�5�V+YD���).��h�����񩼸�lz�Z�g}�+J��$��P^��`?<N���(�����SϮų��Cs�l&K$e�eą���9g��s�8��g#a����V0�
�p�-x��2o	���	+ŀB�Vmg�|�|�1\r���8�>{����D��(�f��/>��7����V�RPiM�$��ը5�1N+~��[���D�<>:.�d�L�3�V-���"�}�Elݽ�-s0�hs!���g��z7Z\N�p��p���g~�C2�����#p;t0�5��?��Kxs�F��10<$��&��P�^|����:\�����4����k��x�8)\ו��KO���o{58:G �
�g�·��5h%|�K_��7���~&&'`�١3�
�Q��A�.0�Ͽ��$��Y�����<Z�q��~��]��/�7��.�����త� _J�P`>\	:�
�?��ܴ��t^�V�I�~u��ؽe���p�e?��?��o#C�2Jd�p�k,F������-��l���mjP\����_c�ƭ��onê�G�o�7��|�j���$B�I�2P?k~}��>�
%d�	�A̮���9'�^m>�g�Z��p�� ���sa��eie��K�uo�����BAK�C���0N:��겫Ez%�#{���DB�a8R*0���Lz5B�(.��Ja��l���	<�<�����F&�DA��
-B&�5�ܸy1X�a��v��on�o����9�
�ux�A�(���2���k��$�b-�f4���T���/!<��^ǂm��t&#�>����p�?��v�T1xY�7�����ʶ�TV��3�-eʺ��-���v���Q!�O!N�Vh�����~�ضS�ot�nݹV2/ N�k�|Z��wj�e�B��0��߁�z�� �a�+�
̈�à�	��1*�Mr*��d��9LCp8���Y_���$6� K��Z����ϯ�gO>A2
���N��^b&���|&�b�����Y��v���<��x|ͣ���͐���SB*f6����@�s�Ai�HaTZY�MS�t���tM*�|�du��Q��C��S#z0�t�*�=E���c$$V �T\N�\���4��H%�0[�Wtld���	t���:�tnZ���#{�[�?�zӌԃ����ů���R'a�ܿ��z�M6���ȟ�MPf�'��4�g5�������sI�'0kŊJ��F��0�G�0濰�/o�rYɤ�e�a�y�1hk�`��&�sq8�q�Xm>ɐ��__�s�^E�P�<.d.���y�L�8�Qr�㤝|,���LD�����d�<c����ҷU�ϋ�_Ǔoz�*�E
�7���z��Û����<-j��(���*?/H.:n6A%��M��9D ǋ���� ���ʑ�MI�+O��IѼ0��#F�z	+fw"
a��8�_Q4on*dӌ���X�y����Ë��$�	��V�Y���1����6f57Ih.��L<�\>�ێ��Ay�V���+��8�^L3���Zg����a疭���bт�PU4ߠ���dP�9.,F��?��
�Ո8�[��8�ґ �Y<v�Æww�������\�l��tM�f�V"$������kh�ي��Ȱ^�j�����d�x� vlކ_�xN=�4��ydrqv�������Λ�ǟ|�vJ5;�CI`�QJ1�f�Zf������v�6�	���E�M�׬���<��lۻf��O�e��5hr�!42��＇��-M-⪊�S�k�ojDT�_𩧟��%C���a�鐉�q�܅0B��|?��'8�ӑ�d`����HdE:@�,X<���M��`���h  ���	ߙ���� <2���rn���X��|V�Y���:�^��#�
]uÏ�)����Qq?r��3�����_�n��z\�݋q�W���[2縘�U�H�������]�ݏd��`:%��j��b�	�:��|2^y��u����.��vZ1��M"X8��O���߇�+�¯s���a�dޑQ�l�¥����!�"f�F���jX��%{��Q�C8��}#���$�SSǃ���8.:�����d�*�DA�jZ�+nez�n��rN6���A��W�@"WCGZI����2��T9􊾈�}���V��Ӏ���I�~Q^X�*��it^�V�̛� �h�[��}��l�n�
Ah4��a�YجF�s�*�2aO�:�AR�<LV=�4�.�����1o�lт1#��`��P�n}CØ��*u]G�<7}���7cp`�H�lz�MF�<$��6�?�+ݖQ��V$)�mN�6�d ���{!�cX�Q���D6U��5#��{��;�[6z���y%/2�����g?{"ɵ�$�.K���^6z��d.�y�`�{��|V�+Z��<�<�������q�W;k�T�j�`�k��S��xT@83��J�a�23�j�� ׊�-|�s�k�˯�@6���]����:��x<>�
�a�Se�J�YM��+��V�d��;���YH&���Q������2�M
9Ac\�Ӣ<>�8FYU�?	*�j��f�2y��J�"YK:���ɟG[��2q5+ݾƠ�gVXG�� ���Ly}.�Sj��Ν+�;��d�E${Ƚ��C��d빗�a���U�~^o�����yQ����8� ��g7^�ʦm�k�fh�:��������c��a6�79���==x���%���T��./e~M�HY���(z�f����b��\Z��9a_�������{�DGטFho�8n��LI��4Gf�?�O���Q��+ P�����j	5`�XX��q��hl�������� ��������;���Y'D���<O^s2�:�S��rY�9�:j%���W���C �(岒�C������PW�� ��1B�����xv��8��_�I�>��3�(W�w+�9��bd<��[�b2��nF*����jw�nrJ<C��G2Ə.�n�fC]MS�d�����2Žoh��~��(��h-�4̟9��b�Cx�P*���I�<�k9��zK`��14��������R�F�7#hoiæ�>���7���ނcV��������,�(��a֜zlڴ���C��ȗU�&r0k��w7��P?6�}����J|�^GO�J���lm�o����w�b�!!ĸ��N�U������A��� ��{��]�F5�v�oߎ��v�1��!�!�
�f4bq�\lzo�^�~u㍸���-���c,4��UNI�[4��]���!$J��6��k
��Y��]=x�7q�/o��G#O�}�p_m\.'tf=L����(:�lAa���U��uc�k�7n�u?��~�k��d�H�<,�a|椓��3�!�N"U)�܀uG6�������<���fq�5Ի�vٱ`~;L+b����t��[0�OAc���S97M�ys���.�G67����8��2�6����Ō��}�=h�ӊ�C]��1�N�����0oN�_ ���O�!J�x�QP�j7"ap| 7����X�=,���Ũՠ�)A�*Bo`�@�B��-�[�r�#˝MFQ�s�������{����'��݀�9m�L���G��?܎b.��J�V#N�??�:uc�ҥ�#��9[�1�J�ܜ�v��a��1>6�?�u+l�B&�K@*Y�K���m��`N�<�̞�����Jd =��"!�UR���)Yj�L�".��l�{�@�.G��lv�]��X�xXʩ������ю|!#l���v��q�5?F<�V$d�4���(��H�"�����|�x&jS�E,�X,/��J=W2��J��A 3�j=n��T������o����% \ں�	�~1��lݰj���\�X@$5v�7�-;RBv9%�aomm��/\�(y!�}��.�l��X��`~b5ɞ`�nZ>�0���v;16:,��<�!)�f�x8pU@V.'���lU��i����
E���ى����I�j�������7>�Nd}�){8��{��o>~ou�柭����\�z�>7r��<�X��^���٥�L�Z�q ?�'ǰ�y�3�����܎�+T*{�߀��_��+��z_�?����n�{��a��Pof�[p�Q�1�΄94�� �#N��W���v�lq�M{3E�
+��q���?��E@a>�,~=O<YW��&s����bN.^j��pP��㘆��3Z�rr�V�I�?���X�)ȯ�{	�x���PU���Omt�J,���R���f	^����K���%�|fE������΋�s�l6-ϟ@�|V�0��j4a��+e,yʉ'�͞HF�� ��!nF�:��~���Id�X�j5���+�tu�ٵ���Y��7�х��#��\옯��Cv�������px�$�
c�
�
���Dch�و���T܆s�H�����*,�(��Gq�/~�x��3�6�"!9�w��D1U��G��O>���N��"����>�4h�%���%<����"],#�禤7uy�=Ø��W_���9�*H��/�Vϣ��Z�8^Z�>�@F�F�]���ᅮ�C��C�C���G0ļ%:�4�42���0�R#�8֮{�\Y#'��J)f���zD~�y�qY�b�*%���`@����N�ŭ����,���`C��h�Y/�`>F5��:�A\�58��FB����.��(�3���փ��	��CAk�h $m�LƊMn/6��6z�/�K,_��@D��\6��MqIP��ۆ�ع/Ѡ���	��*_���l~oz��E߽ '}�O�6��~�fŲq�b�\�
o����A8��Z�'$3Ԩ��u{���}p?n����������Z,;b��g����Dg��o������p9=S����X���蘷H����r�Q�>�;������-����<d�Eї�bqa=y�_�d~z��(��i�@�Q���F�F��\���q0w�&�ӎL�"�$�Xi8*e��U��2� ���F��(�܃px5n�Jyx6�{k1gf>ܺ�<�&v��Fm�l44�FO�/]��n�C���e�aq����??�Վ�y�i�
���%r
�Y����r�DpX.gq�����V�K�a��Eq޷�G���8��S��_�6 �z{E+���0aN�k�C8��#�ӟ�f-�j�ѧ�u�V��w����{�ףwl�!?���d6`��W�ܢ�(2����8���A8;�{oeW}�?[��̜q�I�CB	n��\n{oK�:Ŋ\��C�X�[�R�X x �>��9����gz��k��^�[�7keMf�}l����|>�0Л�q�����7�c┉���uڮڱx�b���Po?����x��ՌfL��_���3s�����+�����2���.Y^]V�M���EsK�<����x�u�Q��6	N�G,\$|��/�qR�H�{Y����b�1�MFZ��t_5�@����o��f���eO�s�N��ǧ��$F�\�{� v�/^�]{v��y[�^ޏ��c���^\,J�n���r�SE�&q0�RHq�kkk��J���K�f����~[�>ޟ�õxǎ�yS��$�C�;���!�n��5�\!2u��-Zz��(��m,4�x_S��r->������������������p�4��b���x�����=�Lhhl��U$:B��F�8���Mɪ��-Q������Dd���زi
*|d�i�l�
}̊��lr;8;��#O~���I�l��B�ڥ�Z�y��@ֳ�����I�����(��,?�&S�$��5"�&!~��&�1B?������b����&�\�jke񡲲��Q�M�І����δ��I�*���Đٍ�6cמpx��g���r�<��3���1����q������~&<kX    IDAT�ֆh(��U$:�L6��>��ݎ��脃[6�`�d���%G=�HR\�9�\�h.8�gV���.���SI<u���50ǹ��#�,�
�ET�BH�F�"�@Ux��G�m����5�MhFE�'��Gc&ʪ7�z?>۰����^�'1�l�]~Y�/�跘;k���XEqC�yA�WZKUTze�X}�CX��c���Cdp��jt�QSY	������v=�w��Y���p8u��0�:�5.��*�߹��+��\$=��j��t(���^�d�x4*�%�� ����
97��]����;�u��o:�rPԲ����Ћ���rLlm�s��IEN^P��EltԊ�)x��7�eo;�0�I�7�n*�n�X��t7�|5&O�(�ذ�
��)7��Í�h[����`�Qz�|��~|��'����5�U0JyL�҆t&!�C�=�QWTV�w(��b��>q�O%�(��a�����&qO�\x>��ݎ9�MŌ�1c�\ܳK�av^|�U��ׅ��I�$�����̨�g��ك�Y<�8��1yR
���Ō��_!Eh./�]����+�#�	���<b�|�rTޙe�޵�on(���F��oٱz�0��`O<�J�2$�ib�.�3 .=j1�9��.���])��:,�Q
B�
�'v���7>Bo�(�.'&���ѻ�@Uȗ�9lX���x�gQ]W�P�������(t
��(.`T�.A��)���{�-��L�;锉�x�~�L�.;f9�mX��0x��a)p��M-'y͉��+65Ǭ��n��ɢ�15.�*} 7@ȿ��Gq�wc�������mC��\��Xy�-����=>48("�,rT�OeP �M����<�t������F��ɢ-�^!}�t�S��\K�z�Ru��xqϽw`����G6����n���,��e̙=��mm-����S��&c��9h0h��B�{'7,�I�������g�Ը�ĤI��P{�r�'�/��{�T	l�V��g�ɚ�Ϸ��F&-Ql"��&�%�Z�d��B������G"��.�8���	��%)B�dR����.������;����5�/�,���e��|Q��}<NKK��~s���ӱn�:y�}�v��E0���.|^a�`�ou�y}F"����/x�裿q��e���u�ڣh����]���ଢ଼�`�Z����0}R-��w��܁�k?��]�RYE�DҶ{,�9' L�LKl������'��CF�ǟ��h�P�Dɱ�+y�g8\V�ǌa��;�� x��+�C��dU4���ʤ����?��a$U,��i��E�^fFr$]�i[���'�e�J�OW{qR�"'*��x��D"��&��[��~��	 "m�ښ��+����?��q��xoo��0��/���6`����·��>���xw����Ftt@�y�O�d�\���̗K
���8�;�=��Og���_��#bv�ً��:!�{�c0����Ͼ/�"��KUH�, �$sD�������E�]�L�&L@dpf.�͎ƿ���ftv�ǣB1K�0�NAuM�������;�ɗ����!DQ���ۦ�:���@�����0�!y���y!���TL�6���0n��!,;�L|��z��)�A91TS���=�D|�b�I�E�B��.O}�D��K���_´��KG�S��K���A7Jx�g14<  ��YH&ݪղ�H�ϗT�����䳯���SաX��:�c��}w߁�͵ҹ��b�`L:oU��p�����=<��xɬ!9��ء"�QM�����kĥ� �EM[���½�3���8����ǟ�@���
I�U��/ס�2�X���9�u�l�
�T��W�s(@mU5�����;k��g^ �k^�������j���1���_tF����"�hǮ�hm��G�x[w��dX�C�S�5
BR�04z��YXv��8��S'���N��j��Mؾ}+��/J��h�5u����T�PQ��B�3�#��O~|*n�}.$�ò��J�iSh�����]v�(�u�}Q�����$�P"�hG@o��0�6Ӧ7��VǢSi�"�uU�b*K�C����G��Q<��;���vJw����
�it�ŗ���IF���I�0�Ja4n';::*<4n�15���ظ��K��o'&���T�|�	W]w���,9�\JԻ��o^������zDFiy��郓ٞ�8V3���{�U��TA�ɧǳϽ�eǜ,ƩY��ށ^Q����d.��"[�I,0a��ܶS (�U)JTU������#Q��&/`��1�) XQ���^x�M&���lj�
?n��F<���ؿw'
��p��ǈ�pL1��_�bp�鍆��&,X8�*�|�歗��i�Ir�-6��m%�Bǡ��m[���$�H�Z['����h�"�#�A�,h,��s_���n��(P��6����_���-������ $��Tv��l���>���}��������'������x|ޞ�4��4Y������3��`v��E���c.�O@ȿUW��c��v����3���뺭���������ו�u�0�3����~������CWx�����(J�(lF
�5�2��ܚF�������*%ì9e�D3;�����m\�c�/%<�d�F-�T�QHZ��qޟ�4���]2�vX'>Or~�ϋ� �'���搜<�5㸋ρ�|�,�nq�H�'@c5ȅz�HU�R����`-9��B�8� �nP���(v�m[B_�;S*!��!�������z<�Z�5�!�n�i���	��E�&�ŗ�����;�P�gC�h����D.Cm�?:�?p�i�"��� pdtP��i�DFF����JrU���è��G,���[��YSq٥��?3Q��I�ɑ�'`ڑ3t�������Jd�,M���	���ʸ��[�ӽ�K���3BO/�|�j�1D�d\u�]���](kc!�n�*��]6TW����c�*�.�\�@T��Ʉ�[�4L�0O<�����xlݱ_:TvME*CUȃ�� �����P�\n�wY$��c�{�=��/��~��7$9v<7�B(�Pp�eW����� ≨˩+p�u����ˤPQӄ�oz ���=�2�"�72E*k-řC5���[1��	H�Gd�gg��ɂr�t<)�H�g/�}�<���yP�ء�3QQLg����p��x��;���~����b��1�zQRt؜>\u�����m>&Vg���*J7��ꒋp��+��v�ri�)y\x<��Q����g_��w���/ƣ\|9r���W��G��X���z|�?����u[�@>��3d�E�:��������PbD�^�P ���!��V˖.��S&���Wa�V�?}����D�c쎻��\���~��R�#
�g���gM��ç	Xa�7��]H�h�R���V�t�i�Ӝ9�F�)���b"�r�M�4�u�a��T@42�)S����9�u
�Ml�Po���9,T+*k���k����a���4q&�{z�j�J�{�u0��	8F"���?���;v�����*����~lڴ	;�n�xI��`��**q�.���3���P�Ev5ݎ��۱��O�s�>�55b�)�Bg{;�o�*�}��ðkw;
9N�_h^��#���[n�*�aL}=���~��'R\���0i���v�o�݇:�����\L����U�J0�kks3Z뚱u�F��1[.�6x�u����	�gh�-�-���Uu�&z�U8�?���(f1-�ų�:[���ӡb˦��y�t`��_fc��H?�Λ���/�;d��DK����i��Y)�yN��	�&	p�g�Ԗ-����$`�#v�>��#�<q��r����HG���S~~���p��G�9/QUc �]%>=:y<���ʸ����.�p�锌����2���CEH"�>��S������򨫫�\�`0  3�#�ځ��
D"Ql۶�-��������JA��? 1O|<>>;��,�ڵk�X�(���W�3��e455�kkk�L���Z���op��ws�7hO�D}- ��o��������S-��.�T�
	(�t��ˤp,�C��ы�2��d_E�&X��$�:o#9s֤��S�zA?�r�0���+6���嵪U�9��L�"����H��\��<9(ʈ��R����-�K��g���vZa�B~�
bfg�h� ��H��TK�Z���ɫ�2���FQf_��6��3�ј��E6Ckc-N<a%�?����k���#���CR�~�n^�C���
���!�`>_\�'�<.�<�8���sP�&�S�v�%�-�L"ˣPV�a�|��FĲ)�[H���
�����U4T���e��5�~�+��c��)�����i�T�M��\���(�e8i����VT�<6�|%<���صkFG���\?����|F���V\{��X�nl� �c�NC��i��N\u�o�(�Ԝ�'��^i���^=�����#���?<���h,�MCeE #�0cj+���_}�>aT�qDJ��u5���)�����껟�#[�����0a3��u���s�D��I��v:d�y܈�
���A��Å��	o��9B�&$�9Qr��9hnJ�K���P�߿�V.��h�_�	�
u��G*���D]�d�q�q�CϢ�3̀y��d5lz��m��[/Fm�[�I��g�P��/pz}�%QUӈ�o^���Z���792��qI/�)g)9����~�7��ӎ|.�l:���&�X��S��D˔�p�#O���;P)cR.^(�`Ҩz0���,?������� ���u$Ǭ�����Op���ɕ������.�Hb�F6�9s��1�X<g}�tTU��o���K<i��G�ƾ�n�h~[Rd�Y��f����i����QF}}�:-mT�ص=r���ذq+b�R�ܕH�
±A��u�ǳ���J��4�h� l������F#��(��^�nw�����˯�E��%����={��o�^|�tZc���%������%���ҥ�K����k�N�Z�@�8V�z��]E&���W_�o�B<��{�<'���/�e�v�N���c��;w������"�z��(.���=�WG.����V����p�H9���i���/����������2y
��4�`.$#CPL�q��eW�����F)v��R��̫�.h�0�Eo�����-@�G/[��+V��{���U{!������
���&NlB�kǞ=[఑��GttX����v;m%��K"��iq�QK�x=�4�cǉȬYs�3˝��z��	Y8qo��Iгc�N���;hii��=�tr��8�9�ɱ�r�z,Z�@"ո߱1��/��vÖ/_�3fH׋{����y�qu%� �>��TaRL@���whh��T'Z�9�����bpp�x^�_�G5$}��HZ;��h�D2�0����0;;��x"j�!%�K�#���u�eS1��*
�t�lh�S+*��L&�_����G���4A@�T2r~�/Q.���n��97�Nj�r�+z�$�����s���L���'�^����z����NF�(dH'F���$	�D�3�4���Bd���C[ ]%�
��u9�	̨�cw� Hl�2ǝ�I�&�fw"���m!�-k�)Jr9.d��Do>�b2٬��ɇ!��z ��GD΋��F<n�<.����uL&��Z�|���}B>��+����D!1̴T���;�vڤ������
g~�T�\q$j�H�.@Q���C�x]6U����x��ϡ�*��8��He�U��/DP�G��b�"\���������{��p
�x�=Cx����D�;)_6U`t8&uuȃ��J������kuE�{.RU��b09��?�C����t^3�JI��Ԅ<��ظ�3BC�eC2��U�����	_��޲|��`y�/�"|�g�8�S
����0{F3"#�P��H�9������:a
��J�y�p����m�Rt������\�lS'6!����>�$yj��re����<M��H����E�^��� _�չk.©�Q_冊�|�AD#��s;�0�$p�4!�t��\ϻ�:��ʇ�6K�X�y6E%�b)���W_~>V-���C�h�8I��|�QQIBM5���'^��?S��`r�ʹ��s���p����)�L2"�$ռT���e��|ϖ	�q���Wއ�F��������6 %��#8�g���g��Tb�İt�hkۑ��T5�a����?
��>o�5���D,R�ťy�7�A,2����+^(����[�[����ٜx������J-X���A	} ����@C}%�OoÊ��Ċ�G��uY�~_�X�|��z�}�Y�4�W�;=_.�d��-��o�v�~K� �t*.�������o��B,[DCkj��nh�ҡ�a(�ٔ�ёt8P���̡��3\q�q�K��#H \Ƞ��+Y�_r=���CE�LD@$��w��.���ą��pdT���(m�Fsk��;����aw~߾=�	��[oJ���h:)��������Δ�l���hnj���(��&L��pm�tGv�ށl����2)��\�����gT�y,)�<f���b8m䉔�;�{�>��S�|�X���1��8�[����bۗ�"�T�s�(�����yT���B,�|>��*�v��5��TL��#Y�q�X�ѧ��0o���%K������3��HZ�cT�g�Q�e�T�1���wo/7��Kp$�Z4G�mV��p��������9�!�\���wϿ9s��y�$	vq�dO���V-!?��{I�������^�r����q�����ۑ0�����0-����fQd���H$�ɓ'k��Æ7�Wb�X���ʦi��D�MMM�h4Z��r%�ۭ*�RTUU�u��H$�pX�f�Y�4�Ua����`.�/�t��4��m�af.�͖����j9���,��u0ҩ�����<dtt�����7::Xy�@�}Ѣ�[2��$c�1W��?\,�d2Y��\��R(x��i�כ�B_!�}- �@Ҭ~���yg���*�5n<�Rƚ��/GDޜ�ЪA�<��V���k�ѣe�H�&κ
�8�Ovn�(�|`穐�Ř1lIs��9r_�!!B�1^&)'��/�F�e�$�c0�(�If}]t��#R�D���:>Z���D#XcI	
�A 3�G�c�:��#\6Z��'�ɨ'�Ҹ���F.mH�!G#E�.
���n��Chk��Yg��U�.C�9�Ŭ����J%�%O���=��l��m���*F��t�2m��d��sq�Q�����p��0���{�����=�D����v�Ͼ>�@�@��Kx��VB�߆������k�ń�h�L
~��.g#����s�*�7,(����؋e�Fm-�rӥر�+Tׄ�g����mR�2�rh$o����N|��6ؼ(k�d�94�1����A*��+���9�M�붉�$�zev���5B޽���p�}O�l�G�Z��@�����YL���$�r{��(�����ɔ�����/������{�A+P�4T9%���G��X���ԲMƻ�5���(ӚE�₋o�k6��o]F����R9��K��W_�E��Q*�Q��,���0>/�ܞ ��&��G��C�����A��E�O^9k6������ua�>�:��>���qt2��t����}�Sx=�P����L&Kq�<�b����|�18�;*+����ҹ�0����f���s���݁�|��]���#>��Fo�>�Z��fNF��ķ�y�v��r�µ���ض}y�(���*�ny�1E�a�^�&f��������sx�Zf׀��M[�a��=����A%5����MU�Ź�C[k�>������q�o;w�ǚ?E��    IDAT,N[
�8���>�2i�Ixym]���Y�smb��U'R�}t#~������FU���a(΢���^��j�l�h$��8��t�/�9���/�HLx3�MM��bRXrM�C����O��&�P��*�k�A_-*t=.�$؅c��r�gb�S��ۃO?�S�M���a`8�D&��_�+���P���$N\� �\}\vS��јxD�Ƅ`����|��n?��ga����E�`32�Ӡ�<�|)k��1��E��A�ِ7l(��X~�Y�H�'��_������\�L&���a�y���a��?�(+�ǆ�{�c�1��itw��n��g���f��]\�y]+�t���p�G����O��ְc�������"��@�V+UV3bL���r�"�<zM�yW��͢C���� �E�c��M�ʆa�%�(�����*��g�BQ��R~����JA����Z�1�F��(
-���%�T2<���̛�=_��U�}�uEOB3����%��J�0��4VL�PU{QSբnc���mf�^6-e��WL~�M�PP����`M��V*��r<ޞ��(��.�|�_���_��ka�	{�nz����j�;_���譜±d"*&!�[]#ߩV�D���@:ˇ�z���%h`C�]C��<Q9��ŝIYA��P@<��}U�'v���D�_�:o���;�A	x�LH��g:��>.�c�������c�Y,�3=�]�e|V�A��Pȿ"#������nb�iQ��̱T0uR��˅$��+�j�2�:�(�U��q���1
	�#�i���:|�v�NY�\Q�v�	�RI�������ۧ�$>Z6��訌�	�H�K���x��O0���~i�'H�2�\r�k����.O�׍\1�x"&��b	Fr8�7�a4m"^`ڪC�i��U5�\tb�c�ރ��["leE>��"z*@<MRmο�|�� tw�ÉB��n�*-c\�U^w�yX4
�A��n�#MJ\	˂��V�����?��������"W7�"����b�<p�R
F1%]rRt�K����ћ΅�/�=���s?�e'u�p�:J�^v[���V��P�eS�7�^CQ�v'L͋�/�|�W��X �$H���d᳗p���ܩ����B"��
Z�������~��q<��05?
�&�0�Ut̀�V�S��ޛ�Du��h��� �ހ�02������n��܏7��^w3(;�����x��$.<��8���ؿo��K�T�ÔIm2���S�6g1�}�i���s�W6�f�D�\.�㐅S/���S�u�X<�8���������aɓ|����뾇Q(jp�}·*�-�%�&��9TV�1��FF�G.<\̄Iy`��ˡ�(�[�9�zg-�y�(� a܄�~�l%�蜳���C�G���FF����GgWv�:�������<�'NF�P��O�@=b�,t͉B��b�`؃�N9�`�9{%�|f1���^Yi�&�PU[�X��Cz	��;�Rэ��A��e��ڋ�+H$b�C^��-͍�Ƶ�J�-�7�c�8Atww
�%'�~���#7�� ��
l�k�r���g������$0�d��eho��h�1<��_�/8����CEG.��V_/��0QD��Gk�V%�V��֝�q�X�b)���L�Bji��B��B��E���5�p�㨗�i�AŁ��H���O��_}]ޏ��fx=�ń���;�-�B٢�p�\*�0o���<�vA1���Ɖ�����eV���)�7�I6�*<`��8�$��_�fΖ����L�O<���,�ea��]��y�h�"K��r�6�-OP�ry
�|6�t�3��V�PE�r�����ϚnK����T5e�J6��GŐcб�0Ԃ�*y�4�s�i
02Mݰ��&?�M�a�s&r�a:���?���w
r3�L`��p�	c�DM���Ѕ���c l�/��+w������δYw�������3�z�+Wb=�Y	�
�:c�O/	�Y���e&������B�9�xXƑe+���0qV�G!�-�.��q"��r�/������4�ᖉ\�H��1>�؉ �
���(��q�0|x
]�-�gM�jX1q���8p�O�����\~\H�70"��]
MEcm>��|!�ǮX��[�	-5�8S4920wp(�w��_m؃	�恌$7.���P;3	�H�����NƒE��p�Q&��fáC������>�o��!b�,���[���KS1��]�c��:�p����9�>�Ъ�yv������hF�S��(jZ�b4�A]�N|�vm؀�
^�<�������T'��5���2yC�	��y������\!�.r�hzʈ&�a�r����h����=����B����EM}3�u������O�[�C�@Gt��CM��H��շ@-&�q�ɎA���+JwM�ŗ_��>�
��R@X�h���t��J�	]�`��W#�²Cw������fjxTG ����]�w�8�K��͜�L�V���S��0�M:	jU,�o���CC�tQZ��6��>aGɤ;����B.����� �+� -׫�ؑ�������pm��Q���zx\M0L�</�0���b���p�I����]���0��%;��tN��.�CO��_]x5&M��R��M0����.�i�Z���7O�i��$�>�5U�c���������K�ή��+���2�f�՗�n_M؏�Jt-�y�O��'�ļ�3Q*$J��H�(���y�<�����,���dE���!�F?��w��B��߉��C����Aߡat��c��}(6(v7`s�����v&�%����p�\B�/�I��Q�Ob��ñj�B�v��s���i�)]���W�����k�œ�}��~���.|�@W�A��Lhi����7����/_&�tTg!��G�nG%�huvd2R�p�Uòב-��;��|Ua��[�f.^���aE�h��ǣϾ�B�	SuJ��GNǽw^	p�-�124*kU��t�h�X�����c��1ˎ@ׁ]Hu���Yi�JI1"�	,G�.���vYGseeŇHZ��9�PҼx��ȣO�������$>��
K�����[�h��"�w�4R�Y�"LC�LJ�_\��cjI~��� ���T��5��p
B�`]Z��geMX,1���/�	�8���r�'cΜ9�M�t*�����a�9�
�A���G]]�:PPl
;YE��.E)8{As��RI+�l�B�\.�K�r���T,��b���rƤI�ƻR����?}]��a�Yw�#�m���3��O��K��Ŕ���ǎ��aTB�[����b���I�s�Y`H~����i)'�G~����JBL�J&����r|��xҳǛ�.�`���g]v�Q��Jg<�^Ԙ�#Ǳ
��7�7�O��:�^Ƭ3xZXTWV���˶rV����R���/��GUP4����a��>�\*�[uV}c	�Mj�P[KY��A:[����e�>�����0��vg�"��)�?]͡���'�ę�����j���J^��+"�+��w�Gu]�(#����bUQY�d�X���>�`�����#f��~�����N��F�\)/\'*$���d𛋮�ֽ��h����	6?�U�˳ϣ�k��}x��;a1�c�2VD�=�� ��&��<� tWT�eŐ�K�3'��k���[���"�u"9��L.��P�fܽ�Q<�����M�d� Õ3��thy��M�D%���t8]�l4{d��]v-��|to5�`�PK�^΢��x�(��r�҃rmx^h�W��v�jY�0���UW߃?���Y�|�_��F���Q_{�o0eb��^c��K��p �T�M�C�<�'�{�P6�����G>p���MD*�b@��΍��(�{_��ݫǇk�I'����|d+'\j����q�������ס�7&v8�~��7���C���K���N8�H��3D�m�
�Zj���O��˖���/��s��i��m�־�O�cO'��2
y[@
v<.;&Om��Y@"ч�G��駬�&�U*DAͬ�X<��>�~�-h�
dr&Je�m+r[R-n?������MI#t�����ή^���uB�>��`*�5�cY���r:P][�B���
�vv� �®�0N=���8q���14ԇP8�}�{p��wc(�G4^�� 4�#�����_{)jB>ḱ �� ;Z[�$��I[�nB>K~�L����j���ۅknjFS�D�]^d3i1[�p�V32�(����o�]�،�ڏ>�'�|J�C ��n<��N��Cws�5�8f�a��K��a��X���/�q��ã�ױ'�|�[y܃�����ОB�H�Xbj�+�eƪk�%ՋXXp�I�!<�ԋx��'E�O��6a
z������R�j��Hs;�V�� #�D�S�\�XtD
�Q�Y�]�xk�|��T�3� QDf*��&\�qK�QlFXn��s�����<?�DD氻��}��r�3m��M�,�����ɍ�n�;Kb<�u�&~]��_�q��n�5w���l�\�V���%�p�8:��XUD^Lf���̢��Z�Ʊ*�Yv�mK�';Oc�VW���c E��-v.y;���ǅ�T�\����=ݯi�I��⍲����aK�<5$A�cU�8��EF�e��q'��1��c+���W������x�����A�in�8�QŤ�H���"`���-��s&cBs<^�gt��͒��2�>�d^~�m��@��ɝ	U��*t@A"ҋ���X�t�lp��-0�9�����/����:�X��:��iT�6�0�py�hm� �*C��1�	7_�;�۽��j`��\�EU�~oX��������!��(�;{�{zPHK'��k�d��Z@tx@ԡ-Mhkm���0��
�a\|�mX��p�`�N贩ȥEݥ��F	�_C��jD�:P�u�̙Ȍ�ȱ5���hl���>�Ǟ�T'm=��!��D�T����o�Ѿ�Ќ�N�d�9]n��*��C��'��/��}���F@�)o3sp����ߋ���6ՉB�
��k!p��5�}a\}����m�y�!'���Y�CS����o��,�߆��=�Cޡ�c�LPz1(��£O��Ǟ�+t{e�Dz���
͏�pky�s˕�:�n�I*�,e҅t�o�
w��>�t��6a�'�⤂X�C��G?�6�;v	:�H1�봐ˢ:@}?C����kq��Jװ�_�yKFA��*7�j��6�Ǯ8�.��,��opH�;�~Q���-�ߏR���nT�a�v$�I���3�(U�࿾{:�yƉ�Sg�s�����N������xoͧ�fLdr*L�%ݷ�?�Dt����a��46��ȹP��J��O>�ƍ��+شm't��K��&L��\��P]S�M׋������.$��T�bG.��bz���~TV���} U��8��ΔѾ�_-j\ ��im��ߞ+ L����	��0�?Xuuu�1��S��444 �N��pm�&��d�c�Aʚe����q��CY�:���!Q2ǝp�+�oف�;��W����L���M�b��0��z��(f��,���洉�P*����-��@��c��
2 � ,Vf"�N�'��ֿ2�0v�b9,=��6<���x�ٗ��V���k�~	������xE+�XH�a3q�K1p�]��qm�ZN�����w�{�",�jRM8�8�������{���4����^څ/6.([�t���p8\p:�� Y�`���ոP�J@��|.�� ��E@���_�o�֞ohU���i��'�2�C�D� ��rA��խ�C�B�,�pa%�[��\Y1(��n����0Q1>:�w�^T��6cdzM4�*�M�@�M����B��?Dz,�{�v��-&<����8��8,�Y������a�c˟�1����A�u*j�v�l�yk^�Oi$��$��A3�ƚ0�R�L����יWz�����[�x#���bi!A[�^�+b�f�\���8:��1y�$T��0��۵���Oqұ��s��q�����{k�b�ރ������1� �Yuu��pV�X���)&��q�e�@��=�2i�,�%#M7�"g���@,Qy:Sp�:=��D��ŅgS[e�-7]��h��0z'1��d��sE����!\v��b�A�^�f��$�i6�p:\s�yhm�@t��0�
ټ��T��.Z&MÝ���Ͼ�Y/ �b	B�T�5�u��0��s	�q\@�벢Z��
��������}�y�/{D��8��jAw�u%��y����e���B��aE��_����t�����O�03��E)=�뮹+W�Fw�^T�*Ċ�Tf��Dv�n_5^~�<��K���	z���S3������Au��b~�.�P8_%�����`wye��g{�q5K��\Σh�P��eBG����pܪ�<�p�F�y��}�<��E��mg;������߀l��&���F�e�M>^c}������Ӱp��{N�i6#G�,��1t���?<�X� U��D����㵣�~_G?��٘2�	5�bq��і�\�����i��'_l����O�s��K�j�>̚ނ���ƌ�M8�9�����-��e�6Iغs�9O�������@%�=7�C�@�vMF���@�^����S�{���W?�i����!x~�:�t����x�K�����O��K��	*��ae���!�̄�&��n޸Ih�ѥ�R<I?8��`V���ǬJ�Dj�$���p^Q��bVXP2�$�C4k
�.]�������x��q�'��RSڂx⑻t�������!lٶ	��0��µ�A�	��l"��ν��w �ČAXZ�(�a�RV�H�7U�
L����8���^x�M���[8x�3g��a3��Ϳ�A���$c|�Yr�8�4=�q��������� ؍��k��xt,��b M
�*��L !��"��Й�e��u��tr�1�jxSL�-�q�q�q�9n�DW{�#���
���W����(��n����ށ��i@���������5V%M̂\l��q���$uAFO�1��9yB�mƫ�Չ���5�	a���;���p�0������t�YYeBp���	�m��VO�E�xS�]��D�_}1΋�<��.��E��?���?e�6��=~{� xlza�Tyrl����U��eG6���JW^q!j�}Е�Xl�j��&�H��ӎH"���a��ϯI�˔�#�7�m�n���ztx�z;���o��~����"�R�t^x6mE<�,8?b�^{�o���_�'�l��7���ϱc˗h߿7��;�غ�[d�P,g�i*�B2�*Q*���_]��H�p�lJ<;��됏Fa����uKEJ�?;��/��b��7�#�K���1��5�K*[�v`�2���_���'c�i���,�$�@�c�������S~vW�&�y��)��QP���~�B���٤�֜n�����`-���N|�� ��F�K�׎ff�#�#�p��[n����t�UΗ��z/M�	�T5������'۠{�)h�X6E�_��2�Vą��K�������":2�l1U+Kު�@E����1V��9������Q>����2����r4pT��da����gw��-�`w��}��.��:��M�<�htT��N=���8����D���,�n%g�h�	�d>�2�棍x��7��� K��2�R1�\:���C ��c���8l��hO��rI�։TC�#ؽ� �~�e���x�����k$E<1 ���������`ڤ�"�Pʚx!�
��8�3�M;�㍷?B�t�H�+"m��    IDAT;�\5�Y�=:��h�q$�OmƼ���
ɚ�Mk�3i��r#����S9��J�ME����ʆ�NE��F�L�14B���ӏ?�2b��/����:y#�{���]�;�+�X��_7|n'V.[�K�CxșEI8\�]��;lmh��9K�|N2
�Ο/B�����ip26O�|Z|���e����n,ޅ����D������$F�س�}�x����k��'t	�*���{��P�2�ߡb4:"�8���ϔ��b�W�&~��g@+��Fl��e�ͼ��3�f�V�i��"2BGQ�4��c�QǊ%�o��/����aL�83g�����!$�d
eI8��{��iÃ܅���"6o���P�EY���rgQA�[v��Y
y�ұ��1��q�>C��  o#�o�W�~g'��8�"8�d�r�J1U�E�ǽ3_0n���o����r��_�	�����i�� |�ӯݼ�=vB�^N���K@�,�7�Q�s,iR.^��i�i�h�L�Hv���1�3#W�#E0ˉ�9JGl�I�:�-��PH�Ęy�Igv����bQ�,9���(--�;��rۡ�Q��������;(|\�;k1��@i��c`R��T��t�+ ���?:f�RK��9U���WG<j�
�*I�
�eM"����O�᳧K��v�H਑�0n��T�l/��:6mމPE�ڰc�NL�2I�����l�\���E1�����Q���ۅl��_{�;:A��(`ǂ�me,^8]��p�5#:҇��)��2؍ �-�Ӷ�S	��9�^��;PP�x=>$"Q���]���p�u�Jn$��DZ ��n��R��r��V�w�߀�P���BHwjv��s%N��o��v2�m{b��۶ms�	'�&���Ķ���^��߰U�oO�S}�������J��/E���܌�����Pt{X��
�WdЮ��9�f�p�rx�Wm�Zb�Y�-��D�$��d�����)��	o��u����>N����LA�o]��]M�\��2�����xA��{i1o��ny��B��a��kB��q�D~��Hh�K�]<L-���,4EW�1C��B&Q^~
�8KQ�P&@�ڏ�	��<l��W��.��Ûo�-�Ʒyb�w��O{�lҌj��pҕ���^�1	I���8cC�U���^Ɋ�)����vtߏ���T��V^p^��C�_$��j�]�J|�C/��qv{���˥)����h���+�m����w2W��S�$А/�9T��ی���B�R"�ӱ�ϥؿ���S�;���3��cۏ��;G�J��y�e��w	��p����	������u��Gp���[{�ĝ�g�ܵ�
�L�N� 8��g3���F3\v/�I�9W��t���_Uer�,�7&Cf�Q�SPqn̦������k�>�{gEcq���QE^��~��T5v��g�Cr���+�����;>KY�~��fԒ�%�6mZ�;������Q�=FaN�-OT�n�Zȗ'E�[h�}B�붴����þ����u�곲 L%(�g�8s�#s9ҥ���;�ެ>F�8'�k����fh������2���E�.Eƨ�q7ҥ���(P�s���䍫&�_�R��sWr�l�?Qv]����8grZ��zޣJ����5�,!�O����-��t=�t���\\���$Ǔ�3�TQٺL�[�p#��>Y\��	n�
8G�/��������8�m�7�c���SV/A�{2�6?r	��H�kM��`y:��%���~���+��������F����q�zk���{��֏F�V�3-�}_�x���j8	x���S�U�L�p�[�����>i�3���1������d&vCAH��g�.���K��$ȕ��Ӂ�5&����4v8��B#�oE��8�Cy�+`�4QW��.н�+�D����j1��a�ipW�C7�'"c��B��D$dE3�H���f�7 s��M@"M����en�~��z���p��[�jYc���I��yY��y���x�s��4���+�O�OYL��˶z�󤦦n/ߘX=���f���Y�F�iںhӜ�U�z��
 �Dm����W.�Z�i�x�x�v��{�L+gp/-�n&������M�f��:�(�>\;���J�ݫ86���vt_�H?����6�������C�'�aZ�XH����Ҍ�|��t�t��MRUQ19��8��ӟN���p�f��&��Zɹ�UM98\R��s+�[Ѫp����׀� �U�1��I�޴��O�<!�xp�e[S�G���$&�aR���������R?�NV�` �"N����k����M�ݠ�s� �`��bf�NS�/� rg�:{埛�KYF(HNk�G�Ǉ�s����z+���[��̻����F��	I���~�!��*��_�	3��Q�%�g ���Dꉹ�x{�+�9�y����l8R����C��o��x�cSA�q9y9����m�4��/�ɔ���=�����$~����LK�w������ �����Vi��9�UcT'��N��s��c��G���G�/e\�o�_����Kɢۡ�i��]?߿��m�Z�w��h�82gh������z�:�g�� ͸��˔��-�ı��Q�lO��7�qNQg�W��Re9��:�g��������*6�~��<»�&�ɜx\����XV�s|�Wʞ*�L�"���$`���pz
���*��/f��ܭ��#WT��ϝ��&���3m��ǝ-9�Q:H�B��R�?wآ�U�fTm^o;�1��o��B�N�v<5T�Չ(�t���{!�s9213�ճw���I��E[���9-���>�x�=�w����y'y�����~@!Qp�6W����Xސ�z~Q�YL$�xx�C�W;jU"}߁[}<����;��ؤZ,	g����w�Ν�ζ�IJ��	i[��O�Ҷ�t�z;��o��Y��)�"��ރ�~[�_��>�w
�e��8H׸'��(����L��?�I�.WK��)LF�"b�����2��U+��:E �^B���#�Ea�ߧX�e�N�z���q\<D�>	=�s�rgZ��ڨ,�~�H�n�~<�|2}|���-3��GR�P6-w"��"�R	"7t~�$z�ܿ��XQ:(�����7�_����2�J(B���u����]8/[8�����`�����^y��QL�}�\��s�����q��όަd��ND���*[��S�p�2�?+QOt�_pYp
��m'���n?��6$\F��Om4�*|��p���=(�#�mZ�ƽlZʸ�����d�wO�"K��<�N�f\�΅#�W�@#r�Z��M�̦��5�?;(��m�^١����6����-��_p��n�Hʸ��E��S���^�XI&ǋ1b����N_�+5�,� ȘH��������s�c�'B��c�|L�s�$�?8�v�K/�9'�?����&e&�!���t�Vy���(Ιq�}�Z��-J6*�g�ig����j��Ԓ����|:�l�\��v�i�û��5����\��4�3�j~(J�Q:|�;X7m-qtن:��"�>R_\�Ϗ|�5^+��(JHVeC�׀eӟ|��̊�Ș��z�v�����k������x��L	�<�v<m�Y;x��4)PY�A��rJKI��]���XW���D�`>��L�'S�Cl������������*�fph�0S��oJ{{�M΂��x��I�T8��E{<v'p�yi����r�0�A��'D�c{��>�Ǘ��})��ÀrI��)�@m���/ci��I	����!���ysF<�X�x��į�M��3� ��
u�g�A3�}�W�J�vO���9�b8�س�BN��x�c�����<����mJ<�ZiŌo?T)��;:W�'c��ǆ"o$��sM��#u��B#=}��XS��ܩ��K�}��l�lh�_�Et��+��%���+���* ��.Z�0#]��	6gus�<�w��{�)��E�麗eN�Z�˩����� ��G�.��1E��:>�Ip�z2OÅQ�F~aWP"��p��O�_4J�)��[-��N��}�����}������/7_�U�L�md��ty~ ��i�侊���"�&�"��Y`�_�9��A��l�*�\��.���?���sN��p��y�v1��J :p�?�V�ڋ��<���,��=Z�q���b͙����w���V�w����5��r5[!�B���4j��s���s��W�ǧrR_
�o1�ȩ{�3��]8
�ވ19�W��@V}��-R\:W�"���}��1o ���zο�xo��7��p�ꫢa��z��^}]�f����|z��v5��� H�y�a��y3!,Ϛ���vag�A�I���������qU�U����F��D��'��3�e�h��`��mҾ넂CY�\�X�?^�&�[�x~��v<��}}��V�z��	��3l��M�6'�*��5X�O���i�����L�'mF܃�2q�b����<�O���j�Q�x\ƛ#^�{��gnAv"_X����گ�Q������*p��oȴ*[����xGa�1ӡB�'�®t/���2�;.	_%��SD!��(t�p�azlZ)<�ڈxY��fev�{	��궉ٳ�B��a��~��DaU��`�~����]����� Z>�w��t�CG��,����A1���fħ�hARp4��H�R��hcY	�۷i6��W�<ϐ��08}:��@�\�u�8B�|+����0���|U;�׼M�x%��� �`#�w���ч�$ەu�(��������8n~�ptyE���̒v�#V	=�)�B�Ŀ��@�o�!!�55����X4
��8�*��ۢ7o�S�tsB�a�Z���] zt�Jb������8��մ�F�4��,Y����E!t�k���������+���1��p��-����\����`��x�[ԫ������%>>el�XEl�gQ��� �JB�|OD�i��P���䕉��C��#?�E�󬗗	�E\b� p	l��i��o-�Tٖ��M�1	&F@D�w�IAؚ��k�}N��F<&�iz{��>�A��Z�Ah��~=	��¿��yb�$�%�8��8[�g��7���M���y�S'��m���`�����j��
����q�=�*	��`���i�
�_DEHG�rm��<�$"7σ���0����z��A��D��j��� ��������PzyٳLp9��������}�ᇨ�xSl��h�m0B8d!��
���Z��Dw�p B�F�=:.?SV����<��?�fP�4Z.�Ґ��G���֟6��'��4��mmy.,7+j0��ϻ�[�u�f���"]�� Wx�~��X��V�W����u�,��l��Th��u��=����}���K�Q�jU�e��o��~?��vщ�;��%u һ;7�6��'�s9BD�h���׺�߀Z�h� ч�SI*�Ck!�F���#V�a��"��;�\-�Bh���՗�k-�9��s0�8;���{�����LJ�6���о-��x)�7�QM���*o��{�eYF��QXiB�I����ż_ �jJYI�Z��^'�iA���m�+�#��MC�ާ�����0l��j=H�Wz�0���$g�l,-�4o���۶�s��x�8v�'���=�CW�ﴧ��k����Y�}����W~�9}U,����:ytY��23�h�6��x�2��G���ք����W��^f}���� i�W����K����X�3��ln�=��&�md`Y?�0��o( ¶{E�mo[W��`���3�/���	��2����?�4^���n�Q�WH�	����K)"�D�Ʈ`B�4gŇ�O���xN�k��X4r���~�k]��'�:a�T�E]�t���q*� (V��޻�֎� b��}\��?�[��a�����6����$�Mf�]�K ����c~�W�=�4�ţ�]L��3�EUQ�LnY��s�Q=Y��E�N0��6�� �R�B�y�;����؝����anCS�>�f~��ʜ�y��]��%��R�%����D�5��9;�~��M�(�f?�@�Lw��ٺ������!L�G@ f��E�Mjo�P�Z"���I'�8�+�����&hzV���9� ���r$�-�RQ"�an##�Cw���.��u�t���i�D��	�L��!��ܦ��t���}>��n�g@.�B������]@�c�8�v����ЎR4s7^Х5Q��,}:�}3���Q�U�N�?��-H�Uo��\ί�8O(J!��h�8��T��y^y�ڐqV�*$_o8#�٦�D�5yn�e�h��'�viŇ�p�ߤ���}Gs��г���LBn�AYIW��ic��l9�R<_�	ZeD�M�!�Qf��5���v�p/�^'ˢ��=_�H���a�_I��I��#���i#Ev���;�GZ��3�C�#R�����
����>���|���)�#��N��5���x±i)�o�_sOt���C�ER��5��e���e��w&�b_���#�Ѻ�����}���p����ee��D��"���Aw{����I����Z�-,�=���ĩ��3���z�(Ohc5jƎ}.c��O����������O�d=a�\�զ8nH�<�b �A��Mf���G}W�<b��$��5��7�u����'�\y֜�>m�/�y4��x�ч&K����C98�8Ifz�q����5��$�3���}HUa	a�F���d��氘V��	sP�����%�k8���z0A�i�Vs�{L���ڙ�JIszq��8����TZ��W�Q{�_X6tQA0T}�=��3�f�����P����AMN��+!(,P���A��p3 ��j�]6q���I����K�g��ڔ�vfw�����%�^�ų�c9�Q�iK%��䔻w��<��r�b{M{�.��pG�D�:G~+� ;}�Ϯ���� �zV�����r]Ze����"E�}!l�KYH���0d�q�w�F"�.�n}�V�0���4�������@�;�<��$����ߚ�^�PF�/��l><�t�i��y����A�0�J�ɀP��k�ׂ{w#^����tvuHMY�^q�`�[nBJ氶1�a����mP�}�Y	��f���\G��p6Z=G���9�+�BH�*b�QƯBq�;T���9ԃ�����	d��\n<��}v���~O%���U(�$vH��:>�L�MQ� f2� 0fr���q�+��V�ѽ�%7� z����7Dw���x}�J���>y�R��k�KV���.����a>{��~�AA~�u-�|��7�y���6��wr}� ��r�n�X ���ט��_ct�}��C{������>77[>��z��;�6 �_�<u�jɸ�C�3ؓ��x��W/�4i	���p�ο�OJ�o�赆]�HH���/&&��-k@������Aƍ�vD�P��R�\n�I0�BnyH��)�J5����YgK�t#��wy�X�$6�rp%���:��͍r{v��԰Դ[��9��E-���?X��9m��B�wb�>!�H�e�!�~�?��+y�����O�C*�Vd�A�p��tY� G��vd�pAg��ϴ��]t��&Y���Wc�M^Xx�蛌�@���9
9�S��CW(�#�ݞ�2pP��A;aJ&˰� ��z�����;H��YaId���Ƿ�ݲ�p�h���VaeҎ����_��D�&��o����m�A8(̷ljj��V.��y�n�J�BKs1��<�AҘJ�O桬(l����vu���J*S���Ê��)�KܕB��/p��緰��w>�D� 59�4��������rw����Cs#o�1�D$��s|�Cۣ�-�.b�Q�r�1�yQ	b�ߍS��뾋��;���}���r�����(?����t�?T5�凚]�5GN�)P(53��&l�Ȱ��M^��ߦ˽��#�q��_�Ƿ���m#�ִƱ�;�8� ��WJ,&�ר|\aB�_#$ g�Y�A )4PZ�<>�( ���R�G�m��y�yr� ������犸�W��B�  .��� Z�� �T�t�v-@���~���#b���^T.�����qEb����bb����#/��.?N�Ŧ�V�*F���{<.��1Hu�[���N>f�Y�T� ����bW���.s^se�� �j���c� ��� �2���X��cp�r���ϓ�	�H�ӗZR���������l=�_`߀��cVVR�v�\re]\؂5&�^(p�#�܉�������6 ��Js���r[��r>|�d���uF���/O>��S!�'=)�v��~-��$�&&q �-
�D R��b 3���5�}����I�|��q��A���.,�}�=;�v��5E���>d�dE�UN���U<So�Iɯ���ǽ�Ij2剂Y��UA?'��j��
����Տ�9�QkK��׏�
#��[�X'�|B�틧�:���D�Ս�����}�R�>���s���?x�7ZN��'��-���q 7�����Qi`)��,ǟ�?�w���98a��[�bB2C^�x��dk�j�|[7�����VV��Ky; f��|G��*x;7ɡZ�"�/S��17WCL2��QԖ.����o�R�<Ju,�Pv��D�y��;�pb��c{��v�O�D�é�[E��	��9��~(.j/�{�%OI�ɻ�����7�s��a����J����o���׻z�l��ž��.XS���΀Q�R Y�4�@ӟ�{&�[�Wx� ]�^mG�Q�ޛ:� �'�7Ϻ�<{����f[���&c%U�>zV��N�AX���b�����f͕U/�궸Y���P}���!���z�w�#������F�e��ԇ'$?� ��۟�v#� ��PB1p��.�n@Y��E��8BTP[s����慼�)c��겦 z�#_3HV�����[A$�r-w��a�H�sY��,u�� �E^�8����f_�\2w~���t�i#��-�VvΨ�*3��l�(��T<���6�Gy��K���m���� �`�:v�Rɴ�_��˺bчhf�P'���c��:�ʳ�����XL�+!�n�pu��!D?�x��[�2 ���t���1�(���j���S�JL�+\�&]"�$J�P�[.\D�����d�����3�� �'2��M�><N��31<�����'�6s ���� �$�L�ŝwKK��'j�RA���I�RpT��#�(6� s#��0qb��3���U�W&s���@`�H:�#T�7RKW� i�[�CF�N�{�7�E�S6��4��]��-42+$Ў�h����.>f:�s�E�m�tÛ�Q/f`L難i�8��nP�yd4�#^=Q����6=�
�'�H� t��X�h���v�F~��#�8t�������ӎ�o�m;RI��2��fR�H̠'aE뗍!�9&y�#9p��pY�+6͝�8��J[[g�]:�: 2=�q-"�C¤&�`�ɡ��}E�NÞ:Y�}=r{P��s��Q2��X�8�Trs�7�T��5���Y2bg34cJ�8�s��ߖe����4��B���z�Ph%�4�4��F�H xi7&�p���K�s�_`!&���>dc(I�'�`U���k�9�<��^n��£����9��b��
y�:�l7����`
k'���i(t{"�=3S@'�N�PO�Kr�S�u�_��+���	�$3�PB��﷞R�xRP1�1e��+;I�
D)��6�a�:7>���hǞ]�{�lo;BI��\�VW[�d��"-٬g��V0�Ԟ�L�(�"��lY��L7m)#S�N@�Ep4�1G��k�lw�d���oCF
�0�,��}!�~\�X~�X����YS���t�*����kOj�:t�>1}c��a�/�fi�)�X��������0�	
2��t�4k|����湁ӽ���B.KԖ��e?�Ҭorh���)#6��Jv�E��,����Vc��Akp�QɆ��3��P���Q�٩aiZǲI%Y$!��!�c�!��ϷlH��?�O��-P���3 8��+/mM{�S��,q�ui}T3��][�+K��g�_�d
tM�)Z	6=�#�����?�s�,�U�;K�<]Y�S!�����$*�Y��l��v���s�rs<�����?�'�-��rF�GGG��t������fXh��8�k;;��������z|��g���6Q�3IFx@�_�U;'�[gV����ju~WA�����-����� �F/#��.*��&&L/�ʮ?��(&4ȵbhrLzB����=p�l��Nj��!PF5#E�@qD3/�В႐�pp�XY��:������3w �L#C~���b���� bX�Qh���������Z!XH;g�X�RF��s>�[��@%��|��4��̫��f�~&��f��Nd��Y�#[:|�A�%}�N�=;��%���;�7��ʆ��}!އ�c�Gk��O;�V<,(*y{O�Q| h���%���������,��]xo�!���%P��<K2�25�����m �Q��)~i��)7��S�	��aQ��������P)�<���7�Z���������wAcm�*�ۆ�&F�*�M�r�/�p.R<~���q����P4(��~�eC} �xl�S���+�Nt�����qV�Щ���Vv��4樠�5���;�_��j��{/UD�6�Ť/�)oL��]/�FRH�G Bc���X�W�fѧ��-�ג�_(�*�����w�|/�&�zǅ "I�p��]�fz���s�����g����q�6J�ڴL|�n�*"0��sX�c#q�)�(C�.�ʁ�r����O��0O\6�Vݾ(6��6�x30��y׉G�8�Kt�}�q�$^�''+f=����3��:��}'�>�p�����ޝ�ƅPM"�/.��>'��g�x�xf��.#�C=("N��,�q��X-)��DF�e�'��ea)��)("��!�������$Lz��=�׵�G{I9�b)�����E��
k�_���	e-S�C��^����P���IU�:�6�Xo��]ܪ*�8�Ya����wB��"���@}(�m=��M��W�A�@7��`׮,7�Ù��r_�2���#jg2M]��%4��.=�l|�VU���e����v4"qh�Z9�����1U��R3��B���I��8B�<H]!�/��u��Z�>/�x��O�l�\���gY�x�"dҜ꾭1�-�̉��q
*�1u]�i�ix}]�"28�Ά�zi��92�Rx {�ڪl6M���vZ6������\E	�4u��Ѽ��3-�����ص\�C3��a�맢���d����n��Hm}X�ɵЕh�aVLu�}�NW�g(�<=ul�3bE�@ �EB���O.��Y\Kw���kZ��	MO:�|�u�LĐ�['�f�^��ǎҥ��-Oں�S���X�A��К�D�0��}e�J-ʖg�A�g���$�Nܺ1l-
��3��QĤ���������ͪj^����o��zӡr�sx`j�>�u���t�ơ��O~��۾/�vLD����ݙ#�a�� _�X�McL�tS��mQ��]��Z�~� E
k�]İ��63s��ў��W8n�yQ5z�>V !$��ތ�o�a��a�پk��L��=��0�ʎ�σZ_G�`�a��W�E�ʷʠ���3_�#x�*��H�1O]ԃ]4���@�!�����x���-	a�bO\CcjQ�ij��<�&QK�gH�\N�|���M��Ar#K����vA0 $��\�N_�Jj��Nĉ=�W��X9� p��j�.dg<͓􆹚�=M%�@�^;����D��h=%q1�Mx¯c��}[6��zR�쇇�c�'ka�*�_����m��%�C��>�<�~u/.�B<�Z�e;@�</� �m*?�)�}Jt�Sb�JI�H�.���_c�B��;��a�����b{�����e�:�%k��#��G��*i�hˆv���`�8��?�V���my�����qGt��S}˃�J�HN��+�}�
g]�֢2uQ�^FV:�gV��5鋶�P)uo�D���e�A�����F�HE,��㗝���2g�l�rI�!���0=�3�����nJc�������1�s]:���	���ϯ�\�>���D�c-�� ������ȯQT�����/�j�U�����ite��I!CuM�:Et��4[l����5�4q�y��R)�|u�i��tS�I�Lq�Ak7MM�q�&��\�?ќ���T1Q�d�e��������d�m��JI�!`t��X�<������|��c��"��D�%�����0�m��?)��A�i��ZXsA�͉�G�����t�w��H���aS�����ڎ����i��a�K �������	�.J�+w Ic�M�hj9Pj��l��(���N����d�5���ߗgm��� 7�fY�=�(bM�>K���s�)�2�y�$�g��B���)hZxq=D�J�,Ȁ�5��h� �Q�<[�$�2"�j�| [�%^E� � S,#��;�E�qυ�h��c����R�@Q�WϞoA��˸�m���V'�0�I�n!�Qo���A��@���9:���C�;��9�#�:�4`�}��s���R�Ԓ&v�;���*t��%oY���,�����S�e�As)�����48ɀ��A���������71�PVe������:����Y|��>�j�H�^�c���>(O���0N+D����AB0�#�pv5'- �d&#���?�W�H�n���m���.Y�`��o����>���	�X�m�׆�bm�I�$Տ4M��h�����7�ax��W��︫m8:a�����ih[x5��p�`��'�3y�P�$�pE�(1�~3��00���	�`��W;5ͥ]���t�!���K'rfb�}�	-zk��e�6R���B`1B���s��$0 	iHϺy��c�Y�ɿ2���[OH��E�{%	�QP�f+Ot�����ۧ	5�cPC��r��y�q�O%7��2���K&�x����ŊR���uB��:r��Ư7�=s��K���#��jo���a�@��-XS�j�~�1�����r�:v�*��>�%��s\����RS�T�"�|�>��-|�:e�)�C�A���2�S����&��E
˰S��� ���&�������\�~���K��HՁP��"���d�p*��h�����B�}d�
ԡiK�; Քq��m�C�P���\w�>��N�u�ʫ�>6uBX�?�Ǻ�-��6W�6��{h��Y7�mRY� 4�N+��#I���M�Y~DJ�岓ʬC�&��>�,z���J`t-�F{���w��{>�0���aD �bU=� �g� ?@DM3��Q3p��
Zd�!C����/��4��tB<	�dsu#�3}&'5}^�k����_ؕ~r��f�pv�H@;|`ڏ�a]�Һ��x�����(;V"�*"f=��2V�;n 
;U<j� �Yx��IɌ�h�7��5�7@뻔Xei������ϯh�+�
&�\+M�b+V�tS�X�²��$6����$yTE1�&�Xil�<�$�c���jX�bͰ)15<]=Z��j��D|r�!�h�Kj{�F:,hw�y븖4��&E���4����-I@��6\x΃B���:<b
�����6�L���^zݸ`�~����P'J������}
�l��)�Դ$FF�%�@�2�~�$�WК�(:��]3b�����8kA�Cc���+��`���7±>��2̐zb����*���;ߘhF֏>��LN��6�]���/o�,�wSm
0��~�BĽ�E��q�P�'��V�C=&K���q��[p&V;|�` :�\*h,5�ث.�[<ӥH�`^}�x��uc��j��GM���jH��9Q$� j[�� 7�h��i����pQkd�dN�(���MTW���t�1!�,���L�;A�vV�N�QJբ(��!቟�lJ.��z��6�Őbrs ��I�dW#rKsW�K�$�c�x���.I�Tj78jV�i4�5`��Q�f��4r[��b���u4�I�5?!���7���=,�'m�ؽ!�:؎�.V���vTN�,O-j���#�N�q�j�v^h�j��EN'�Bs� �j���]%��)���!L8!��ƖH�IY�@�����}��-jA��=��Wo%����*��ej��.�Tܼ�e�������ƞ3��Q4��Fݚ�z\R���:Ö��.L���\3
�)]�Rw\\����1V!'�ל꞉S�5}.]��,�f�֟�+�M>�C�J)�{� k"/���@p��lNUV͐�<R��k����V�G7r�k$��"_M*�tcM��P�N���X$�.D5i�z���r�X
�A0#��.>7��k(BE�<�1E��gn���i����K"nȼ�*d��n���
��%�r͟	�%]BFb|f�AB��PSM��Na�>�[��Iٝ���Hp�-��(�xRcj:�����/�V���K�`+7��F����S�$ʖ<���?3��Γ|f�:�a�ْ<\r��H YH�a����N=[pf�=��Zo@�t׌3�g��t��B�����g+Ls���ʎ�u��TB�F]|�����r��� �V	�C�Az��Av��؏i$��!D�b�pزyM���|��|��]�����Rfd�V��h���i)f�>��|/���=?�`����f��i��o��y�d�4�徯#M
}�<����m�$ܱbi�<���]:)�-���F��K��	��g?��<���M�$8al�9����0?��3v$�L�Dm�%��N��+)g)�3s����~-��L����E�/���l�}���m�����=Xi�o�_U������u�:��_��Y�/܌��(�4�M�KNJY�N�� PK   "��W��L�h� �� /   images/40f7d2e4-4064-4959-8822-d1932a7058e9.pngl�w<���>w�޵ku*jTՊ�U��ޣUTc'���(�*�V���3�*A��J�#�nl�+���<���>�?��W�\��:��}����>��bf�� ���h�@T�����G��T0C-5P9�o	��ָg�o��E��x��l:�`�������ݧi��44pcy���%�S�C��_K	��U����z���_:Lq� F1~���_AgC�̀���}z����Y�x��e��)x}B�}��e���y���j�N����y�-�F�\�� �[�2D����T���H�<��K��*�o�<��������������۳�_����AE�L��_"�>��۞�N��o�;/�?WAM�{uLy��l 	�ȡ��W��W'���Y�>�J#B���ʸV ����@�[�{$����
��L
����M�f�3��ʮ�A=F����:��G���@���-؟[V?k6��: O�U�9|��R-��+%O��y��h�4ТӌZ��K��KC��Յg�Kf���ՌP3�)6q�alW�~�d��y|���{�~vKV��f��u�|$r��Kޏ8�d�OH�G{��ޤ��$�����fD�1$|�݋~K`*�1+-��`��$�_x��˥?4�Ze��i���5����Y���w���F����M>A��'��A���_��  �r-��;�R�B��V��
[6��5�&��^Hȵwnl*:_����_�nL�y?�9V,&X���E�������&���T���	L�q�FG�wˡE�4�
;����5-��M��l;
����:��Z��1{M��)x͇�]u��*hQ��/�'���X�w5��V0J�J4�~a�]�� �DҐy��X��eR��Y'� ���9�7}��3����k��Η�/2_g�j�c?��ժ�&�D\�X�<<�e���S���8h��m�H���ҕ�i�����L.vL�$KjO���e�px_̓xݪ>��=R��mUR�w�0�����EJ$ݻ�ZI��K�w;�un��J�Ͼq_�,�Ps`��+��bt-�j���{�$&�B�?n������{��A�(XO�`=+�CwH5h��C��9p���_�E�<�g����mR�&�[pZ�]1s�.��N�~�A_��ז\���^��w�ϧ[r~�;Λ�_�^JOu��8�7�p���Vƕ���%�9s�W��T�f5��ĭt���ؙ���V��q��ս��v��p�e��t�xX�0�^�X.�J���W�:�p-Qiv��԰��C�.�߲ Qg�M�����~�kӫ϶�:�j�|��,@mn�^�����S�m���~�^M_>��φ�k,���u���"�Lh[{�RӌrTB�����~��
|R�(��X�W�9�F�S��3;�ퟪ���{�&S�)�VV"I�ӂד$5R�n$��o$���|�t�9������\���x�u�B���Q���������W��F��@�f=����Æ�Z��R<��W�I��\Bh��MiVw��#%+��D�r	_IBi	TD�#�n~N�����8�r)���,VX�%#�]�*X��fld���VM,�JhY~���TxM���ӌ���z���'3�X�j�T��r�pu5g9G�0@��n ������yv�Y�㓣��`�9�x>C���7�_�72��~$�܋���4��Ҳ"j���49ZYV�����[�;9Eb����q*G:��y^�<���i���L߷�����P\]]��p�΁;�~!W��D��74�B���>��!������(�?�JGk����sz���@�O�;�i��4��\[_���["�7rh�E�[�y������W��|q}.6l>�l9R��D_5�0���u�mf�m�F'�Ќh1��gu��u�j��]��f�f���9_n�޺�r�N�!��	]3��W�_�۠�G��Qn���K�{���:iΖѿLU�L;��͑'�)�T+kX�W�;::�>R����|T.ϞR�eMA��?�7�Y�9�ߑl��vD+��X]L�e��z�@׵�\!�q�S�u&q��A?'8�Iz��d��O9��Kz18=є�k�l��	��b����ϭ���Ҙ֙��yjG��C����ޥ���y'�i�L�T(yM3�����ύ���JLdD�2=:K��C�>�Q��Id�Rë=�� �rs��ĸ���׼�--�[���~�������{���怜 �=�Ԧ���w�p6��k�2>}M�n<Yy�ۑI\`�Ig�Oӌ�i]�C�J���z	���,����I�ˏ]��ɤp��j(��9��p&�%G�9��$����.,D+Ѿ��^5c�
�V��16B4��咟 hf�x�D>^��s��Y��[~���P��f|�|�r��r���oEE��VW�!k������m��4@(S������;C��#
vC
|� ����*�G'�.�>��Co��3�V�
1U.S�Ə�	Ot�Y�&������������D�@���i-^�ٟ���|k�7m�vDF��n:��$�	N�$i}X`3����G�\�O��Wy����#��gw��� ����HI����ߤ��	��p�RW2�{��CϾ�ڒp��q� ��a [y�,MJNϢ�Y��
5x�i���L�� ]��%��,���x���i�:7�S��w�PHe��WE_�����i8v�4�����ɦ\}�a���E���@a��$��A��X���y'xv��mF��㬃��Yh�T��o�QMz]��X���F��q-��8#˽��:�D(Ɛ�<���'�i���a�/�A!��c�׹�M�>zM��h Z��&,^~���u��ײŁ�a�c`b��2�K/x�ccW(&�0��K�q&�9��Z.P��CN�yU���C���En����������uqܤ�N�u��zT�Q��4U���<	�zi�H.;��4t���]
ƍ(֓�2�'m���F{pȷ�	�6��K^����!� ��������
�h�3ળ{�*�	T�R���'�[�޼/���
���o�t=Rڸ�2�K�����V ��69���t˴�qjp��'��*��7��t���0�\��N�@�t-�U��U��n?x%zm��[�����Ϋ����_�a��x���v4�WXRb�Eh�z�|��y��s���y��F���|���I�tլ�/G_y�S�!7r�Ȧ�|(������XLh)0����`�`x��*���6�"��t^rQ�`h.Ȭ��b����TE�uع�k-�~HE�l&އt�I[l2�k��� ���ӂ��\���}��>7-M�%I����7��$��	�wR�/� ����ߜa?Ed�,?��1�/*he Sb�;�M��ݚ��� �u���u�����Z{�Zq�=9:����O���P~@La:<��-�����v7{;�32r?|�	s6S�K��W�/;jsԏ��Jݗ��Ky�a*p�,���gy��T Lހ�E;�]l���Ux����@���}�N�Μ\㻉�.��a�i�A��X�"�t]���g��nX��r����(�5(���O��}��78v]=[R����X��@���o��!GkS%f���h����o�
t�J�{��e��s`O3���H��G��X#'yHE��������#��fC�	�0`(y������w���@>�<�����AV{����9rS�^�E�Ek?�tp��]O��HXuIXl9I_������#X� .E��S���]Ca��e�{_�TǞ��7�clKń����?*�η���:[v�#�0}� ����bP|0T�*rč:��7Ii���b�Ȧm&���U��J��GF��D/���nN�L��l��Wd�R� 
�`O�_��e�㤼y�����2�K�j��)�����$K8�:�\������A00���g���<�q��3�"GQ��H��b��	'���&w��T��\����z�L9[rO�}�	'��)��nx�uE�ˋEž��b=�-C��i�F.�(�!唫7��{��������#��F.	�<�M�Ԗ�q�cz��yMM�W���W��G����&<П>}=��&��7N���-�+�~���ߑMRq�kz!Y���I�U0�t��Ǉí���FR�g�r$�K�E?Z����_��ӌ�م���E<�Y��\Ǘּ<��Z������x���{����M�AX~\�`��;�X͂��a
�(-E�O6�+�����������e�:�m
��Qd����j��&�9����J^��d�Gd$8�+s��cߠ�Kw]�+�%�͟�;�Z�֢<7�>�z7M𖎚
��J�n2)�6�T�����@x�p�&��K��I*�$�d!����ߢ^��%&Hcy���H�Ax]�	�^��X��=y���	.�&����h�Ȃd�K,�<>SY���l��X�8�G������������۰���
I��0�;Rѣcjf�&�T����%͓E�vWr�M1�(?Cj�|Y#qV���Wts�a�S��"����K��P�4g����NklZ��\�h��M��E[�Swv |}��Jζm�է��:>��%��U�͸�iޮ�%�U��J��/n�vz��~�����a+����u�6��ܓ�ym ?SP�\d��/����0ܴ�s�e	������,����"F ��C}�H�?�,��Q����)&O�%�I<�J9���=�A�N��7 ��*V{�p^~kn��꒖�l�۔(ח�/�?dxï����p�4"�5��⣶�2�#TI %�iģ��(k���+,~߱�����?��5����#�m<w�!`2R�Ҍ�$l��v�K��~�==��WWIa�ؿ�3(7}�0 "����=(?~�c��GXȶ�Eg��p���'MQ�|�ʟ����24�>��&����Uk^�K�[%�6�7Zp��y�R�Y)6�S�W���;�p�Gfv!>��g�`R�J];or���l�3�=Fs�)�@�j~%�n��-�w���%�����Mt�b�7>��W�����ebff���x�OL�4h	�5�\$pW ��B�����h����D������ru��[Y���,�0��pL�bu���'&,�ˀ��L�q	��	s��k�kv��R��,,4�V�7r��C����>�x��KC�c�<�͐���=�+�vvz)N�[�@p������$t]j�K����u�V������B��K&|T��u`�:�*.*7����%,���&��?#�����s =��l*h#���޷�ؤ��!��0v�W��;�/ۂ�y��,M�d��se�҃�.1���e��7�F���fM;'by�k�M��T�?���a�~�1��=��~���[�ױ����7Bn���B�Z���r��o�c$`��[pe)=Vg)6"�!�WϨBZ��3�ѣ�ʑ/z��P���(M����:/h�D�*�ʸ�<���>J����%^��b �0�W�9�-��o_{�;���A��&�1 E�Y�{,��H��=�AXtMe�����Gy�Dǝ_<�����X�ǐC=�f��]$Ou�b�:6>�A�R@�2�i��4#�����=�����7!{�na�'I?�)P�T!�re� �~7W4{���V[WƊ��z!أ��������#HEy���������e�Hz֣�iп����b4� 7E:�U񰬬l�c��lԏ�r����!u�X�����$nP��#q��xz, ���$��y�v�CR��¹���'����@��U�7@<`�?�Ok$&����j��Ŕ�ʹ�.��I)0��_�<�s���p����5�I7<8��^���ku\>|&T�E��;mW�7O^�!)פ۔�k����RW#�)��\�%��C�ݳ}'�[�����g��9��.?��}��>�=�wĩ��{3h;�}y}�
�=�cQh5 pR�m��[����@���d�����ۥ�ન��~��moE���$������s=O�`�m����%��O�_��{[e&�?=��B���é���N�
�������d&7F`���(�Suu��g}�YWrcn_|W脿$�m�Q�c�䈤pw�\�}���"�0���B�ݨo*q��-yo݇ۧB7<wg�g�u��Ph
d���޸�v�r���zS̶�\����ա���g�����Y 8=����u����˺15td�!��m �&�m�pN٘S��1Y���I���7���l���˖7v���eUvn9w�`��u�8npG�uDꗎ��Q�8�3	+����j�6��hWNs�V����u�#R�D��������/�E�[��R�t�C�������>�"	� t���#�47�.��e�	ʊ)���Cxt
�Y�����
�T�����KIg~��g����(z�z��d2��.� ��k�����"4��� U��Ԭ@�؆D�T����k��"T���1`���c����뵠g#�c4��,N=�;� �� x)Et�W#�ۈ2�=Gh���/>�b9e}�@���+O��}�(x�O�T��kN�}�>�!�ť��n����i�2�7�i���<��QMI���M��uN�	Do�]4�!q8�g{��
�	�1�����Z�}�4��	��f1�����E��/p��|�5�zד~ΦK5�b�28����tME���%F�B��0 ��4z}c�ݸR\^�h�sI)����'��>@��)ߣ��&�%@־xG���3{��g�)U��5Q_�	[1[��tp�"�m���mkten���nhד�Y3U_�Ȥ��:bl2����?܋�@���S��9Rwu2@�!�����{a�������՗ ��GQQ��do�~uM�\��{��Z]У��g�C�[`sx��~�?��~Ѭ��?�f�Ҙ������p�{+dRn�v0Z�C��@6K�!�EZY�P�zCR�Z����t��mK�u��R���oa�Uʤ�{��j �#�⃁�ƌ}[W��*��7X,֗j�Mcp��Z������V̓ߥ�����5�:�%k q�����-]*�%�w�m��2��4Y�5��@���܊h0��,���d9(����wy�ɿ*��[��|C�GN����R�� �K	���Hи`E�����"C�Y�:zD/C��i��}}��0G�u�G��=A�Ię��17#k�QP��0�Y�%�<���Lngy��vƛb�ӍMUk�u��l�$`5�ܯ����B;2M�r4��,��Li��_�V{�O����hG�'��,��p7QW�
�xdT�2�mr�Z��%J�z�|H�źX�)�ll��G�D
���G`C�dj6�E$��Y��#�{�c�����Q��c��~�J��ɀm�������|#ak�w�Փ'5݃��}A�^��cT�m=�A��q����n��t�m�Z����>>>Eٲ��'�3s����tTV�SB��0=ȁ�E\g5��m[
m����*�V�� �Yd>�P���Wp�kӀd����D~��� N#���9ZPS�
41������[1x��������#��6�ڣ�`�T�ms6�Y)�AS�:7c��(��$��Lp�_��_��R��V�`�w��JW�(�k^nm�P�^I��ٖ��?"TUG����6��蟜mh@F�m�|���׹%ܲK��&�����1Q���CV�~)8�ѨĎ F�Grͅ��V8l���0@���{�?�,��E�N86I���lCTh��)g����)�Ր��l��#Њ7 '� �\?��o��t�p��)	.��a�MZ��9����C�j����ak+E�;��Y�K&��У�
�09������tLIGI���G�;�� B.����A?Cf@b�޸@��A`�;ԝˣ�
�W�M0w��*x����-=���q�Pr�^��
�b�\O�����ޔ�{3L�E"�^�BT�)$����~ʉ<�6;�p��toȏj������Ŕ�q�NVz�������
���-�Ղy�H�m#�;��2�8z��f|Ǭ��$y5O�1�r|BO9�V2���%8�I>�9��EW�;�������gxN���Ct�-~�O��	�1�	������	@b4Y҂��`kd�9b�?�D~c�7�s#�j~f��f2p�Ξ-�A  ��🉠���)JN��y!#'w���w��k�^^=�2�]F��HH�R,C Y\��X�D�z���9x�6)s.��l�~�uvS�u�;�Q9����aG	�_��ʲ��H�%�V$|�p�qf��d�g���@���~-<�H�uq�D%�7���6g�����s �(�?t�I3�V3��\��Ky��[s��%�F�ʠ�x���]ջG�,( _�h�ȯbR�Sg$��Da�f=E���K������uϮ`8�pyF�/��P$߲�#��}�~Y,z��xB���Ms���'4V�N���9Z���&�>���5����x: ��*ge?x�"��7��|Up%y�
�[�9HtrE��]n�LUq~Q|��'��6��D��{���~��ԪTT��R�Y�i5��"�O�<
2v����]�_wWQs�i�{rv�RE'%�(���E`j�?�9Y�O͓���)�9U�`�������N�|�]��*ZO��z,e&␥� �: �C���t\3�ʴ��<�{
�!Ȣʺ���PMU]�x}�r��Y�y_%����t�Y�[v	�UX/u�r��I�.��ժ����Ѫ9G#f�uMA /A�П"���T����$g�.��hř*�x�j���Ò4n�m$ }[�t��+�6�%*��շb���o
)�2�W��6���gp9��q�	z?dgЯ�����\��0]n#��,ڮ/�����+�N�p�7�Z�L�m^yrun˶Yg�+Ic�\-�)7���wь���p�̖)Z��E��yK�A!�7�i(�Z���i9NUܼr��������9�p���a'_]���a��ܧjw +M�Ϝ���q#{��q���7�-j�}�F�UG3�u�5y�+@ǐ��L�q�n?�0ȗ8Z�ӌ��kV�݃\���ҷ�YÕ�����"i���X;!�BMjI\�ω�\9����� 
!�^��*
{�W��	����<�W�0����x�3o���t��㚮�W��	SQp�]Ĩ�]!`࢏���>A�G��?J�����n�V�h\���c�}����Oֵ��f�v�j���^
s�s�9�3q�$ZO�6�l_����ū��,��C��J�λ��-l�@3	=+�kf�1����b,���J���y�I7�I.�g�_�AZ�q������E���|�Z����C�Ξ�ʽ�Nm��Ub.G�'��?�����}qR�����p�����u;�&Е��+h�ͦ�Bw/ōj�GF-�к�[�6Z+!G5��������̝��L�N��Թs3�HLp>V�J���\7��Q���Z��-7�,��V���\�?W�)���Z	`�9�!%w��E��N���$�0��5PG
�V�H�Rl�Z��e���i&����}�FX��z��ޚ���������)ɦ�7hqtb�OH����n��j�X��#е�T���E�ڢ�W#��eW�8����>�RV�Jl݊�4�'����Iѵ�Ľ���i]�y�_eP.ъ���s���ua�J�����]{���w��֍���x�[�K\��m�'jʙ���΅��K���V|�+DZ� 曻�� #���q" *	�b3cӐ�)���w��� ;��N9���=�]!iY;w��	������ۛ=�ɠ���k�x=w�:����~�S����`��	����$'��g Ɍ�[�����
�e={�F\/ʌ�L����{ P�S�W�� di��ߪ~j�.��p@��</��y#%3�f��sٷH�tIkRȼ���<�p���Qf%8
��
����2'9��X,,���IB�w�lâ����1F3B�p⅊7�)�&�Bz�m�?�U��FGMe25�Kų���@�m�F|�$��^$�y�k�'���2f2d41F;4Ri��=�_=�z-�ݠc�K��)�����zN�^	ʄ/�ο+���L�e�\7��=�Z�i`Syk�������뎏�^\�u(���f\ǫ�8���f����l)�v���f{?�,]�`}�h�G��79=�t�Hw��iH7(�?�t����ڄ�؋)��TP��򣢟�̺�F0����(�Ny=�C�b)mpo,�?�5��1|9�4�0q�h9x�^�{+�	.�/!p��[R\��C�F�ߧ[�a�?VfT�ϬL��>;!����_���~}��(���[r7	W;=�H���٧)Vɱ�n��
�:�Έ��H�o������ ��U��h��<H.��$e%�pR����I�\.�`��)y�>/I��|3�W�a����*���9�C��f����-z���?��/O�%�V��ˣ�J
I�R����} x�����0��G�%�G�'���o/���*����;E,^��띉2
n��4]�/���E{ՄL"��O{S'�ԷޗAB*��C���U_svac
˚`�S����#�/r�[;�S|�|���ʩf4���N^�U��M�)���X�z��t��	�@q*7��%p�H7�TS>�26���<�-9�(=	ܻ�+U�'E�W� 1o��+�:�����R�w�jv�������r�Nn<д��1�2��py��g��1��i�E��{���̶i�M&w�.9@���~߱T���OI���v9a[<��'1�fh�x�B �_���X��J�
�}2>َ�Գ��� bx��W��ǧ/�.��ߙī���4L�1����dq�Ç�ϻ뇫O����@�665����9����ihT:
�[*��7�m{ȼ�y��{8�c�Η��$B�t}G��Ln��-���B��A��|4���`��35hH��&P�>������Юx8#��V����m�a FĲ��"��A��#Ii�p�Vd�o������p�5�C�M�ȭ���r�Q�pk����P�j�n`���v����I��T�K��vT�a`�uɋ �f���U~��@�ecjf>s<�Yl�F�L^���߮��j	�=/��oo:p�=���L����!�M����g��0�Ѕsx7��k�-�S \��Ŋ�qb���A��=7J�/�����ȣ�?"\`���r�p)ܬ��N��{V	�*��Q�ȷ�ܕ�Ȼby�?|�@�'~��:�@>�_���kD����N_<e�����o���1�\�Q`8]�z��'����l  �:w��;F5�!=0(U�ZME������*���w���5���?�+��/�oU�*Z~��x�J��΋Rƫ-�@�M�F�CZ�FyrJ�Kx�v�S�Řʆ.���G���s6��Fk��'��k�s⎹�Ϛ�+�gE��c���y�����	�DE���(e��oZ!������+����['�D`�+M�Ƴf/�˲��0~�v\�	��4sL�r��� ��W&�9��{��w��DEcY+va�D4B�1�y��՚!wi��E��b$�4EP�b���S�vo>�T/����CD#|���_��
g��OEn��ݶT�C	IuJ��˰��/-O�O5LL�r�����N�壞��`cpY�����H/[)�2�{#Sf��n�uqpz����Ť�Y��O���="�ܝq�hq�_�#�42�~Cފ�B97�KK�nj=�]bCke�gR�L���s�=����{�~Ǳ�;>_)S��e��G��+Qq���%����7�_@9z���>���323� ᶦ�:�M�����K�+�Ͳ����@3�܅��g�����6��/P��:M2	D�,�Q�[�������ܪM)��$(��)�N�j9�=�.۩�E_�1+�}Ǉ+k
��zgh�q��$����'�� ,��L��?�B���D�N����ꬭ,�	��MS��	�Rs砻��I��_���j>#VR����3�R�}n�:����~ֵ᧴?�߶���2v�B��x�o�ױP��Ū��|{�oc����菌V�>���brh�V�L_��,�h��%����*Ȩy��_tR��=��,��ťb^?�ֽwχ��&u���(֨1観�\5��������ZOO(<�GH܊�d#-�h�f���r���Q7Xڴ�g�M$�>�4Z�ᧅ�0����22��i�bQ[��r �-�������M@�W��9�q�� �qWN��v�ٝ�D����BW�2�d�5�2w�tLfm�Fw����M�O�����@ܞ"�j���b毞�u����� ��9%I��悁$a<�I/H�X�U�!{�����!�E��D��2k��J�d�Wo3/x�X�Gj�7��:��O�a�!nB;'�D҂���ۅ�X�q�ny��.�pM�{��|��U��2���G������t���J*#�Jk�Yl��rx��j{��P��Yi^Tne�<���3�J?E�Fm�S����X�j��3�_��2����Wk2mZm�A�u�{Phyeŭ6���$[��-��ltɅ�+6w�H`����j���ȝP��h.�%;b�FYT�E�|zr��Mwx$��*�Nٸmm�<AP �I���r�yc�8rjl���v�z���4,��%�&jP�K�KM�m�S
�aSp���'�mL�u��4-fo���
M2ӳ��j�h9�y��`�K&�<� �X-����ǜ����ѲCz�r0��8���ӯ}�p6N�*ȴ�+}���@�Ld6��ޭp���vΓ�����5�+��G�!̈́�ߗM���*���F���� �Er-�6U������ox���ҥ�Uڽ�uF��yўL�n�y]:1�f������2Aat�T�j�E��D:��fa�%�uیgWߐ���qhN�l�9��x�B�
�h?�O�H;nB9�e����$��Z�d�T=���P���`n�!��/ɸ��D@��C?��� s�,����qXY`~������)�����֦���?G��1����K�Oсاh�X�����k�Ui�B��@p��5��Z�C�o�k'_)Z�hT��QTI��S���n�ܸ��Ș�;tϸf^���t��u���Q��e���Ha�W��j%����ۦ� �<٤\��dL�޴�uxa }篧��ۈD��y�˰v��i�[�oL��yd;N*`�ψ�������#�����t�rO��ô����>����m���_�HT��9w���sL=d{@9�A�I �Ґ���-s�z����]� Y�n��D��K^{��?]S �=������z��`�ĶḶ!�x-������#��Qd���a�Lr�j����pi��t�df!�C�N@��Q�wYp�D�$-g�K���cp�=FY����O�J��IbķI���`�/���k[ә��_�T3
��.��k�7Lc�-�v�N<R~넣 ���|S�us3���y?�����\��|�S)�*�fOn8ef���`�J�����c�XDf���.��~ǩ���&p��6 ~3N���I�I��뀝�ɤ�;��@ƚǤ���&kG�~Z���Yw�SW����:	�7��a/3�!޴GH��� ��%�/v��iva;�i�+�}>��F0C�����ȋ9�3ᱱ`A�	$N�����z�A�R�a�YhG(��3v�z����T�nVLm�*�	��%·k�s�4�@y�F�e��!�d����FD �w�������l��h���	&�vĕ�;��VKHj�k|�8T��coq.!�kRȤ�^�\Rڧ]�p�ʹ�;=ΔW��YMLn��w���p[��cB�����0�m��Zvw=�Z���u%��Xܼ��-~�"�������e����TV���#f�(������*hbff�Vn3�D�>b�!�k5"|)�����he-#T���������rY�!�˶Y0�&�0��ۜ�-B�+Q��l��>��s3�V�YUbz��vx�i5�[Zh�#	;k��Y3~l������k����^�6�M����sX��og,U�<���ӟ��n9��T� W���E�D����msl��|���,P(�� W�����A����4h�,��R�V^��+?�P��X�|�$�-��X�dH�8�y����Fm��N����SS�&�ߟ,퐏3W��M����x��Ǻ�}�`���b}��cG_e��4��X���"�M6�L���1wPQs�^��{H�V>$�f@��" �v"_����f�$Ԣ��g�i��!�Ixv߱�9�������6Bl����,[��/.2Q�)v�N��0���sJ �MAd�3u+�rA�0_E���<���\t6�Y�y|���/��s��T��H~�Yq-Z ��/~��ߊ��>�s_{qʨQ��%��|H;��A6�`���2��eљ+(��D����D�t@yk9,q�Pt�-�s��D����}�Ԡ�����.�L�ϥi�Zy��զxY������[=�aԁ� M+���D�D��[��=5ox�^�4ͤ�����l��eb��o��^0��]G!��V%EE_!��<6Usdg_�[<�ݺ� �j�cT~�}�:����8��HV��8��k�M�8#���_=U1�	A�Y�Q(JT�b
�s��������;轒�!�v�˧e�m��u�H���i�-��R�8hC_�s��AAo�v�(��99�lO��-���[q�<4q������Ϛ�3�X��PQ�#S��tu�)OE>��=4�@Zl�>3l�Y���@����cmE׆�{i�>�ո<H.�L�C��v�m�)wp �0��bF8����� P�����7��K�1EU5��7([�8I���E�gG+<��{}�Ӣ_�ږ-�[�m�������p���F���;�4���̶蚖�N0pd��`� �ǋ��P"NZ��ޑf�qM��ď�se��ަ���y��&=��x��.3�����r�>���{�AtЛ� !!��
�Y�S��x���''�,��>g�Fu�a5�!�2C���&x/e���輏��8_<D�uG�=�x��}�[��,]�{�ǀ�_a���Lf��#�&�xu�)`x�qP�0�˗�y��C�KTIz����j�͸�0������9��9y᠓�B!�k�K|�4���"���^���<V$P���W`λ6�|A΅\�f�� .�jV&K���_����9�9����#N�)_��6��|����u��{�h{� �j`J/?˛/d�q�S躊�����1�����۶$:�Vݝ9�f�(�$�bnx�P7�<�T��t~G�r��M�/�Tk�kђ���m;��n���~Kf x��O�2QTpX��\�oû�$��O�0zjQ+~}K�)���I��:Ã�ae�mg\�Efœ�i�3�j<�(PS�6�U�����rT�m(�w�-����-;���<�>fN�޼6��9�M���󅋋�۹X(+�n��βû@Μ����P���:��8�`L�[�� ��T�g��m*����*�E�i�覍���C i�g�o�$������k�x�\`m��S�h�#�P��т!���`?�=221k��\�1�oZ��n��C��Q�'G$�W�$�I��oPD�׹De�/�v��'���%��B��ү7�P1k��xhRF��J���}` x�ܴB��%ede�����7띄�$�Rѷ��ф{�B[~5�Y����(�gUm�=/ٖǲr������{�
�%�ſx>�R�b�"��y� �A���=ʬa�&���!�hM�io	
tpȧ.:���q˺�L�-?h.[�6�$\ś����GG3��#1��Ɠc�Nl���uDE�����=UM�kә��"A�
so�T� 愢J�l�� U���"��❥�ܞ?7�,>壱#��|H��r聱&'{ج��[��%�7��f`ΥD�u֡�`�����w��e�{G��t��g"WB~x���H��D�����Xj�t� A���<�u���)��;��4[=���}�-���>���3��1�T@h���!k<�!Y�G����ͽ��8�&o$P��=��% KzŦ�U󃺏:r�l�ܻyq���f�\~tF���{�n�c��뺔u�Q���0���%_$Q�f5�a�ڔ7�#]3I�}�#w���]�oj��cB�}� �������~���ݥ5 ��$y�%�V%ys�u���7�~Tة��r�/�(X�5�����HC2z-?	���νү�����,���U����M�����i�g�Ґ��ۊ��6fj--���U�?Z�0���+֯�����yi��<;�V,Y�;�\�N��孑�Ht��?K�����5�~��W(�����ż�r�S~" q�_sw��(�=��5�>]����jd�2nޫ�e}��*��/��y�6��3J�1�~=77Fˬ�.�A�}�f}���.�1x���դ����'��6�ܝK��3,h0���d�G�K�Y��
��F�3�v�K)Is�c����S�����Fe���&Md��b��-��j�niI\�̼3�r�뱄F+Oq�ܖS�N�#���m���T?��3���le��D�`��!�/�#el%� ����afw��0���EV�ԹPl�
;��6�H�l�d��������,T�5����­Ɂ@�۪}�o՝��X��a����2푯�������>���m17q3͌�I��k�w4"�:���d�	��!s�����?e5��\|W�,	<�Cp�|�@pwwwYl��[��-�������w�}����TwW�Twf�)X�W<�v]�dw�]^�M��Hy���)�p�^��~	�XWݔvu��0>� K:r�3]��-�dڽj�(i���߱Q�tx�F��w��.��y�hX�V*-5���i>(ͱ�p��&(���"4*'�ņ0��(I�܃\N7[+��b54���zXr���j��?�k��8f����X���X�N�_}��M�'���t4#'��;r��k��Kђ��Xfc	�u��ل �xIGG�0E�3���>87�xޞ<��,����� Ҿ����Cnֶ2Vχ�V�W��6zp�t�:M��x,#
������k��_��!8�B�J���\f�٘�Ji~:��C�B�Z��}��-Dh۷]����x��߅n0��"�>��>t�b��TQ��@�� ���(�cT�Bs>�E�/۫I��2H�2���D�N>%ğF�ԇ���Z��\��t�rt�&`Ol���32��� Y�-�נ��0��(6p��nU�Z����&����#41N��r�T1�ʱ*J&t:߃��eH���κ1��s�joƦ���#d��%�=�<U8�������(�۲����yP��v(���,-,�^��A5 )�o��{D����6����q��;=�ΚJ�����=,�ܗ��y� W!B,,�C���Ws��
7�#�Kշ!vҢ�3D,EzS�8�u�]C�]�y;۞�a�w�L �k�,�*��-��M�{< V�|C�=z&]Ys���`y����,1u<#%���|�M5�J��d�m7ޘ�C=E`ٗ��8�%�@�V{�WX�l�fP�W��w5)_��
m"��H�~�װ�~U���s)>��QU�N��ew��=Vi�9.б6|��6�[�{!����r^�N�Q�t�%0���;6\FvLO��kZ29����(����ui��N�m(�h�\���K<����jj#ĠP�~}/���!5�v,�})K㝍�1�픔����kC�T���5�$B71X���W�>�� }�뼻G͈4���i�W	mC�W�uJVL��L�{��u=8 �����	�i�hh���}���H��_U3m�WǍ.����2���߼�tP�n�05(b�mI��_������xC��n8_��ˈ��|�`�V��-P��d�y�I3�K�HWUU�#�Ƴ�n�U��9qHO��ћ{�1gA�
�H��h�J�:�|x�V$�]�E�|3�&�3���-��`�
I����^Iw�<�b�*����1s1g0iK����)��k�+����":(��ʺ�{���DV�������,�$�������6�(ߋ���7�V��zVf�� &v�6� 밅[&0�Nk�/���c�v_U��)�\u�(N�|3uR�_�|��FT$w:�l�6��8�����#�=.B��7u�4�Q3?S�F'n�r& �?O� ̨w{�6�r]Տ�v�k��%���6:iҳ�/#.;B�K'��������.���T�L;���+niUM����g���"�޵<G9:Ɔ�I����j\�a�"���9�(���1��f���y��Bx�庖�Am��R�.���ݔ�a�37[��i6�ӊ`�6H����2�L+���E����y��ۦS�3��1'��K��)X����|�v��5hXEwn�$���ZǪp�%^J��$ �N[ȥo�I��V��}L���P��	?��j�O��s�?��N��=��������*���+�lb��I����B�/��a?|63����Q��:�M,���q(ǟoc�]�q��^V�nz��B���Ӿ�k��p�5�1���#3�N(������<4����k0�Aa}���G�O���_��ȁ��[���ҒhӒv����`C��N@�ْ�3�8t ��ջ��C�y�E��$V��{O��n��z�ׄ�<$5�B�`����őy׷&W�o��\b��e�k�̼���s�9GZDESMٲ������S�[1 ����2ZK+k�8Ľ�$��3�O��yD�+kx�����:���1��i�\}����483���]�E�w�[ -�e��q?�3��$w��ŸE�=���>���[Qâ��%  xȏqN0�o"���H~Hf�x��;��5S9���$0���ʱS1�.">��o�g�4w�>������k�/7 �4�L��5]��9<��Z����C��B�=��Y$/�Ab��ݜ,4���Kf��?7�#.��-�I��=�U��|�+�5j~~�؅$I��l8{����QɈ�ly���d��+|^��ru�"K��#ml�+g�?G�����ʄ�߿�E����# �p> h�?�U��pm��U��&�'���3�ٞ+�㛾ԍ���t�/68)� �X���1��N�Y��0�o���HͤҫZ8 �!�F|L�����߸&������Ja����&�x"קf��ٚ1].����	쬹]��9�,c��.��9��ՙK�?��7�[K;���w�=kY_$�ޞ`�z�_��C�5�4^i`�Q�Ja�f��`�cf2f ��e	d1���Θ��a;`�U_��Ȥ��y#��"��RM�u�����ݰ�L��
��0>�qE�]Խ�X$(]�m%���R�]"wXc�H�D�ͼ�F�ٙ��*ծ���v"����ZHP\�GGF8w=\�u7]�6�j3&8�͖4]笀�႙*�=1sS�.X�9��(F��V.�=H�i���]榋LDӶ->.��bI9]��x�'���u&��1HH�����<=�t0A�o%�j]#[���hm9H�;�촚m�lh�A77�*p�[��~\�a㡋<�r�:Z0O,I�����}?��S���$��p�y�|h��UU��97+��������� .��5����H��^=��h
� ����j�������1 t�J�d��G_���8O����n�}��Cb���l���d����z���nx8&����b����y�t�}����{�{�EӶ^���b�����Z�I:ͳ�� �,�䇊�۴��8#��,����7A��nש��Q؜�͂ށbus�|9!4��\x�ý�bqW� �039�)�Ɉ�X�#���iF�������^6�Y7�K��Gk���|^Ams,��Dv�Z����t��ó3�c�z[E�Y`knA��/���or�<����T�yq�i����|2���`5^]#�T#�k ��z��/��=��P��Ah}@�du��K&%-�JH����r��VG}�ܣ��7 i���p<6�O�GYY0��b(���Q�R۽+���)�X�(�
?W�XK�������34!�a1Y�>�G{�th��$��?}Э;Q�k(����4���t�=��q��̳Ҙ�cL�5����!Vmk�yst}ai�2�w��֠�!��|G���B1�+���/]��<Q&o�S�s7���|Aa^mA����|6}���md qt�ef�wd��i;겉l�Eӿ�qY&���!e3Lz���J_	C	��wlaM_�ܹ~6��`=z��_y\�`3�[t)�T��M~��"��:����!w�o��j[�z���=^mvV���>>�c��_nX\]y���������y�(�h&m׬.����g����:c���G3p~:�CLsk��ի��������]�u��R��FR��w.�X{6��74g�* ��פ����Վ���R��0�3��{��<�au2F�3�`G�􅃒���(6[�Y�m������ڍ#z�Ӹʽy������D
M MY���#t;� ��D���임���r�<���3KZa��ڻI���Ƕ���J���,�sI��U!_��ܕ�h�p����k���}�o%�Pc�$��<�4��rxE��f��Y��単�W���[�R�/��Q�;�GE��&����w�����?��	x�u�IM��gXD�7	�g��ZF;6���7��ۖ2��������b[yT��H��@M=��N=�mEt���&��<��c���ϯF�fJD�\�-��f	�v©��$qV�	���n?9����V:�)^k`��(lnN�"��,k}h�w[����������7 �.`@t��q�dN3��;�Ɉ�h�a��j�{��j��2�O�:g8���;MpS�B,��.����z��M�� �.%�P5��ƑA#����=%ñ��n���׻	mݾd��ρ^��9L��@�6���Ok�U0�Jo��N��#��L����+ߠ3��^Z¢�"X�F��iiR��q*;#v����$�H�&0����Xt[� �o�%[0i;����O�<�l]��v+��t� Y����,�>$�՟%!ҁ~"qE+Ǝ#�R�y+d՛[���o4���0��.@�X�E5:q�L���ը�}���yؕ�w`Wt ��,V��q?�9��ll��N�/)T�� �������������p|�����$�<��ۋ;�2ccb�=�.�.�b�T
J!�<7����$�������
�4�߻���5�e��h�Εh��n=Zdi2����xME���|�h�_̧4�Y�5��\p[��촩�����d�q���ʧ��V˧;��h�ڼs���(�������E�+ѥ�_�U{J18�91TY��3���\&�{䦱V�Ҭ/ﰙ��1Lhy{�[�<}f�0C�����f��ݦ�G��:	9u,�w�����(�w';���H��ר(����٬�ی*`��ń��BLOa�}���m*��(�Zy�W��,t�F�!?��mK�;9�{;��;Ok��������2�+(@}�`�p��?�E�4�����)���.��y;O\���D��+��~]p9:|k �a�C����5�"���n+�G�����5���F��uq��f��Ԓ-�4��-ߟ���������%]���p�a>cb"��N%����Q����%�,
h��"h�OCi���q�v��e�4%�h�`^w �oZ!�R;c�cfBN'.�}�֢P��=�A�t���ɋ�7��VU"ژ�@�D�lñQ�e�B�v&
�'B��.u�=��{!�X�|$���BAq���~����{�]�U��-�UC���va���?��j�L
�T�O>����&�@��� R��5'{[[E!�d�N͓�v gc+ȡ
�4�?��̡AE���ԗo���䒛��Onk���,�1�y��Rd,H�o9(��~Z��L	��#����V&B�w^��X��p���m5x.$�!)B�)��K��z�~�9��P �އ{k�"\�	�]�`)�ؽgW�˷��?=@�2�d�v�Ӡ�%��po��C1�ţ>��T�"��I_R�G�7�8X�~��Gůq�s�r��!�p��ĭl�;��� �]���a�ϒtB*���%ߎ�y?��my�#8)�����M�i	Ha��*�t�֤Y�3�_Ya�ZW���opUM��DI�m�l���8�}�6#��8d'ɩմc!�S`��얚��U�x����W᠓��6�E�T�o�ռ���늉����p3�jF4sC��ǆK�2q��֎�]��$X�����aIn����o���5�u���=)��?@����&B?W�������O�r��''-J�;� ��-!���퉍n����Q(����$�~Oi���0,��us<^�?ՐU��\��;�����;XbBmcA��F����"�
�o=���_���S��y���f�"�]";�n�k��<ob_i��\�"ݲ��ɦ�:�����b,a⭕�e<�&ǒ Ц����ڟ�&�Gf����BX�@�M��4�Lvh������[E�!Ͳ���nwn�9 ��-���J�b�r���,}[3��������9p�-)P�����X����Զ~���1�f�YSwC���_@�	���~�Y�b�m�3𑹻O��C�"��a�\H$Zo��g��y!��4jy�_��җY�	�=��ip&<ICF���i�֛ 7����~l#������V}$CU�_=�ͻ���j� �"J��B j��n�x���._x�@w�Z�	y/���v�XZ,��o�p�u�P��Wf�2f�%RRb�l�ʏ��(�����n��Cx�f���v�'�&TKR,M�d��*���tTU��v�g��]����ȤG�ͬK����%��w���I˂�2��6_ߧ��V����V�J�=MS�q�o�o���# �[����_	-m&�}𭊖���%"�q�F�U\A�4.�w�	X�_Înoή��q��)+���s�Q�(�b������q
��\|��g'��lφa�����JOu���]�#��3�{Z�E�Y)ѥ�CJ'���*��k�^�ZH�
e��"���}�q^G����E ���AZ�+�NՂ��!��m�X�$��:� �������$4鑵u���E���2����~U���un.�"D�%��WyD���w^e�0t����;�H?���zN�����y�]<���z�q)i��,�~R *�l������.��0G۶6��&����9��H*�M������]��]���)�6��M���{�LHd��`3�o���P޽�P%O������x~���������;�ݓ
>�j�ϸ��>D�Eb��
��zL����x�6��٩��=�bǩ�s��;�ȉ�@^$8�LҜu��$%���$�	,���J����!��$�]M�T��0��7��4�2����!ҿ����!um\*��+�5���;��7]&�G�r'�Ru�^$UF`ە��߇���M.�x������]�6A��n>��/�b�zZmvv~�f���+v~4Z�sm�Vc�U��XlE���>�yv����Ȭ[;��:F�I�jiGc��4s���3�b!EYj�͖��	�sߙ�X�f��15SF��Ci��Bd��5�C��N�UГ�{�_@�p*d2�m�����<.�z<����Կ�w�W��fY@Rdz��b�J5��C��^�f�7{���	h#�n�WIJ��@���ú*�w����x�u{�v����������z���^[+�ؼ�wok���C��⌾]��NG*�T���������@`��rmJ/&}^�ƀ\̬��bՓ�b�3�����YIj�2��F�:�^G���9��:��j&����J���{s?cD�P����@�ҹ ��O[E���������z��t��c�=RRo�8B�a�
Gz�ܷ���eJQ��U{��e4���:t�w��{�`��u�<7^������J��f��rm�iU��{��2}Al�����Z���2N�H`m���p6;�}[�t��k5�t0���[c�	,[�F����� �]=��67?]��yh�[��'q-�\D�j�;�b]�NOUXqL��
4R�˭�f������:�KE����J(Pb�KS��=oQnl�>��K(�RJ���=�U�Sm�����xI��ڮ�)�,������K����Lj��-�C�c����b�(I�Gݻ�M�r�w�mt���K]�9x��-w�Y^{�j��G�,W	=&'M�ws-�H��b�N�u��#SM�#Gkzp��3�"��oSqoI�$�Jktx�q�pr�sNDI����Ie�:#D~n[�}A���~EZ~R]���j��^�q�9j�_t����h6� \���I���%��YUy�8�P��u��w]�0����@����P1g��Y�kE�ƛ�"���86��?�ΐ�k�y>�͘�Su���gד��Xҵ���)�����鑓�P`��A������Z͜��Iٺ#�u��I*��w[��P��
*�3$�U'l!&\�9��q5N��q��f����*&E=a�Ȧ��z�L��`�Sa~�N	�Y2��9S�2VnO:c���0eC�Ev���3m��m� �"���,0bۙ��O�s5"7��/E���P�|d1V�wG���9-��][$?���k�aˇ�v]��=n���0�QY���K\��d .���F�{�9��&f��Zj���FSg�:�n���̆#M����Gl�Ā�!�j��[��ԡ":?G��wPlo����P�\ZH�VvX��X��\�w|Щ�o1lч=)�r�ϝ93�ɻWIl�/O��j��J������ �Ɩ�R/��jF����uf�` ��Z��,qG>�qaћS���txԕ/٢��56�~���&&[J�7�cՓ�0�WbZ����k���V�!B�?����$�t�[,�*�2�OVW�箩[
G/!�H�h�����U8�@FR��&:g���J`�&Bg�x#��9���G@�����0���ȨY�5��yj]R���}ʯ�m��R���s�_��7y�N�@0���kFl��n�d�e�v���Gٳ��z��{��=��R@�����rp���7!#�����Z��i+�`.+r[7/d�t�{҂���Z�7E@��	n\���x"p{k\c<m���-�������y�G����'������	� i�Dlǌ�ܹʙ)R��0�
e���ϔ�ې���k�3����%5��4Wi�U�H�]c{z���
"D/w��JX�2۸v�㙞c��ϫX@��p7\t[���@��0�����ė9��e��`�z��eZ'��NT�/v��Y��Ab%�&uJ����q��+5���]�<�`�?Q�CQ�|�ˊO޴��������-�Dc�ܐ��)M�;��<�*����>�r��^$�˳�X5@�j��IZ�A]Bv���[dB�)�Fu�s�kO�`�q��֬HnA��N����H7,��b�#���� ���6�Ȧ��?j<U\A k1E��.f����J�i���%�2��pB����'�L�����Z�ӿ�^,�Ws�X�g�ln9	J�w,���0F��h�1f�.v��eQ���%��ݑH7�&�f_�1�����VX�A׫��ô۵u�1-�-��DR�W3�yo)P]��C����o�_NYo��U+f�����J(�$�* *�,�����4�%��R@�[����4[3��l���{�ڪ��/I�?���}�H`x[�L
�L{sR+_N�"i;�7�jrLz���u��ϸ�j��I;�S�p��~o,�3�<u����tֆ���{T���o�X�{G��+�*A�9�Ñ���F)�
Y��@!=SG.�Pm<_�;�����d�wC^а!8q4m}"����fQ��ah�&�P��o�T,G���⣡�a���P�g�o����!�u�7���U�wԑ
����Lk�i�N�l#�H� ���Mn���i2*�g���gJ������HE��fc�V�s<R}����s�s��ֵY��� ŗ����#�^�� �b���0�Ĳ�:%�'NFߴrS��m8}Ȑak����
�:��r/>���UH �"����[������g��>���A�<�z���z�p�'����̖�1b�����m` �>�t���c��"pOl�cY���,~r_�O��Iw/G'�z���yK�5��:�)�=Fc�!Qak7b��*�X=��X��Xa8h/?	�R��#F=ǎ�쉟J��h���9�,�
��m���踻?+ʺ}�y�ﵷ���Z�b�=��4'��:�z�<��׀K^U鮢���?JIOg����:�U�J� �7�d�/ݦ%{���h�[S�?��_BNڠ��(%A����".a�[DL���).�h���l�1�,W�<��J���|�ؘ�>Fa]�y�+J����F��&)��K«���I�0��+&-a�b�K��n���>���ޜ|�ש�p�Gl.��d��;��besW:�1t�H�Ek�nZ�d@b���/�%vp��,�P�Q���,h�&9�b/�HV�#S2�7@�v�������~0^Ե?�CX�c��<�_ټR�!1~=y��I��b���(��eo�z*4���G�����߿�?~�B��G?�S�8>���#��YV��/U��s��zOx�?���ּy����w�Z>=�}P�KC�t��,%����l0����i�"�-1��ε�D�-�ϒ�o蠨��"�81�O+�gkj�����P��Y�!�!�{_�ڰ~��$�b������Ţ��]�m�tV>�BA�g"� �'n=ȿ!)�%e?!Qj��U2�y*jO�Z�(K�������C1
GIt,�N����#�kh/Ć�Ӽ�N@&���o�<R��{%�*��򤉱�Ur�Fk�|���4�6Xyh�`������[��P@��C�$��h��#t�H��m$��l4ArJ���ڐ����\]c!����'&����{���^	OV�T(O���G�������Ě�I��~��ç�%_���gT�i���+iQG�ҋ!�J���[^�Q�T�G�c���4�QI�9��9����ol_}��0��ъ���#'x�IaRQ��kv&��x@3%>ց	u��x���8�����LO��!|w�m�}�"O�z�D�r6!÷..�I�����xQ���5v�>��] �}}��ιOW����=/;���/�_R�W�L͇k�}S͇G��aj�5����ħ��4A�uw���m
��1`9H�JP4�b`�ذ�X�aFq<oHU���2��.W�s�C����1��W�ֶ*�ӌ+�V�Y#���Wc5�����v��#jZ}�D��jۤ�ul4���W�n��z,����B�壙\z�pW�l�	��H���z`�^}�~o��^�?7��}�>@��~����A{\��l�dVq�F�+;7 �D0ASp����+���S-���R��n�.K�G��g�=�`�st�q�rZs�l5mQ3����R���6}� �j=3v��_Ӏ�T�)<sUX���7�>�L_��]k�Ѧ�%D�|�0N�Uo�7h�S\�;5�9����uq.~ǧ�I����#3�Eܾ���J�E��<��L����,͜��He���j*rvÀ����؂���%�x JG=���O����K����F�DaS���X[��4q�0ߠ��օ�����+���F]���_�W�L�\�F�%�<��嚽�G�uܸ��^BR"WM%�%n_^&��V���̄9�_�z�\t=1�m7n~]/@�<3o�U�� �`s�}��nn�N�>�A��P����?�XOf���V��G�=����n�eQ(�z�vG|z���0� �����zA���$˶��輸��o��i��"�c|��gԔ��:�%~
D��R�g�а�lcW \:�<���@�M5�yyM_#��P�����#�Ņ��� ,j�E��eǙ���B3kD2����8����u�;�@Ʀ���m=sB�MI98�_��d讉G�w-�*!��,Ho�ZG/*��ي8+���w{�̿?�;*���w��"qw%��%"?��m|`k�>���l�$`�x���-�Ͱ���{e�����hx8��٭�~�'���#c���f����
�v�5�h7���F��֯/D�zZj����!���x�Z/����[��2_>c:�hH���n4�P��!S��|a���Y�\�{����������"D��+���f�3\D`ǯ�o9�8Pɍ.cU 6��_��D�����g����Mu�7��d�%�,1�-g$��Hm*1��^�C���G����o����P=߯?��?�I����x�P�P�s���B�����p�~��Y?z"�Q���.�3�j�ۊ�UH2���?�G�M�*��2v/P�?�*l�.o
��uwx֐����|�w�w�6��p}��"����b_� ��_cK���am�d�G��R]wSg�[�������N�ݣV�ŸJ1��W+�i1������QR_;��W��ru��.��_,mz�O�v�+^�g�����M�Om�KO��n'�>+����Шi?�:�8P��4���u�{K����%M���V�yӱ0eIv�lMv0�n}\�*��C��)ה�:I�g�
Nm�'t��ˉYn����^��H�[ V�*��-����&.Q��nB�#�u���7��؝&cy@;�E����:s%6&���sw'�i^uN�d�陿�S����x�6�����|ơ'"��T�w� ����׀x0�k��0��[
,�{� �&���.�;.��>��=I�C`st)HЬ��c����";���.,,ٷr{/�j�!��D��W(��`9���V��FW+&I����V�w�Z�O�ONGx����]E��E�_�c#�E���\3���Vר2A[/�����ε~|}B�D�>v��P�*�j��2x�3k�Ø,�7�9����z���M��{H��a���/5ZcjQ���'ޔ�#T��J�cun���w�(��h-��
�u�;o�,ٜ�qP�Τƫ8n-�.T�;d��%$o�x) �"��/>w1̸'���n��9�+v�n�>��\�"WY�P�rD���m�R�.f3!�'�3/�ۋ_�\'��c k��8&{�t{z<9<<����P��r�ǃ���$�<*�[^��Tt#��0oQ�bd+>ط�^n�����ݷY�o�����e>\i�&)�k�m�\%��׏/ϋգ����in>�`YmN{�휝LN���zޗ0=��ʦ(��l�b�8��IdEƟ�j9~�[�(G������i5v+��'-ip��}��A�v3|e��4�=�_����}�E9�O�{PR��.����Mw��'�j2���oLӲBc�
�Vƶٍ�]�+h�ͥ�1�;[�$�[^<�k����M
�1(���44����-�1껵d��Ο��M�ݗ�'W����)��֜} �C�ệK��-dj��O��퇩*6�9_�??o:����R���T�ӕ����^y�{nX�2���9��YA�n#D g�ޮ���ɴ�i�1�(�o��~���T��c%�u h�H���Ϛ��4�e����]<�lR���������Q����|3W
x�7K�e#�Q��B�w΍R�xo�M��Yil�[���E�q�����l^N2�h�g���}�*A2<�a]1_���.�P�ҲX�T���Q�E2���*OC��Py�����������5W̲-�%V�S�1#�9�tN����-�PT�F�F�5��O��T*��JΆ9
b��0Z�A~��v�k@�9�`e��Y֦��:�	;rAaH��S�(ن��Y��z�|"2������i1�͞�� V:�8�ȟZW�9{�T�Ҥ�l��x��2o�rG��O ���28�i�k���-dKe�A�8�Z��3�/s�c�s�����!�	�p������	x�4�uj��s�"^��o��°W]x�7�BQVOe�k�8��"�I��%:�: ��__`O�w6NK+��5��}k-4Qgv��ֱ�#��%�ߟ��v��5��ν����-�m��(�h�X=��;�1tSQ��<��yGx/�:.6��2���������g��X�Ȍ#V�u�uV��i�B�}��IN���F%�ۥ��'k�jr{C�7]���}� N��^Tc�s^<ZnID! ޶��$�3[��=1�۟��Hxa wGDs����o�y9�qr�#66�L^_������{��)�������Է5����ح�`��u)���=O���r.eW���,rkn�%K���&B����j���;�������DG��ƊRO���x��2��J�����\��:b�Ŷ� �<`v��_3ŷ�o�������*���¡�M��;�_�̀G��G�}��oW<���L[[.�H�Q�iS��q������n��a̜݊E'�0���p6J�A]
���ӈ��Uv�������U�s�I��o3������,^f��v�G�����Qcz ==X2�cH�r������$��	b��I�r���R�=���qEX�G<��+)� [{+r�a5����n)-$���!f�=���/�3�+:�[��1Xbv���S"���^��z�������h%�)Cf޻v�M)�Em�\7��Q�N��j������yժ;�ft���,Qv���t��������	�Ы�H6Z|���up��"���L���ţ����o��z��F*�n��5����̧6��{�V���[�bMA���Y�	e&�4��,E�7�1�� ˉ=j�DD�.��Vӱ��>��i)������� r^�G4J����k˥l���zj��|�'ڑ����k��|�?��
'��g���f�5�ߚ�w��x����yFCãQ��P�G���l�x��o���;�UHUe����-M$T��Vm�����D��.T			�u�SA��TJ1�܎�"�hoE��V/���|N���8�+̱�٬|JR�����9L2�C%���3�B��5E̯ɛ��a����x_��p|�>���t����ܨC�(�O��e�=B*�b^�Q����tSat���r�Ÿ'2?7�ς�E����b�`�k�!���2�@}�`��VE4�n�����O�Sb0E������v�_J���1��u�{���\m���A�jSY&�ʻ����u�����SGϭ�k2
�������(S�U��8~�M�ѹ|�#�э�,��9F�U��\d��Y��{����v�	�z3�ٲ }�M��Z�cϫ��~�����X��maݤ,���Kr��y�r˞�:-�#`�<:~�gY8,�\<8j����B�����7yo�����WHm�{��M��ئ�IK��{F��	���VܐA��o��������Ҫ����*G���0����Y��"�k7\	��q��p�1�4��7E�9uI��L���M����R�5�7k�����u	z�F~�ڷ ���ͳ��r˱*7��/���G8XT��7��������(�Bu��+M��e��0��o�yN?-{�Q��Qh՟�����fzs���,/�eU�J��*�ϭ~JAaԭ��1���;�	s��a>4�h���Y�O���d�}��*��I���� {{����J<���� E�u7���o�@rƇ+̛Sޟ,����Д5T�y�3|�j>�NF�8����I����\�b�R�ݷ�-�+�&���/om�sBC����a�m|������mO�t��'��l:��߮V�����O]�[/�PE)ջʎ����P!M�m09b(XooV�+)*
K�̔��T�T��;̀��m4B}�[�ڜޣ���g��]44뵋�x´?Ԑ"���(><��jNO�Q���I�����������kG!|,�+fB�g"��uM�k�ج��s��j6��ՎP,;��;��`�v!��`�P��~���l�n����p��X̊�a���'x�z���1���xo��\�Q�8�Z'�kK}߀D�˹��l�q�:i��#4?�Rf��O-����U��1\���1o��|kW��� ݵ?���d�OXρ��M�83E�D��^W���N��?rA=Gy��χ}z��Z����_k�x��	N635�{��HOE�nǞƯI�������������-�>]ȧ��.Ag�!��>\�FX�(󩕱�` ;�����?�?���[���>pF����O���k��HNRse)[:ĩ���S�=��	:�v��vF�?&�\0F�e���P�=Y"]��!(��D���˨SV3��ڿl~7�������*!b'�!�XߎWkM�b�説fEAńT�;�4����(��4r��]�7҅�����pݚ��K����p��SZdZ�D��o$9����9l����q�����YX���(O�3���;�i/�'!֪�nr)]��6��cw��K����]-���=���d�ef��21�~���TW2�>�:�
�5��m��c���}	5܃��>��+y{ㄥ�������v^wLͮ�wh��w�A��2sp�E�`w�&��^g�N�3�?U4}��L��=Q(�F2��kq!ŅOd�1�i�3j�^�n�·$x�1��i��`��՚� �F�ǰ����2z�-.���(A� ���/�X�pڟa�
�Z^Q��a�%jh�) �H���rcB8W�^�����o��]�v��$�ܑś�5��AJ�&���|0��IE��Cg 
<��<�(��I�q"�!�D���_�O������f!��r��Lr$h��}��>��X����+�]LX޶�_O�gj�v�r�9�sb��?��ku�0p.=y�<V�͹^���v&�	ٓ)�#�Y�S���{��ɝ>ko6乹ّ�B�0􃥴a�y蜄�U�T��f�\u=&J�e����r?\��e���8̧R&�݉�� �Z9��������m $�6�(�])��2^�o��o���F7��-��u�2�^Վ��KɆh�,� G@����>�֜H��j�йUm�8�c� �|���k�#=#�������m#Ҷmk|���W���)<����t>3��_��ĉS�����j4h���ϔ)��/SZZ���g�ӫ7�Oc�������w�RZiG1'r�Mmرy#�>[Ī�Kؽ�g��:�U�ճ3�D|�hߊ�߬���-|�:�Ĺ3'����v����_O�{�Ze��&�ٲi=OO{�˿$77��w�����}�^YC6dJ8DFj�<G�Y�z-=������{_
�<��3��ۇݻRVZ�*��)n��\F��Uede�PVd��B�����_�t�<��K�U��j����S!"�a�`��s]���t�4W	�G�d�.��Q6���O�k1��dċcžD�Ao�j�+R��ԩ߈����S�>��ߎJg��ś�v�Y�<��~��D#�=��[�b��ݴoۖ���;�>`�M4i׏���QP^��l���H��^%k���� E�&+^�}���F5j����l�_���zvN＜��=����׍�_rn �����9s&�ӥ_l�y�J�6�;P/;aäQ��*�"�i��k��=��Z����b��_�&j���6���_�w�H�?_,��^��1c�#�=6��x3���={����F�:�����$�gss�Qh�M>��4���{�mdg&���CUe%i�i��.�-VJ�����/��I�<��+6�T�(:�*oC���a�4<e��߹��ͦwSX�@mN�LxQ j�@(�w�r�>}��?�
��Gjz�$b�3�7�ό�p����b"59��d+�M� ES�-[Ƶ�b��s�̫�лv��W^���S���� ';K����ʫra�촧9{�
�l�Z�nj�#�Ƕ��9�U�%$�����>E7a�r�8.�Siw���F�Fu�>���"�4�3��#j�
���L��NN=D�F��ؾ�4�����_/�۟��g�^Ǝ�MfZ�lŻo�%Y��Y,\��)?Ğ}X��|�A?�N� D�}����Fj�J�Y���Z��9�����w�A�Q�F5��˥�N$��i�3�j���?j���6>	v��K�p����|Q���k���^CH�Feb� u��hU��Ū��0'i��o���~Y"�D��-	��'��痣|���k|���ؗ�M�1u�x���Y��\PH����VV�^͵�J>�j5C�=�>!?aY�}�m6t�<�PP���������z�s_������$��衮���e��q�k䮺��[���Ǹ���gn ���^��WRTt��¬�[N�x�y��wl�jR'���}�|��\��]�۰�ˣgη8��b ��J�	�֠yK����)�p}(B�.�8{t7aO%�^
�8�.�&�JNreU�T����6Cј�z�Y���Ɋ��ɟe��H�j�z\N��q
��h��p� �~K��Bx&��m#Pu��//=q?��BiZ�W����#F�*>�F���3h0��<:y<��ë3^�Å����&��L&#� ܭk*nܞ���>p�]�mL��y�Ժ(�nݺ�=aC��m~~�p�N��|]��K�ֻ��x�3�@��'�ãS&�h�<~�	�����W������R�^�zQ�	Q�t�7@�֭���E\+(f���MqTV8eZ0����IzZ"-Z��/�L������-,��kv��۶0|�`�.���Y\�\���ןM�7SZ^��%�s��C�;��{Z�kp��9�n;-Z7�����������Q�|�t�[6㻍�	�}2Z*��8k�$�"¤D�@' Y|�H]���ZU���R��0G�g�{��_��e���P拂|̪V�\�(��?����E�H鉶G��B|z�nFDk�^�h2I���-ӣCK>��6�F�'}TJ�
@x6���t�x�u�L��ښ��U��2�Æ*�E�SK@�K�&լ�8���M��Ͻ?s�G����t��3�|�M�z��l]���=���ÓG�������77 ��wO��+���5���ް�bic\"搃&5s�uk���[��_��\���Ǜ-�j���u�^�����*�Bf�EK��0�->*
����i\=��We�$B	&�� �P!�������JI�v�������=r�\8�Z���:=O@�Z�	��*#����%�ra�J���ʂ�4�3���_�&'T�l�b�f.�W�
�	h�����e5�;K�����ڳ+~0�Ͽ���'�����رY�n��'U7aѲ����1|0?��)�d��%5�ϝ;'{��F3�=�G�C���CbR<�׮�d�G�>$%R=a���^z����瓏>d�(s�	VW�������+����\�VJX��R0��2��GO����9y�\�u�0q��a���ٱc];wc߾2����\)�Ξ}{�N��n�
q�;v��YPP@��&ebE_�&MX�f�L�6��}{�.�FFjə����-^J��:�W�>�=��%e\8{�S�K�wq/T�,$��B贆(��ty�K���u��iv!���qȱ�5�Puu�}��6�J��V�EA��M��á�T��l"�/ljU�Oz��D���Z*�AN]* .55UXfO�%�ٰb	��Ge��y���T�==���"	I|��j��Kz^}�B�^��u<��*�>I$jū���̴x��uU�)q��hd߾��������yמ�5�u�۶}��
�{����]���<pc�����@���=�>��g�\�ӹ����Bn��L4��+�_=���;7]\;�v��z��7_�mǌ��5�Z\��!�2�*R7<@��;r��%ij5�p������h݄3�l�U�<:�k��-����>�ٳ�d�p�2��݄˧�� �Fy=E\��+���ڵ�	�5d�gIv���HKL������6���,�	|��"�>z�U��<�Qg���a��M\+���o�Ƣ/P���ˆ����5��ڶ9i�\�x���6QG[�D���&Q^^���[��K $z�5t�ҁ�8+Uv�����}�&mڴ��p�r�
^��d0����f����o��!E֭k��ŠSa�����s���h���n�B^~=|D�xy�>�qF��3�ͭAE��_�'!)��'O��#z��^�����&$�S�.�=Q���J�y!
SW��f�I�I�]v;NG%V��aĐ�����Y��d��<��[��8�m枻'R37���ߒ�.�-gZ=ހ�,�l�	� �1"�Ѻ���^�.�[�q8$,K�G��>�P�T��
�y5�*�>�K�8�' TD�¦7�դ�ǎO�$����I̮E�=�����T�
���a�{1nX�|4�xM�p�EJ��S7�{p���k֒�m��c�8̩��n�\��}n�U%r��B+NQG��Z�~��I���s�S���_��yiu�˛�:jh���O�>��¥s������]�.Resa���0f�S�����q� ����[����]/�������F�*G�u���@��42��g���6�[�`ZB�i��+춬+���_.����˽����%2�Tk-8\^�-��WVҼ�Mx�!��_�g��j�^E�JM˼L.��M�ӵcΝ;M ����i�N,���g砊��D����J��z���"E�����������A�f����^aCR���p5�U]�rѽC{t�
�-_D���گ��JMie�l��u+7m���Q��Q|x�KI3���H�(�ӡ ׋�0X��E-7>�,���n/N��ΌJ�}�Z�f��n -�UU�Q-"��E�X\\,���^Ѻ$��D�X���D-T�[m���Q'�#Z���T9�ęM2�$�  c����X�b�:�J��d����AFv6����$�J+�9�Ig���,��(\+����M�8�f'@6>!���2y�ɂ��F�;j\�2�]���9L�0�z5��}֤Zuh�<4��m�FeY	�f�O��s"�"���B�O�0��qM��T�Qc��	�3�	�d_�XP�"�Fڊ��5u���<��<��:���V3ee�v�]��ՊVF�҅-�G�F���X	�0��BmM���lA)�U�݅5p���iN�UOŵ˄�v
���_�nm��8u�<��v��~��oA���O�`w�P�
f��p�-��������G%�7"��9^�q���඘�F�ޫ����$^��d
չ��b��Q�S��~���!S��1d�>3����67 ��vG�����[_o/��p����6B�J�A�D���Bj��"&׈$��VS\RA �P\i�җA��'�Je !���P�A}�ť(�8��H��0(aRU�Y��]:@�Q�=�~��^-[ݾ�j5ks?_J�Q�d7��U�F"�H2�w^���I�In�l�6�q���� ?���}nE�$�l�~�O�v��آ9Mr3X�Ϋԭ����%���
|/,��'�˳�3���$fV#ͤ�FZ
�F�!�Q�h�_��l�P˫^�x�Y���<u�/ʼ�%Pc� *E� ��-LN�Z��(��FD�)Z�D,���o��V)	�q.2 ~q?���V Y@���q��e�*�!�D�)t�x��Dj�,�P��9�Ӡ�t�Ɩ��!�����T�L"(���3dff�(�p�[�&v6����D4��FNz"��BB�JFD�z)$';��J+�<S\�.�Ҋ*y�׭�������%T��`2���zQ�d|{\��d�˲� �UUUI}��Tjծ!e��"9YH�8��Qv��Me�CT�q;�r�E�\δoך!CȌ��� �������?�N���@�e�崓�� �5=��:�c��%�t)��	Tz#TZ�Z%�A	�/�N�Q&k�S&�E�:����G�N]�/)&�n��?Ŝ�Ftx�E[��V<X�o3��>��g.j!��0�A:���x�,%��(�x�!|A��Cx�
�E�1��<tט�;`�_`J�q��bn �_�Ѹ}���ۮ9o��L"AB;���@�~|.fa�)@-�O�� ��p��p��z�	�V�L�b5Q^i��s�Ҏ�d�Z�l�Ue(�6�e$Qr� �;�$'+��k��Ġ5k�1x�����ڂC�Gc��z�&H��Ǳ�[�v�
�}�.�P�ƍ�
��kiX�)�l9~���M�(��Y���KO�����i�)ڷlIvz:��Q��9.��>��C�P�^=����&1�w/��:-6[%���H骑J`Մ�5�����g$�J��5	�dE$/ ������K���t�e��&�.R�⍤R�4�Hˋ�R���'��Kؗ
@�,n��7 �l�"�uy���^7o�~���1>�'HRb^���ߏY�P^r��G���2�IN��B �f߁�|��v��D��J�~bRnG���Czqϝ�	z*Q+vU��A]�>�'D&蒤%l �c�{�P^VƂ��Q#'�ʲb~a<h/5�%Q�z&f��Z+;��_�Y��L���I�T�p��ت\���ә��B���%�FCYy�|�-Vn�Ո�J�^�9Lv��(eg�F��Q)�*��
5��s�8��%ݡ�'lH�+�8�,f-��^xm����F0��^\<{��]��j�Z>��3�������D�JH-�XK$(�o���_�_�/���D��S	�d5Z4�#b�"���)a颇V�/����t�ӛ4T,!/��c��[�����x�����/��d[�c�]ѡ�	{<(��`�ۍ�����eGo6��5Rg]�5`Pkqڝ����Tku��&��d��\�3C�OW���L=x6�.��S(8w �N�Ly�����gN��ǝ�HʬN�7�:1G�,'+=A2�Z�6*��#/7�vZs��X��wnێNcD1�(�Hϫ+��۵jJ����}4�M��r�z�!�=/��_s�r>k
����^�O�g�}�Z��Ԇ���ONZ*A�[���m��Ir� �̴TIhzIwao*��D] �H��~em�I[����R����Z��T�KM����o�n~�z�\<dee���ș3g$����㓀D{��+�����"�E,*�]����&#u7f��-z��7L�=���Cpb/�L��K��Z*+�����h�	T��Z��E�m".����sԪ����QqU؅�8��K$�B����JL	�����~���4�ٳk7߮�@b����Fj�����IO1�񔓚����e�����%M���zY�Z�JX-�f�����rE��7=3=U�siI	qq�v�K�\��rqͪDH�F4��k�m�8���p\5�6&`�����̚0AGj�����O<>�	w���?B��2{�<�,����ǓY����V!5Aa�����񸜄�I�Ө���h�%y�`�BK��8g���J'3gE�V�#�b�B�.����>2��ҿ�Lw��oD��g`���>�}� �    IDATr�j|yD�F���z�Ho�Մ���M؍ޠ��fG�7���Ъ��<>	�n������ ެ%⯤n�\�?E�e\�^N�.]���F��fpI5�q�^�_��dV���ųD�����S!�f=���M� k��d�n;�0	!7珲a�֮[)�V�6k�Y��[,���1�瑔]���M͛R=��WK��y�{�h�����g/�����ڵ����u��=r,M���[��hb�'�L-�%���"j2��٫$�fgdbQ��GQiIT�D�}F�� ���).*���v;e�)D\D��VQ)�.�$& ]ԅE�B�/� /~' ���V�I�_��b�n�^�7^����łBԔ�zj��~���h���8tz����жE]�y�)��A>[4�������V�c*�EF�*���+��bR����g�.^w%h�XQkrq�,:��
qi<��dW�c��[Y��*�j5��R�zMT#ު���@^Ge��K/D9��^d=T�t
���t�*W�c�A������)�F躋L� ���ע�x� �$�A��&$$Ȓ�x���k�p��5̩��3|�����@�ϡ2�&��˚�����r��ZlŅ�~��tm��G�H��9s�%�z.�v�g�$!�!uD.���Z.�P�х�h��ylH%;��.�(�R�Z����JMX��?�F-�|�
.��*e⨁㟺s�Վ����R�x���{���,�z�jB�H�	U-o�ڈZ������
��!1���V����W�dn4X$8	G.u�K�t+���W�6L�0�>�o�~�&\*�g���h۸���[{�h�z�"f��������D�;��*5���+gN�j�S͢��8��ﻗ�+�a0�Re̠���+E�h2HͭE��O��]��l��wf�����^}q�},�fFK"ղj�����3r������Sv�Vo�YQ�I��g��V���ĚG(�ZV6��J�ŋ��iXR��& BHז����������
�ɿ|EF��?��ɓr{��ԌL�Zw8llRRҸv횘��q<n����)�-�".�1u4q����ވJ�q�]|��k\^�J�����ۇ��w��go����кY:>�y�R�8i�"i��Ë�d���ZB�L��Y�D�.�� �Ȓ��|�>�����3e<��L0&s����̮Cy������{ �ʴ��wN��izr$gPDD��L��9G0gE1�a]]Úִ��3���4�����9������z�z���}�y�ٕ��f:�s�p�����6�"�����s��S�DQ����(M����&R�T:�r��� �K��dȐ!J�P[�@sS�P����Қ�Xm�%G�F"�QZT�H�҂w9��TW)ЌG�8]Vex�$��w'�}-#��H�Y�;kQ]#!:��E��3)y������F�!���_�0�P'ɜ�SA<��_\�n��s�"[�٤�e�u��͙d�$���+��>@�a���A�&cC�+_z1ͱ����=���l��O9���Λ���`I���[��{�ܥw������,N�ٸ�%e�i�����XrX2��AL�}jV4�O��m�Pld��#�¦뤻;��h�}˵���Ӭ^��^x��o���N(؅I3�W5�h+]�X<nb�#j�Mgs�*ٴ����M����<�cAj��-ă�$�m`�)H*C�1���]�m��-{M�����瞍�H7R�wFh��{�p��:TkS���_T��bG�9GL��_�'	]�N,%�	�\q��,�M��`˖-��mfs��L	�C߾}ɤ�=V��hO��6I]�]Z��B��� ���:�sL��VT* ������$�H�2G�*pp����c����簉L�Hc^�0n������L����x��'P�KP��S�]z��Mx�b� �e�}�V������%�[�����rani9�X,����D���<��r��8|������y�y7�Q�{3�W!En������Z����H�q�Nd��[��ѴYI(�G/Ns�XJI5�\��HDU蒈&�T"�X�}kz�q9qجx�N�bn���PX��U�:��.aܑ��qU������"���j=��d�D����k�|D�qJ~�VM����=�a��&	k6u�2��%U\lNȥ��awc�2J� ^����ɒy��Wִ���m���n$��'�kX�]~<v'2�?s��K-���w����+���=p�mK���1t^$oGOd�'L܆�"�͌��c�p���������A<�"����j&�%������:��f�?�T����(��o�x�~f;�T"�����O⛯V��LB�#�C@.������p��#�1ge����dJ
<��g�m��֍�,lՒ�<t,�6���X��x�_j�q�ln �T�˞��vPZRA$�!�ż��)��i�0�	z,�{ٲ�g�>�*�SJȂ��բSSVFaA@�A���&S�5��E��d�) m�F�����Ѕ �R�2&6�CI������V�+�jjj��󨖾$�E�q��}>���s��i�0���9/՜��:����2o�[��s_|�^��͆��8hh5����wY�i�*�ib�*�l%��+�e#���uF���e]66r=V�"�%��"RF�!�i?{	{[3��槜yލ,��>���(x������y��ٲ�G���^��
�M4����s�UPf�^�]i�e3v����y�L��R�����l��*Xω����bS��σ�aWպ�Ӊi��.�
�;�W��y2����y���V5m��i��� �Վ�I���p����dg�.;n��G�f����L'p	��Wy����dr�~M����2�E���S^���2=�]W���%�f�I�N���'a��#����3���k��������?�����1qNG(����`&S��*Uz"\�3��L:�N�~C9��E$�EtD c��}~l�"ipn5O,
�;f��By�ν�B�}��L3��y�g�1�p�M�����`�TZ�����IkG�/_͡��9G���'����r��ש�^��U�Z�EU�ƻٶu�~�3�<�$�X����}��uQtw!�x�Pk3�x���J|5��#D��1��JcIg1L[:Ju �$ik�%��a�Qmf��)9T>�ݰP��(�Jz��]�y)�T��0�{
�*6��c�"1�RAoPf�� %�2=���ck���/�n�@��gr\=�t�$+i�M��&E&����˓/`s�1,643ũ�f0"̝>��b�V�c"]'Z֋UW��\͈AN \ Ī��\F�9+��������]���:�$L�|���gs��7Sի����N�;���[n��ֱc�V�>'�D�8����u5����9z:��M��)�/	;�(W�YdL��>_�ekK�v�)��\����QVZ������ҹ'���a#���+�ǂ�e��s�xz�*Dk0�fH�Aê'�%�hW�|�\�d�y��8ٶ ��l~1�`٬�;�*�=�2qy|��$�idt��cGǐU8���0Hf�dE�`8��v�(���p9�$'�6�:q���W6ŝ�pڱ3n������,i�Oq���{�{�M/}Q:��ȡC^S��'C�Mt��f�BJ|a�z�h"KSc�{�~���	���G��
kފn�OY�sS��hY2>��n��VΘ3����p�M�;f6w�xu��Ȋ�H>�����U-~B�9�E�7��.:����g���[o���B�[�F�hee�b=���G������X�j5�?�[�:���2���h6

K1�~�Z��]�Y,�ם�`O�Gpf;�]�!�ZO:�L�&;3lJ&%�����V-ۼ�cg�4y4%c��P@V�z��zf��1���J' ݣM�g3m��*�G�b|��w������=��9�d�ݣ0��%nB&�j�--٬��!�b��5=�5�N&⌓f3���1�p�B�Y͇�I���.�M"х՞°tSp�U�:�E�3�T���x�J8l��V��ɋ��lh�����'�Y�����bsi\r����Ow��U^��͛	E:�H;]��r�8=NE�hk����G���"�ݩ6�mm��	��ٞ�l���B���+N@Ks�-[w�����W�|ڦa�B�*�W��9|E����7�RL{����t�D�o$1��O����腸%d,&v	pF���js�
x�n�pډw�Ԩ�mbW �#P@kG��"2�8EŴ7֫9zqe��H�g&��c��g3XB��(�|�/@&*����U:|�8n��[�����+��3�_���3o���O��w���7��'�f�q�����.����ڢ$�A����]���x�5��]1��z�����w(��!d>�xq�	'��s1�M͐�2n_��>��̛=�%��+�s�H�j�������������;)--e�9
��͐����,W�q	�uI$�
���'��~�׮a�Mw�=d%��G�ۣ�jw!��ЈYR��)�,�Lb�X7�X�+K�H�C�D�פ���ىvK"V�j�
y��=t�b���������ֆ��U,�}�d�.�K�-@�N��ɊP.(葩��$MZ�{��U;�^��9PD�x��+��4��2�H��q�Ӫ�/��3~*���T����2g�xfN�ءn��]�� ����|���J�]Q'Mq�h�3ح.�W�ki��뚝h�Z������ha��*J��*���,$g+㹗>cμk���{�i&����E<��C�p�tB�m4��������]v\'��6��-4r��S�3�kt�	��,V�&�❭ab���ށ�aU�?Q�Bav��MSs;�pC�:(��ֽH ��g�@/�\t�1{{Íi��b�sX�	Hv��/��p��kd�q�KE���qE$�M�8f�0�nb��uz�f��"� (n|�	n�]�n���Zte�[TX�a�H%���gu��[t���hohR��f`�cH9��)�>p��w�������B�}��|^��λW��i����=��1���6�/�A�r�DԼO7�8ܥt��F��������{��ޣ�|�46�e��*�~�av5%z,ał3���̂xO=�$�>�=����aӦ��Ң�a:���h���ıǝ��)9`�HfL���bg�����d[t�_�Y*�c���[��[����,Zr/���pU�J��ߋ5��������y�R]a┹|<M�+�4�#��5�OG�$#�ܶM�˧<ǥB����[U�Z�R��۫R�lv'n�K��1ɢ^\\��[g�ڧCW�/���U
����.�[S�ȆF�o����W�˿�eS �&�.�!�wi�+��dJ�#�L�9��Sx��7qz}d̸2��z�������"�B6�J>c#����?���Ƭ���q�LJJȫt��P��ș膃x,CSC7��W��J/��B��B�V���+�s�����V��D�9�t�T:��1zxo~��{>[�����{H���PG>gꔉ���M0b��z*��P�k �T��֮a��݄;D������95ϖ����}�ۻJ͜���{w-�~بd��U���{����J,*�˼��b�	����T�
?�[���b�CKc>kq��bjYe#R=ql3�)2��l=�?qS�+:�X�Ds;�����EL5v]6m2�ɛ�\v�^�K�ꛔ���립��b�
�ӥTF���>��n\t��s���r�W����ASS��^]�쫯��9�`�D-"SˠeӐ��fԂ�E����j�v5Ö�9.���,}��;w��r�9)�Տ�}ga%	���E8�I�,�+��_U���^��N*��Q.s"���Å��e���L�8�O:N��/��2����+/娣���8���SJ;�����BKs'^r�X�}O�ۃ$4VL�-��ҧ�����f�����<;� �!-^"�-W������ןb�N�UW�i�ŰŤ��3���0@�߫Hh;k�0���SY^��|RA�u�
] [lL�('�/�$af�^f��s{��	�0K�����.ϗ�ľֻ<^���sy��aW2�}3�������2�8��pyt�'����з��q3G`׷�4�e���io�Vnf��6����'��3j���6Eȓ����8����x�HmXl1,Sɴ91k)��e���o"M�)�{�5f�8��ʹ�yh�N�9{�ٗH$���=�i��8b"���n�h�[Ϗ�70�y�"&o���nbf�������W����\]�ۻC��<V���9�Ѓp�zR�:ں���rY+���6[6{�P,BU��\���G�F�VL�[B,o!!�p݊5oǁ���F�������������d�Ø�S�]�B�r{ˋJ#��j�H�)�(Ô�T	��d��\�U�a7Hf������X(��_��[�������%O&k�Y�zlx�a�:l�����+�͗�����\����o~{�
����_���]SE��U�T��R]���ćJ�w&�����M�Ĳ.���x�v^}�\�)'��֭��?d O����c=�3���t�&g��rݍ��d���c&{�x:�4���LVT�[p.No���U�5}�����3~�裴��)�g�^�|��:�p.��Z>��[.��~~���IzW�PS#��M��"�b�aϢ�R$Z��F���"]t��l��3�>�����ۿ�J-r�1s�}�r�8%�E
tٲ���'������P�@���k�Ke-�2J^��*��}a-چfQոH��R�Ku�#}����o���U[^� ����tΰY�J���MЭ�j�������LFGك��0';�CG�Q8���1�d��2�yɛ����e��(Ua���aq�y�)�x��r�p��Q#	�W#���J:��]0�'����J8���k+�Y�p��<�o��8����5�DS�a������x�HJ�<�#!v���G��ݭ|�v=I�Jw2E�j�[���n�鰪�8��IZ[Ȧ#:()qs�ac���6L�sG=1�9�5%>�'PRޛS/����/�R6����D�4�8��4���hX�{8
H��y�@�?y�6�����ID"d���T�ײ��� �y��.!۹�<%D�q��Ie��F�d2N��O2��a�b��Y3�S�n\��2d��3��ѓ�>��]�^�o���?������v�
��x剏?�����/>�#G$�Y�I�2�P%Le����b�wV'�1��=��V~�i��s�Տ2�ٜs�����g0?�w6��IY�� �g3����[�x��֯7��������N��0��޵c'����;w��1a��̜9�ѣ�r��CU�y�X��7>�P������q��~'��{/�R6���5�~�鋯gSP-
0��
�K�B`���E0G�g1�Qb��9���R�8�:� Z궰���T�c�MF��/�6�4����Ś/>#SVR�*�M۶#�n%#33j�/_"?�0�`���Q�T��*my� ��H%�k�.��T�آi�����H�/�+_R�����(.)Ssb���*�l���;�"�H���<`� �N=��?��^����o�8�dS�D��y5+7Xm=<	�Ѱ���b�K�YK��tNm8Z;�q�
05'�\�L��g_x��ʦM����^y Kn^̖-_ѫƥ�w֬�@��:Z��̜>�>5�j����1cƑēYV��P���/�;�!n��x���ۉD�t��I�M�6N���U�5~���}˘4�`e���a��Zvl�S>�"k��}�Vp��L��G�b�:�9�Yf�FΎ#�a��H�����I�v,v�R/��,�B:P"�4cqR�Ң'�B2�$����ƚ5����(�(���/��\�h1O?�4���^y�a�r�Y���Op�Wp��ת���0,y����ژ3y�s�~广��n����������G����/��fܝ7����p��'�V�N<)���LP-��beKǱ���^��a{���H�    IDAT~�Ҋ�DÍ�w�}��v��g�$�(#��csX��:8{�$���~n}�$�!f̝�7��H8砑#��˯�������æLf��8���8�ؓ�6q �U^�rｻ���ǳ�~��ֶY\��a�\��|��w�fly�TW�|w���jR.?�dÑ'���o�m�(*U�ǱCk(rk|���x��L��r;���Q������Iy���8U����BBTh�D73=�2#W5�M=Fi���|/ /����L�K����+S�����	n�LM^W�]�\~�O�&����$PPDCC�bۋ�O��:BݔT�������[t�����qd3<��L<��'��e'�RNs"3S2���vى�ġΦ�ǥM-:q��V�������)=�f�U��0]쪋sϽ�0邏(,�{������ﾓ�"+����H���e˿e�����k5b��*�j��|�"����kXlNr�M�
�����Q�ڛ�[WO.�����ʦĤ�����b���¢gH�"4�ե�6��+��*\P65}z3j�Q�~��s%���y+�|NٮZr�\["J6֍f�������݅�n'�H�7t��Vi��rd�Q��.�=��/��f�w���F����Xr�-̘~4�~�=\t1�w�vl��k�U��V��[�,�ȣg�N��r�֮��'�\��
�G6f?������������+�/��]�]�G����Ͽ���;o8���$��{	v����
J�+��mW�.��ێ�e#�uS����-q����0r7ߴ�];��sg;[j��rSyg1`1�̟>��3Ρ��'j�i�P\SMqE5�\���{�lnV�-��:��o��G�v�9���-�&S����Rı��:�!�H��-{�%>����b%k�8�&�f�J�
K�͉!�.b���\N��"4Rk��	��F�İ���4Mu-��䲔(�a�Knx$��&R5���z�i�&��xU��Ţ~�����%�'u���j"�k�m�Y�
���k�׾t7ѳ[�����s\jk�D,Pt���hR�z�R�83����.�q�z�o\ɈAVƍ���7*	�r��D��Pճʓ���d�d�ҳAz-zR%��2��e'�y����-��o}IE�Xj���;�\i����g���l��C,��Jl����૵?PU���fSYYL��դ5��������+,�v��[@(�$��MM-�z	�Q���tѷO/�k�q�,4�瑩v'6N;�4e�#�������;ҦHm�7��ǟ��W��/71]�f4��`�[����p�\��|ޤ���\^��r'e]dw*�E��R	<6��fL2d�I�.��~�]|�����'w�u��w7{�En�m)���_ˑG���e�����Q�O>��1����q�c�)�z-���GOy�ޛ.��_|����W`?��?\����A�u�c�w7�{�+8л�"#BkS���~�'৺��"a'�q�D�{�h�<���M;s����'W��<�=�0�����K���b	��XO3�A��x鉇hnꦬ���m[))�n!�]]�K3�ѩb#�*1j��_���w�!�2v{���
���vZ[�j�,.��.����?��������1����L����=8E�TPD.PB�~;�F��1�(��P�)�����my��I������!�L� ��sO')-.T��ή�d�l.�4�� T@���Z����[e.� J^ ���ޣ?W�ߴ����}����9����;!���7B�r8�$	,��*|y�d�g4'�X���ǥ{bf8|���1��.?��"x��p�IŚՌ<��(��l��4���n�ў+/�ӵ�� J�.0��L�-�Wc��]�%%NNZp:�B��ws���{���%�6����R�-�>c������1w�Te��sG-4��>���l����Mr����B�k��f�,6�ѓ�#�5����c�ٹ���݊	^�+C��cG)�6}ks3����Jx���!�8b�|vv���X��Ӟ��HS��d"���|��������\���\^"��b���CX�:yR�%�DB����R�G]S=���C<��|e���(��d"�dm�!(�~Gg���a*�	T�U>��r_0��������
���c���������yխ�[�y���?���	�/��	!<�B]RIZ���$�%�X����P-w����6v6X��Η�5w>�z3v�h�n�Ec0Ɠ���*R%��)c9ﴅ��қd�I>Pٗ���g� ��-Ic}$�������pʂ����䠃��^'���j��qQTRLBR�t�J�ڹs�bv��7��۷r�K�j��|�7B����$��[���QVYC��!�RR衽n��Fn%�z�3h� ����d��Z^�,���Q9�^�S�R-�ʆ�bq�h��e�)U�*z����d~�d�T%.D:�PO���LJ�j=���&@*�}v����6�>���L�l>�:�� B�'�]��1�8��Sit���O1{�$��y���7x���0���h%�c5ܤR=����B��G�ұ�
]6'*3F���|]���QΉ�]B$fㅗV��ۘ>�X

�L�6���Ɛl�E펯������_SUُ��6��g�0��~�=Xi�;�Q~8/����FyU)�1�.���V2�,V-���	v�����X]�ں�*<'�);ڢ�b�.t�C����G�0L���{��nPuq����S6�t�8)�l�&B��9
�\KG0��y畿��ǉ��TW*�m���t���>444�u;յ�G#t��0f�p����	SP]�Y看�4�j�E��t�ˏ��bu�ŵMX�ٸ�@�+�8���))������ǖ�`���wÅW��Y|����������[ZZ�w=�����~>���e�P#V��[P��-�H��)�����U�T.��F'��N_�(g�s���n��{��WT��O�����b(s��GN��J.��*|?�L\%��W�+*&�L��Ј�ˣg��,9&r0W_q9��ɼy���L�R⿥HX��W6��-�M=Nj��0o��wy�eַg�V��$��왬
:�{���^��Hs��6�!(��Ku�D7fw;nR�ۛT���o�Jw,�.9�yS�$\��3�}�TȺ�U�2��*����O��<O���M@P���U <�������^i��i�o����<G'$wݰ�*�Ff�}{����Cu$�,f�I�I�׃�K�����y�q�LL��[�	�EG����T�,b����FE�겫��p_|����o�<��� �H�[%>Cé���*����`N=�l�æ/�SQ��c�����3�q|�u#?���!�˙p�(��鴎�[͇��_XLEu�%��I�}�{��k+��+NGg7�x���V����B:"��� �����,i�n�GT���۷+�E� ����9��ٺF�X��9?Q�`��\�l<H�����������҆�Em�"f���88�ǭ���~�\#	Z�v�J���w9��sPџ�n�	�mQ~�CHu6qSy�7u�)R]q����%4��Rv�5���%�Kz���#����S�r�5.��]a�����+���'}��":�?���?���)�s,'�r�uo�j����b5�3�\�9����
���4uxc�F�y�s,�B�x���६��k��Q�KJ�I<��i�8���5u
]|���`�T�����Š���-��҂�f�:���c)�bN]x���nim���\���<N�`JB���I+:I�j��w^�����n��FC�q��]P�VV�ڡF.���hlU����5d�g���&�Z���>�҂r٭K��-(�~6���W^����e�}�7߭���+���3<��?+p��O�}�/W_}5p k����_~YU�R]���_������[���Ӆ�>g�n���z�e��*O62���k0` �?�<+W����K��G�9�������jN=�Z;�t��r��������yGMLUa��eA
\ar)�l�H��8�^��4V�X�D���r蓖���������FV�r�g��������V��;{�nc�L�K�a���减�bp//f��5���Q��Fv������8p --Mjv���a�6��n�tEZU�ؠ���V�cS=�w��"�m{]� ����K$^.솝d��j1(�9�Y��
��M��~�i�m]�>`�r��|̙���,��!>[���!.���6<�<�7���W9u��8�p���	�A��3)*{U��J�u��g�;�$�	�A����k>�ȣ���?dgK︓%w-������{�K>@FΥ�`"�H��.a-i���+�����O_�����,�;�o�\s�����������_���=�;v������y�����Y�{��|�C���DK�!W��$I�$6�����?>���3��ꥏ��W���Ȧ3=1�+]���C�U�������~�/+�Yp�1|��J�����`ӦM��v3ä����+�0f�f͒p��9�8eZr�E�y�/L�2��ӧ��)��_��Ĭ���������p�C|ל´{U�ޱw��k/��"[TB,�F7�8�)���*G�קZyck���;�;�P��q�Ջ��۵����q��W�'��u'��駞�7_'
f͚Esk#�>���o]�`�F�R�.�"���|�~�a�/_�F�&Mbǎ����J�6{�l�W/U�^ȫ���'�|�_|��ŋզA���{����|���7nܨ�lӦMcŊ��~�T��ӧb�h�8�eJ��t�C-L?�	#ʙ6���f,f�bcK�Z6�W�T��S�6���]�\���˒
]Z�F6�#yT� k�Hw#%%���	ʑ����6���/��.$g��ç�S��o?e�o5r<{�r��q�&���<��m���o ]�,���drV��~k(-+Q���;j�����o%�2U����e�\RR��v��স�ɸ��^S]��'	:��iv�٭��m�A�TV��q��S(�=�w?���>Cs�F��'���gS���x�N8�$�Uܬ�K#�;y-�����Q�8��n�Sy������x������1}�L$�������NQ��]3���*�;,�C�GA�k�Wyg��\|�ʹ�DN�aKv�`ִ�����k�����_��������g�������3fM;��Fz�WN=i�H���Z�,�\3��"�8[1�?�Ľ���|,g_v;�x;y��n�0��Z�?{�u��>�1�&�������7��x�MwRQV��S�5{&C:��;w���ҫ��-?�����P\^�Yg�Na��sθXU�W]��s�;Km�x$�Z�m��j_��+^z�5�y�|�����p��l64(c��>��{��f���Q����E��W���_�s�s	6�r�������p�
$ϲw�>���w,��|�z������s�Yg�ᗟ8��S�Ỵ�>�$^�&�0a����1���
�6mQ <y�dV�Z��p�����W�~]�y����_��E��
]�]y�;j3|�p&N�Ȳe�X�n���8X=���������[4w�h�L�-�����%�����[�̝ڏ�s'VZUvx&i!v��jv�6C�8�	wA}i9��U����cY��c�J{]����pJԷ�9j�X�~�EY��&�ȗ-��5k�:u{:�l޹�qc�0�%;�m��ݴw�q�).�������F~��W��6(|2	9Å���*�dz
�Ǧ��<'>����J�
*�6����?��6>t���~޼���69�f�@���i	����'Y�f3Y���i�Ț�Zv����0�8��Cku�����gL���J9P(&��V	ہ>}�s�-��|����Ex
��+��֥�����l��Vq�3I"�:Ł"ZZ�C�����*�o������Ţ }�i������o����������[�X�Ֆ�G:��t-����g���p�N���Hg������fmo����X)G�|Kz����-�0h��XW'.��ۀ�>��3O_���_��9�s(/�`���).."��t��xCϡ���74q�57N������ES\r�e�5�[���3N��ϿRȡ�J"gǎ_)).��-�	����;������#GRw��qe,cO����/� &�:u�cQsf���#�w�'"d�Z�1� "-uq����n���+ǵ��2:��7�l:�f�[6������뵟q�q�ID#���GR�x�g=vm�-�1T��}�j5�D�>���ŤC�SSS������	GR�z�lk��C��w�ǫ�E��\TUUҧ��Q#������?#��aj�,}މs�S�{+�g��ZB9|E�X/�p�a3�)U3�T����4b������)1��n�j3).�Qpc��X%+1v
 U,l\��#Owg�T\��4��Ng�SL�mdt�j��<�l�+��%���_e����Y����ʸq��4u~��3��Ӧ��PK�����Ҋ~6�Q��6lT�q�.��ɓL�0�����i5c�z-�Wѻw5U�#���u?Q_WK����}��ۧ��ɞ�z�n�A�j4��#O^Ha��Dr�|����^IG�F:k�s���Ț��3�B�nFП����3���?�����e�֭��w���)/��no=n��g�}��?^��g�A�a��`��3UǦOi�z�ۡ��T��@�r�;e���~�R,6��>[Ōy'��T�t��gO{����?�w���?����迃[�ۗ��uۧ��	L��s@u�fL3���U�2������y{���v^z��q*W��9G!��IN�]i~�nl�㏛��/=��O����?<���x񅿩
WHS'�x��!�9LݞM:��n�wA1'�~����c撊DXt�y��W��{��E��5��������ѣ��ǟQ����~���Y%1ri�w��g��T���{N3�p��-Xu��C��#�&Դ�"=�y���C���&��λij����Ey��g�f4�����%�b��;�����߱��/��@IM�I>��SVS���pݍKI���<0�矸���7�y�n{�E"I~��)��Χn�n���w��h
�6�;m>�|����|�BQ�+;>r Ko��֭e٪l�U�ގ$eUC�47Ii�ƺ�5i������
�Mz��}uY�ذ��XԤ����*q838]�Wf�ndT�.�=3m#�i#�PG�iS'��w����qz��d��7�og��ٌ?�h!��ˏ=��eo���w0z�!��4{��2i�!*�v��j�PVZMsk����%؝V���%mi?�,v

��,��s�1%�>N�>Uҟ���.��-lۼ���e���3p@5�z�����o~������*�C�L�1��α��Vn��m��Vb2���7���O?���qŸ�Pa0�r�c+)*R�����j�ذ�,V;�@۶�d���嶥���F�?�D%ż��9v��nK�Z�{o�c�r��cf��?��k�p�u׳�{�U�qڅ�ўw)�_G�Kdk��u�y~K��S���{@��n|��U���u��ic�a�(���&<;b��J%@��Ƥ��4��@�He��������ʁt�S*��)S�b_Y^��3���og�c)+*��ۖ2�_j�+T�ʴ#�c�{2��b���_�l�/�1s�	x��T����I.�``E9}�����8�J��?�@Me�?��#�?>��W}čw?¶n+I�A"�D���
g1�*�iOCZ�Htao�N.��x�x�V�x���;R�ܧs֙�PW��������0C^Y]�̣�p�G�f��<��g�Z�|�����ZD�����=�/�[���sgM��Oa�'�����Nd1�&�2�C���Oxw�g�5|n�|�~�名���?��9����;��8���������ޡ#�Ewب�*�֛.e�>�t�m|���d�%�r4�CFr�Cm̛9�>�1�͖@3��$�h�t<Ϯ�46�Aޤ��Iy�O��%:�j���<C�F�
6�l���R���Sߺ�^�J�Y2$M��7�W|Ű!�<�(�U��f������V��H�    IDATq�vFҒ����i��RZ\Dc���ر����0]!���J߯[�����P�	"˳{l���0�7���w���آ�{ZΎ�� ��8XIr2�~������|�'�7wQV\BU�ތ8t<%��Ԓ櫟ڸ��W	g
�Xm�&�u�P�i=�F�'�NqШ��t�w(�^�*�\'�fT�W��`1t��>��y�5_~�E�+���/��%��I���JE��'�zR���f&˙g����x��g��s���;\۽4�Eȓ�����x��k/<�����?k5����@>��^|��+�޸yڥ��e��v\�ZU5f3)�_�,ֆ�g2,6�����ش[c��%��QЋp:IF�qټ�0�#�h�3{
o��'̝���駝����g������W�Oaa1����5��6����w����<J[0ȕW,��*��U=Ju��Dg�Cc}�5��ٗ�p�g���O���o��CW�X{���Z�$�U5�KK�Ȝ��$�لѲ[�΋��V�+�N瞝�r�>�G�K��]t���FU�N��K/?�Q#G`�噿�t2��j������#[~���W���>���G*gr�e�p`�rZX��j6l�AR��v���<�ަW�\q�ͤ�(����٧���~�W���������R��o���+��������H��:���cYp�LU]KW���9��*��(!�FKt�p�$F��2v����Z��%M.�#����ޅݞW)h>��T:��p+��k�,#>�:�E�$�Q,F�t.�'�"+.u�̼�W__Iqas������+�S�����y���6�pv���q��ۻMM�t�X��[?���]aVQ_�h���A/�%^Vݗ²"�>�Ɉ灤��y���
���M��G���j�_9��>�덕�2y|.N���N�UZC}g�����߶��)�x��"��3��OX�բ1���6���Ib�#]�}Cy���iV�]ݬ[��G��o���_u5N���︇/ZL2�͘�8e���}�y�u�dYx�O$����˯�7l���{�q�Dm��a�Ut賦.�㍗���^����v������)��=q�u_|��Cn��T��i&�4���L�Ѭ�;�Q�fS�c���,�z!�-.�}��wV�&d��x��Ri�qK6OMQ!ӧL��
V�X��1ƌŽw��u�\��QÔc��7�� �H\i�;;4h w�qE�9o�5�T�0k�z��p��W�p�x"IJ���p��N������7�ֲ�<��k����h��hd3a�Ar���2~iɛ�:I�7�m�U����;��H�鮯UN[��7��;7�8r���^l6��_y��^��2�b�w�����ڏ3�ċ�=�ѳ���G��(����??� �?�0w-]�S�oۡ|�K��X���3�(���znY���ٳ��t�%�T�ч�����G�)x������Wl�.�����f9j�d�L;��^���f��'_�%���9��.�n���̟=�c���c7�������#:1�4�ėI�HgbX�y���N��KKYHs9t��ck�1�bB#ĭ,�h���dƅ�ۛ�^Y����^R����v�]9wWwu��Y2�(��8��� "aT�1b�4F�9 
�������]9�����}��u�]��B��jŖ�]{�>��"}揞p4���hJ�h��^�ࡣ�+.6m�ACM�Ǎ�)o�B�/�\φ{p��2��dV�lf�.��NuU%յ5ҽ�`kM��-�(>�Z �PY!�_�4܏U����&䥼�-�b���;��*B�rjz3a��q�֚����t�������o��Uo�����GM��1å���K��BO�d"Eɤ��e�;�'RTWײ��Y��C.8�"a1�>ƌS�$pӳ�͈�����{��BU�rBr˭7��u^zo%���f�Zν�Z&����i�>�o�է���^���m�/���	�?�S!�e�}ꩯ>߸n�5WNႣ]�{0�|�;c�
)��d��'��$N��A4����Ư;��x��؃�Ɋ�-�)^1�q�x�I>_����GQ,����*;�����}Xx��Ȥ�473n�x:Z�d~����Q,&�gYT���`�g�P�2nX_<N���0�P-�5�r؉�lش��m]�2�D�N��A�8��[K�^�B B-��)�PJ*�\�d�n�F���% �t��][!����W�ȣr�gP����*�2v�y?W^})��>������{��XZFfV�}����\y��9�w�_�n�0+K/��0��Y��Gtt�Idu,v;o��&����\~�E<��S�4;�b�)�&0b� ���
E�~��bI�@u̱���xnų��e�᨜�8-
�y:��t27��V���bt���݌/����?�?C�|<r�=�+��=��b�C��h�sٔ|TE������a�R�P��_KB�^*�u�YS�{-�drv�F��_X=��_�1q�X��{��������k(h����^+�O��R�T������'Ғ�b���;��I�^UT�%AO�;v����X$��f��,$G�G��$1r�&Qx���WGy�M�^�|���|��O��j+B�4��c&��9���������
�EM���䨰�X0�rP$2�v�/<_�����N�R91zO�3�S�d���Iv��#�g~��]�8��.��7߆�n��܎��b�қ���QR��c��f�\y�9��^���7Ҫ;1��;��N���=7\9�d���ïC�8����n�n��?�oܳq�U������<�>�`-n��;63��)��<.��[C�Jd�N�����p�#8+���Y��=法/��W�-��ϵs�c��;�I��`ܸ#�j��`����-�d�J*���/�ɱ�����K[s#�q.<�d��-a�%�L��x,�a*�}�n6l����M����类��������>]��jeD&9sN'ִWfTz�jVJ���Fj|�`f�)Se�����tFH�ø}v�#wQ�.Ǣ9H
ҁ�nV�?}��e�M7K&� y9a�x��}��/^������co��Y\Ƹ1cY�n5/<�,%C��z�z�1{�������QM9v�tE�a��;Ѕ�TQ�����N�����Y��@�(�7	iY�����g�L���ǖ݌){�>u%V,��h�rD,��b?-���c�vM:���%z�n=z��̆���u����4�����G�m�_ϿW�F8�N��,Zp%�7}°�!��|�U=�g}|��&�B����j�j����M���A���PU�PP'9=KKK��aIЌ%�x���,I�����#O*ىb�ӻw�jj����yw�67�v	y�TT�����xٓ|�a)��$"g]���p)%�U8z섣a9���c�������K�x"&�t��XeR^2���P�f��������b���v�X�!�C8�
m�2�l��r�8b�^yo%Ɍ��<��o��ւUH)nꤷ�ኳ���P��\�a@������}���|�WG̻�D���ʵa.Y�ŷ8?��S�N!�K��h�f�A�R��+o~��7W�&��;��0G-e�#,�n6?�/�Ɔ���Lf�ׯO&N��K��Ti�Oz^�B<%������{	�F{X��X��M=
���-�����Zz��][G+[�o��+���7o%ᮄLS-R�x,G�_��h��hTJ����(��VP8�{+6S��r�J"��δt���l2s���C�lgJX-�%]���^���f��%	���q�]�	ǰX2ٸM��`��FD���E�mM��ҹ�`�4��$S8m2����U��7O�W�bBb�𕕑H�ɤr=�v�����_d���=���X�L:�S'ɝ7^C&�Ă9�s֌�t�n� (t�"<F�,Bz�w3�Ũ�;%N�}7���( DW�ɉ�]IYy~��΂E�RU[G���:r �vo�/���Cwn�D����j�bs����ˍ��y�9��#��~�x,L$%�	�U��3̴�w���N����NW$���6T/��B�/�F�27�l�H� ���ѣ������$bQ^�}��&���
���c&a�ʙW,�Tփ�nF��7���0�T٠G����&�9r����i�.<a�*>?1�;u�@|��}�[@�� �����"S���d�R�l���W��������e]5|�Ѭ\��W^|��/�M��G��W�~�7�Yp�_�����a@?to� �{���'�=r��Әu�F�c.k�[v�Dٽg�Gє����j�Omlw�-�ڿ/G��$S2Iz>SB��t�yT�|�����H�ע ?J��@u��-5��U1�6��gP��F�+f���+6��E������1G��>��%@DS�8ݐ���f6��]���,�n>�P5�>��tkj	�ͩ�Du����ԕw;��G��V�`���ln�m�0�X�f���cT��JA�Ĕ)����,��=M�`g�]����@s3��.,'C�%�ɒ�0|�H�"	�(�>�I�H�ض����Z�d1���ǌ��^��[%��e�Ӽs�����4?��;q,�t֫��U��3٤����${�1U�12"覨3e�0.8m2�޷�%7�è!"�v3���v�T!�rEY@a#�b��O�� (��ҋ"q-/�����E���x��MK�s���q>=�7�폭����:�8.��	���9#U�|�m{���ێ!��J9���4E���ni�۷� ���a����	���j��]�������nqR��岘�V��<�	��ؓ�r7VA�SU�l�̇k����i�`1L�x�9�p�lk)�sV�LN��fQ�9j�.��{�%�(���,R�Q����ج����%+_Q%���^y�b�.^�vV��Mfz*]Ġ*�(&�c`V����8��?�EI1�,���5�aΒ[h.j��"Hq�2�]�r?ܡ�����O~��{m��u�m�:��s�����Xһ(�3h��ۥYJA!*yIz�l�ֳD�d��x��S�[L��Ț ݣ�l<̻�=��s8��s6�Hn��.l���SVڅ�!&����jvH�p�gLt��ofok�3$w�V���^U�LXJf��WU���tXT2���J����Ń?��S���死Y��V2)���.L.+n�ƪ����n�#O���MQVVA)�'��J$�̕��U�~��=��ݾ�Y�����=�z���sIٍ5T�I s�݄������9��+y��gٱ�76|�-�M�2�]v��v�!��5�=���̤7��sfN���O���3p0�LV���{<�2��f0w�"f]~�*H��8�F*ӝ�.�O-&IR3)��ȧ�84V�N!�E)��gN����a�BiLz#vS�٠Xa��.S�J� ��bJ�^���n(r
!��%�LU͒ճ�ĳ�����=�����l��EE}����޻��=X<�"��B�hV��c���vʼ�|>+��>�=;����(���v!<{�6�̔d�z1�$�)`skrZ�N��@���f.��Y��n�^XU�����a��X��#b�,6w��J��i3/�����)��!��ɗҘM��N�b��e'�ӞK�6@$r�x���b�$�E���r�;pG|n^@�慳�\t+&��y\�ƟdH�hf�p,EI�Я�P�n�.͘z��ͯ�w�	9a�	��l�M�����&|�ϥsg�?��~�C?to�a�e7��ێ����9�(7F����l%gn��F�"��L<���,�h�����w�yٳ��T���P��J���믢w���q
��3ϼB{[T�'M�EMC1)�(�Y�eE�.B]���>�����N)����e��I�cW-rd�"úU&�9]V	"���o7p��w2���r~�i�_�H�� �Au���,����?����<h8�h�����s��f_ͦ�h<�A˞f�FM��w�{�C%c-YI'�23^��ʃ���[L=�,�Zv�}��;��R5*�+em�k��cfM��ң�HV���T���SW�f��O$0X�nA١���>�&޷W�Կ�GBs��N�������B�/A�0�*f�-=2Ij�R������1A����-X��z"6�;"U�#��*��B�&�d�
��ꪅ��M9��B��{�����Ϊ�t%so|�U&M;����8�cF�1�ٳ}N���������E��Y����7z�h���G�P��H���H�͈�z39=C"�$�J��-8�\+u�U���C��c�I��t�v�~��l޴��MA��.l��1��G�gwX!o� ������ J&M�E�W������d�\A'����nÛL=���.&A�31)���M<�GN�(}���+>ہ�����*��gM�x"L{4���C�z���ݡa�,$DL�Hx�q�6L��x�$��6e�{/�w����{������^x�/|ද?Z���KgMeΌ
�(QMY���Y#[H��l��Iq��V|��<��:���r��n⺛neʴc�u�9,��&���L7��3g`s����<��+��bb��aح"��� 6�F&�=�T4E���f�~؄��>��,'7�d�N���sY9"U�
�h�E���t6O���:H{4��K2t�0n��.�b׼�]f����y�[L?a2�|V��9�F�ƛ�<'�>^��)�㩬筷Wo�q�%�vp�W�����3O/'|��T2��egђ��p�x��78~�i���;,�s5��vpXY��K>��k�~���Ϳac&��QG��O����d��������-A��o��N��q?�͝�e�]@4����1i�h�d�#�tZM.�B�(R]����,� G�f��粔9����"hod@mS��a'��1�"���+�W���|�{="�dO)�jy�p4a2r���;#�d�/z���|�n;#'���_�q���ǔ��3���|��5�����Zxw��hf�|���,'O=�^=k�e�45���QU�_.
M�d�L<�%�����ew�9��PMu�]�5rt�[Ȧ�T�W[6n�̆���͔�ժ�&����CFO����NG��ȗ'��<J6�O3S�v𹈤�F�0Wr�<���Y�=���(l�}�ŒaH���\��k*��+�3j�X������À#F�T�y�^:¢h��ѻe!
�BI��)0i�4C���ڃ7]{8��O~���.�0���o�p��~٭���m¤qGpLC�cG�(��*)���WI���9���b/���dˎ<g_��'_����_�Mw,aٲ�1�,�4�D>�h5�/����/�;�|��ΰ�b��PEC��\2�"��E�j(fM�dK��/��F�fgw2�
�O=�\� J1#u�FA�Q�� �y\r���h�eظ����:©0z� �þPf�O�=r�p+�y��g����L�<��.����{�.:9�y4���v7��$9�I}^xa9�=C\;�j~X�5�\���&4�������o3���x�ͷ�i����݉צq���s���?��s�����1���k,6;#��pD�:��>z�Ts�G�ݱ��$�_��]�ys��L9cf��+�ID"�0�DE����G��nWt������?��4�!&�4S�>��%�10	Ȓ��"�f�
�( dVl��%��%]���K&2�f����6�"'=Vg%�bϿ���8����*��`�ϹgLcǦo��ܓ��?����ǟ�+�����n>�s��x\6Z����F{��AY������-�3��l�*H�ģ9�6�ӭ$Y�D������H��1�Kv�^� ���,6&��UD���r�Ћ)9�WY���J��M�=��{�>���%�	0?[����/ll�W��3�C�U|�ط�2i��Ȣ���Ï�0a�H��}��\���<���9p�l>�Ⱦ��e�+_�E
%��ơv�iS&�x��9�ɏ�×wx�~h?s�X���GƏܗy��/�f�I)�؅7����h�eݱ���_w���M�~9!!    IDAT��n�'O����8��í7�"3�W�x�p<���F&?�k��g���RI�B����b�u��e2�q�,�,�����,i+C����>���߳;�\Q�hf�Ѥ�	\�B���66����� س/�R	��&�,��,��9�8�kho>�{O>��睍��t��9u�̷޿g/���w7s�W�7c�o�kle�q�p*%>Z�6��A���A���b��6Q^�5嶻��s.��ݷ����0����% G�m�ҷ}��T�;�ﯕ{�!=�1�7/.�i�M6���R�͗����!�)���p鼅d�.2�*�Ndu���������X"��n�vxK'S����fΝ9�1܌d'���V�<u̚���Z�����Ԥ嫰z�d1;e�P�K�%5�� t�4h%�q�=�`�;E4G�D��bȪ��Q�wϿ����|6ͬӧ���W��%r��٧k�.��& ��z>��f%��ѣ.De��L>B8�&�U�K��IkT=/��G�3*F�b��H��Fc��c[6o�n�`�9)Lr�ಫ���	�1fҩ̻�i�v�ș<d���P�`�9��V��.�v�mm$�)������IF�4�T/�"B��xn������9����o�lZ����7��w<�cO���N����p�w3w�R���Oe%��PU<��s �r��Pհ�K�Xf攉��k���!|�����?�m߬Y�w��3�0�����V����DO�$x�8�(F��tV�R�m;�x���5��������^�w���^��VVV#u��6�R (��L"N�mg�Q�%�J̈��Q��Y���NX��@2gPV�KN��P�sr�������e�!���4(1J9"nm��Ӗ���r��z��g�˚�6�b��	��P����/^~��N8�X&Ʋ�n��g���s��1��#,��!Ɵp*ކ�|��WD��tֹ$���x�{��<��}G�ǁ={��k ���?��o��!�������w�z���`��Q,��6��3�L�}9�܋�p���v:�x�q,V�z�`Xߞ���r.>g&�\��}(;���L?�|k9|�'�uf��D����!�،����<@�
�b�薒����(��@2�m�s����>w՞Nj�M�
�r+V,[~��nqOm�8V
2���խKׄ[� �"��N>gE��	�|�-=���,�8��K���;�61a������~��9v��X��_}95^v���o���a�0	� ���&����]-��(ᰙ	U{i�YI]����5)ta�&�e�"E���od��]l޴���Vҙ���]n��	��"��Lyy WY�������n�)��&���J��Vj��v-a9�]v>/8'NY�	���$�� �,v��1�b�1l�0���+��rP]ӓL����C�輿��[n抹��o�Q�M8��vrT�� ���n�Gd����n@�<��r�y���v����a@?��w,���-m㏟8�Eg�Ēي��T�H�Vq�-��a�_�^�]Fy�?�m�Йr��G��t�Tҙ$kWl�t`w�	]�%�H�I�Ȧ�Tz]9b �RS� egEE�,���y9��}�:����C���젪<���Z�<vy�R�.��;O��'2$�
�m�I�j%У/y[9��p��ij�]����Ъ��F:y��e,�}){wrӢ9��5�V�|�7���`Б�ɻ<���DKG���~���e��k�w��qةo���w?����xb�s�:�r*�ըf�H T@��{�����t��f#G�{���J����З\�H��l��ݗ�bH�
���T�����	OY�~�=bYO��.�_���É�t��f)$�h�$�Ab�<��NA��00r���G1���SL%9�䣘q� ��*�V~�cϐ�	���]��ٷ����$P�GCYw����R4kI���w� �|�C6�����}�ӫ
����c�v�b/�[��QG���mX��
�ͬs�c���7��ʋ�����ߐ��$�qs�]��cӜ��Vr�n�]��QR�����D6�EuR*u�ĳ������9��,���dZ�,��]D�J{XM����T��˂ؼ<u��z�h��	���Řر��">�J�C�n5�vK*�Az�H��.���3g�Ncc#7n��.��3f̠���+V�k�N�n�l�����s%T�_�f����Gk����Nw" �_��륐)�D?ݬbŖ`�O���7_{x�~����K<��͟����>��#Ϙz4�NB��'l��b���
&�j�޽�#A3��*�t셫�>Dm�1|�������\�"��F/�8��38�)\q�%��Q#]��+82z��Q �K���Ύ�w���}�Q���^s5�~?��w.=jj�A(�)\n�L�{��w�����ǟ�ԋ/������͏ݰѾ�R�fB	�)�����IN�����"<j�BN���_w���0�7`
Tʈ�\"I��[��&ȃj��ￍT�U&w�/��6�D'g��܂��g��f��N�}	%!�R̸�̾���~O9��:0��wEHw�`7R]y�o��E �%�c+V3<��2��ɘLd
y�^��va�B�
b��T�-���!��0�{���v�Y��b�`Nu/N5�Ihؓvmkf��tt�S�1|D̊X���,&�jA���ê��v����D��u
-U��N�X)*�ذ)B�T��]�ߗ�&��Ŵf��+��:ԯ�X��}v�mE��k�,{]��R��(��u�Բ�׆�i���BV��\�D<�͔�=%3�j'�d����Yvi�*�7���8��Q-N�� }�Ɍ��E��E�EԊ��9�N��Q�H�aWW1�A1b_n��e� ���a��}�w����z;�֭�ӈ����{�-�y�f��@e{�c�3�tRx���*k(�]�Hkm�S	M�To��TG�p.��ӏ?���8����|�����tÖ	�>�K&����)&P��R;+�PĘVS�l#�ߢ#o���_���_�T5T��)d��V���Yᖥ)�	�;�E�_��O�Ygr���i���1�]D^fS�.�v;������{\��q�?$��e����q9�ح�27i�y`?�u�ضs��{9K�Z�+k>��O�h�i�N�������)�P.fJ�0&�̽�\j�r�I���-��v'w=Ċ&�"�;�ř��5��3�<��~l��Vvp�#O���[|8�U��mً��*w�x�x"MsX���r
�ʾ(U���ڕOݿ�r�A�M�;���u�bQ4w%�=��������YQ�I��T1��!�Ĕ��)����LQ��c�s&6v��hsdS����Y�9vd/�uA�=��؄Uɐ��3���f�	Y�h����MT�̂/b�l�lh�3l�,��{�s�V]�"�@?���*F9����}�?,���@��M)�dܘA�W�2����=�a��n�:N�S&�YT+�l�p��p���.��� G�SM0ntwȆ�.��
bw��e2�9p@��9���	Vֲl�#�u3-I���444p�Uc��Ŵ��`�JG?1ʗ�q!K�o���#�r��\��Ȧ2ilV�,�E0�QG%%l=���W^�����	���h�/^���˻�J:��d�>A�T�P"�Ձ�jCu8P�R�J:+�J��U�J$C�;�[�z����w-��?���?ܡ��o�`�ϻ��o�o�~�%gǕ���;Ŭ�X<.cM�l
�Sq�p�]2;�(�M<�Ŝ�����~���]D�>��D����K��rzA��N8n�M�=����#�`�q��l**�
U���7�ѱ�����?�Au�M7I����/;���<���ZI��r��s9y���9~��g>]�%���O����vwR���m���RB�Χ���(�j$��&���,Yp�RF>���廍����YBxB}�iv�V�����¿����c�/�m�V$�<�����������1�_ov�����&�k�棘MX����rr�S�'�r݀�%��	�t��A;K^��]�Q����#o�c_� w�`=%�'w�^k��Ɲ2)z��O�PI�M�Yz��Ck{��@�I_!�B��>�7s/?��O?�#�2��,���;dי��$J52'^t�h6��&F�%���)�CA7��ktE2�l�s����x�j������a��x�?�P��T(ѷg�����ee
��2��*�d'Z���?�ć�}���eܘQ4��U�6��وF�R�!��.�Ϧ@��#
a���Dhi��m�^�563h�p��:��=1�<���;�xl]����l�c�9���]ω'���)���H�D��H��S�m�t��Akk�m���_��Kz}�,?��c���лOٙϟ?�>��MM\~��<��t��a���8�M��
f	��>X�@4�-��q�Z"#'@ZyE�*��Ӝ����>~��O޹��?��v�����g@����s�u��>o�Df�Ա�;��߶�x��\.��a��g��{��U�
�
���)�{p���y��wX��7���&n��nN>�|���"84+yF�)�޷-��	cF��GϺZ�N1��6�WBJ�U����[�~�]ˤ�ל�s%cx㨭�¢�0]���"a)�Ɠx<>^{�Mz�a������7���K�c6��Tɑ�̗ξ��z�Ύ0󯽈��
-{~�b��a�V���J�7�P� ���R%�Q#�2������ �N��Kӎ��w�be�`	�3o���r����x�����m��k�@�Sd�IR���_MQ�1���x惯$8ѻ��=jx�g��pq���9��7H'�U�����a��~�m�[r5�Q2cQ2d��r�^UWKN�K�	x�e����u�T�t���&r�4W^u	'=�'��݄CKp��9q�:Z�%(��� �Tn�]��E�RM��2��ɬ��ps{
�d��ZNm� *�zq����g�����`[3�߰ �ņ��A�䱫vR����,�q������w�	��I�V���)���޳Wա**�!م[�6PJdsI��[ٽk�MʹR��Ŵ�g0�c�U�O�0Y�lܲ��/���^����=���A��Ü9s���+H�%
���X����SA3r=6)c�(�|F��(��ʵ���3�=zp�i�q��E���=�o�z��hh��+��Y����s�u��)ѳ����V�A,�>�[z"�KI@�V��K�k@�Z(��S��C�:q��O�y�ه�iw��w��30�>�����͜�5'��E�cq6���/����5ҿO�lNn+y�%�t9������_��`܄q|�f-�`[v5��*��TH��Kг.���?�Θ1���]t�7S]Q�����0˃�<d�#��륯�˯���[�s�]wKW�N��5�\��i�����~�U��C�5TWW���m̞=��~�97�E�l ����H��BFWp��$$�x����os��|̹�|lF3�h+��r֬��?��cN��j����?S�T������{��aܸhׯ#������9�ēQ�A^_�1SO=�{ﻇ�|��>Y�C�����%��I'������3h�x^X�%9����j��ewK�X��u6��5��f&L����u^��^{�#f]<G�?�b'�����(��`9Q��㯐ni�7��R_Q�9���q/bB>r�p&�e��(U�v�%��+C��0��)<��1�͜8��.W�ghli�N�>�FXĔ�u��ʱ�5�i����ǟ���(�R]ӗX*OK['[��ƅ�]ȸ�c��^<#��d�bN'�ODط��~�*��=6\N�a�ii6�ƾ��ٹ�w�2mo���[�њm*�lZ#����?��Ï����9�{9��y���} B�~#1Y�2�M���p�)��ٵ��];W���J�d��m*��B���C���.:t�,be��x_���2�<�L֯_ώ;����k���3�0j�(�y�]9f�����]��$����LK�z�BG/� V����0%*���USGA1K_�^S�N,��S���c�Xp�!p����,�C�X��΍o�4b��q\5�M�}'�b9k?���p�d5�ng�9�٢H��bq�������/}�7�M�޽p�*X��:���ր�-����ZcȀ:.��|�]}�L�9=�m[7q�3(�:�d��`���:��4�_LSK;��_���g�IN׹�+�?�'N>���h�Y2�CU�|�r�|������_��naCx���� #�FM6��$z���^~���\C$U"p1�����)�˯[�u��������ٗ^#PU�q����e��������`��}��m�f�Y�!���;���3�7w�^_���d�x��2z�v��,_�4}{�����,{�YLBf��8�SX�Ŀ�T���>HFd��{�m{[����򺥤�
r��M#렐�P^�k��'Me�����m1�jm%�J "Tʫ�$\��s�����	��'k>&�QS��gg�PmN�z�yg3v���z🧖��*���'��v��9��3�S������;R�<�'���w����.��uY��m&v��������k*C�ʤ{�܇E�	�������m�i��Bȭ��!�L���n7H��2�Ld�o�}w.Jfk ��##KE0@��=t�wH���hh�2����.�d��I�N���g��N;�Na�X�Z5�;2�{ｗ/��&bWL�:�x*I}}=�z��FC�׋/�(Q������,����)�$����]���mR�':t���Z	�bU&��&�M��@�9��/���~������?��;~��-�Ϙ>��gVS�܎͍"T8se�Ѭ�+��.X���O[��D�˜��p��O�܋/���;g!�w
w%�����$n���d�Ё,^���P˖�Lφzz6�%��+sI�٬2m�b7��q��뤱��7�����9�̳Y��c&�ƌ����f��'�`��s�%���Y���<��J�X�<!�!?�R���T4�ߢ�i?ȧ�Ȣ���`��C�R�]W�]�vKy���&ƌO2���%�Z�>c���|���Pӣ�PE�4��lm!�NK&�J<���̺�
^y�E��f~��$I	��~}����}�}�*��;�{}�h2�ؑ�9�,�{N�o�OM��j���[6I괅�|��wL>�<��@�F�o@��s!-�ۮP-�\Q�JE��Iϧ)�E|h'��G��V��E!/s�I���T�TSA��s3�L�b�K&�勂na�?G m"��A��G1i�V��'�V9Nȶ����)v���o���璸]��4nO����� ���a]��zFD�
�y:�I6х��f�I��˄	<��S�3>c�Y��e+;�6S��d��	B�г:͍M$�E��}<%��N�(3x=6�]��y]�sYi c�B�E�ʑ�*�^
	�e;M�ϲ�*��'�G ���|�����PQQ!��`K�ԟ;~��G9����_U��lk�I@z2.\�t~?%�CF�Z�Yi�#v��aQLb�NyCy��O9��o�s�!p�������,��o���y���j���a�#[�
�Q�(ܫ]ʗ0�Ĩ�Iыv��M&Z�T���V�?�
�DUMe�j.�j.��\J�Db��ia���㶛�>�d�ψQ���l��	J�R"���M&������g���hjf���rW>i��̛$�������Ɵ���5���S�8(��;}��,��>���$��}g��D���۾4����X�����q���j�ZYP4�y��ӦK��o���:;n$��T��+��NU�C�~��b6�ɧN���Ob2)���JN9}K�,a�7����52����g��m8a���FJ���x|��x�~��q�̓��楄��8vʉX5ѿ�D��g_x�}Mm���'�u�\,�I�Dd�A6څ��b�[1�+��$M�r���b8��{{�$�e3._@(�)
EUA��X�g{�;�$�Ma�[0�YF�R1Gg4!���b��MIQ�XlҵO�K���	�1��]M�ݤH3�=@�    IDATkN�[fϻ��ڛ���Ţ`��19�h��-�~�-��vEt�J�b6N:��QGc�U���g�a�u�qۭL�q
;���^�_���#�E�f���1K�T�l�LV(2l�TMz���,J�=#�190Y��Egl��ی<A��]C���[8�	%�������źHL)�^��(��T�K�L���#Vb�$8	B���ǎ��t���.������vɈckJ|��,�nR$��#w39	�g�t��-���C��;|�;�C�Xp�]�~�u���O�<kz;F�E�Z-B����&r"2S�KR֊�V�}�ɨ1�p��E�z��;�X4���}��Mmt;�Սa	���.ȃ����3Ϡ��O*Ӊ��XPd�G����m�)��e�$:-\r#v���.�T�6����cǌ�Y�n��Ͽ�T�*eT�������W�]×�6��!�4�N�d��E�[s>�+���Σ�#��T�X�Q*dp�\�cq�{6p�ig��켿j-m�$SO��Ǟ��".eCfT�۱N�p;���kX�ҫ7�t�.����|���Z��떦.�/�����t��2��������ı��� /���^Cׁ?x����;\ĳ���7��v&��]qH�a��G6��f�QUOg"�IH-�����C<*IU��@e5�t��It��)����&j=)w��d���8��ߘ4b�(j!'�T�*(
���t��$�	�ʤD��Ev��dF�zw��!�R����.�J���=h�2r(�t��\ds�6'�B	SI�k��I��2��ξ�9W_��իx���9�����#h�z��JTo��^ U����:VE����{ϩ�`�<F�(	o�X���.%�C����1���',��e.+����Fgg��ob�!�K��BS\��<rz^^� }э��f�Ν��)V�K~�������(�� ���)�p���z*������*�М.�C��젼�V���,�9��c��l����#��%���g��{��\����g�u"��TZ�8z\%��A��t<��pVU��p�cPƽ��Ć_��_���Ϳ�7�]Ɍ3���Xy���8~�)��5�d�,l8�Yf�8�3O;���Ȏ,�	K�P�����.�({!�� �P9��\rٕ���Y����?؈U����J���C0���=n2ٔ<L��*H�<��;����|��n�f�����(bRu��4�x+W<GM�KAtS^��V��uU!v�ه3X�����O�i�^rEcF�5�̠" :�.I
�UUKs�A�e,���0]�4Kn_�ٳ��'�Yؽ{'��\"BgG���cq��$����w?��b��i�헞d믿QUU�ju	�Ӳ�w��%zOS钙�w<Hvo�L�%Com�9���	�rJ&銦Y=K1#��P&~�����a��$�옅�N&�X���^�DDz����;[��I��_/R��'��$S]r$l���Z<RN&���+�ўy=#���յ2%ܕ��:�'���
��~�NNX��44�"�L�d`��B����T��ܸ�:jB�v��L?�$Ǝμ��8�p{Ȏ�3���u��5�6V�D�E>�¢�P�"�|RN�y��a�M�l�������3�j�kR*Ih�KQ�$�"%[D��V�5�J�E��E�B�N�/c̾�}?���_����]����5׌1f�}�����~��E���k"x����Q:=fG��G�,"�2Sd&ە��7��nڴi��ˊ��mۦ&�a#��b���o��������{�q��1�{����ٶc��Х��}Q�F=�������.����Q�����d0S�Q�����X�ZA��g��+�6�ׁ{`�wV�:W605#�~w_G}g%-�{хJф�d��*�1����Z.\��r[��Nf��s<z�5?l`��s���3��I�u�=htI�V"83��ya4�Z���_�@�ZeMuv***q:�
S�4!0�ZJ*KY���\��Z���3����P��$�]M�EWԴ/ӯ?ę�Me>��Nc����h�M�-Z\�
��3�����P?���aCX�f%��gꔉ<t����3j�$�Y^��):/%�.��ҥ+4iЈ�?Ŗ�~f�?��h�#|�շ�4�o0D�Iˋ/<��FF���wv��铬��3�zX��˾]K�:㒜�xWI>�IF��*B1=����Z���t�ы��lV����%�����S��g�f�3��(��Q�	�����
|y�X�o�������7�������v�{�8v�w�ёӧ����
�6Ė���i�_������iiܠ�b�_)8�o5�ωc�ɫ�N�_��L��u�sg�ٻ� �V�W�NQ��j5Ңes�?HZF=2�r9y���� ������քVIkK�	�k ����$�<<�`w�n����]wv����];������S�hs��Դl�k�{�<^2R�\>O�ì|��~�nK�i�QQr�ߵ�D��љ�����fG�)B���51*�*d.f6�ǏW܎�c���/2�|�صS��E�.���x����7o�"|
In�ȑ<?b8m����҈rؓ��4������l-f��6L>�ڔ4%[��.���⤠�����~��3'�x�i�.�ڄ^w���O��j���,?ƺ��JN�bO��	q��1n���Ӣ��_z��;�b05�l�&����3.����_XD"!��:�4j�,`O<:��%@C���D̨��]m�d4Ek��J����Q�������i�$%+R��H��� �>��׀����lD�&iN�����q���X��D�TAI��5��篗�t�BÞ���W2s�\��z���Df5�G�?�Β�6������o���Mt���,�O��8w��;u�^Fg2��Oyo�LF����^��~���m�k�>f�"��?u�/7��Κ�!!TU��?����8l�}���O୷g�l�����&�Og��;����?�]d��,�`!52uc�=>R3�	�ʲ4�_v�믿N�zв͍��ȯ[���k���(Sy�Y�idg�r�����?��}ƌǕr}�>JӜL�,��]�����Bȁ>222����cO�bUUUÂ�p�|�^���9���O@�ª�k���n���]M�Z��xԇ�o#7�iEVz�P�KVI*dEV$���*8���2i�jMT^�!95�-�~����)q�(�X�'��رcس�7�6�C$�Ӿx��;;�����D�\����o�����Ђ���%��#~U�3�ڂ^Q��Bt����,]������+c�U��޷o_5���+�s�ؗ/_���g�y��S&Ӱ�/�M1$b��n.�ш�� 
��h߀%;W��5�Z�A��tQ�C�{��&WwO�kW~mB������f�r�l"�t�%�D+���K��|kv����>\J0�UZzv��������}�_���S�/���`Щ���C���+NI�JMXُ͚����Q��m�b����j�fe�FBaL}b5j�ݳG���2��gK+߳�%S�	��Hn�<�ф���f*.B� I�u�yU�Z�w4�v�΀���B���پ�7{�/k�]·/f���D�e�6�g��ÒSIk�i�̝9��^�����c�9(+�&59���.���U��/gշ_��������F^{�5��5���ᆛn��}1���h-I	��&V.�G��eێ}� �咅Lzy����v�X�y'�"�L��#����ϩ�t�w��g���i|�d�k���C��T�BB6�����ыV7܈���o����އA'73S���VU����(*.f��7�N_,�!�Qx�kW�TE���*f����~��%4jB��=��؟J1��6�q�����vj]�EHNM���s\)f׮��~�1j\~���2�4n�A�뚨��p@V	Fn��vR2�ƵVTѰA.	5'�PE�n��r����^�H"�U9�n��Q�_�̙Sl��#�W1��4P�}Ea1	б�:b$.�Kr&�`D1�����N���ĕ�,�Ү�������?н{w�����֛��>x�`�f9p� �ϟW?��'Oү_?���[�7��������).��*R��ք�����g���e�ר�Bk�(c)��{�3��a/Ձ#��%^����=0�݅o�?Q�ZuĈCgD�)#Zz�f�%�"DAa9>��HL��S����P:qq��lܴZ�]%+=��$�mh�6��ؒ�N6�	KT3&�C%s�c���P�ɬ�<
�h�jW(�*�6���D�#�>����U����2I��XE~�]O�H�4*�s�h���6�\#r�PH�uf���!��f"e%��l1[7��o�~��Ճ��NVP�ޒ��Sgy�ɾ<���h��#Ay�Þ�ýeޜ����/�a�h��m���G�֫�:�&M������t�֍�����]M��6o��]�M�~������H(H���M+?�ܩ�2u����z/�π���^:�ѝ�G��^���s�E�>�����D�����0�u{�};w��3�X��;E�����|��w��?�7܈���-?�@�;o#�捉/���*��ѿqd����=���K}�)GO\���è,��w+>'3+��/����և����@$΋c����WHNMQ��7�2|�r��Y�`.?m�D��0Y�l��#������x��Q*W���4v����d�4��҅��8q�#�.p�J�̆����t��QE�m��d�:�ۻ�UU;�7e�.��u��VG��=).������l�N�v�n���R�eƌ�#9�g��۳��̨OD�#�РID0DBd��U��6��R�ףt�ܙ����Ox�ؼy���N����~�S�ӧOs��aU쥸������+�L��N]�s�T�ܓ�9-+U֯"[��M��5��}*�8OH$�u�G������^w�yu��&�:pL��x���Ͻ��[�B�v���qJ���E<� ��@��Հ���H���\ٵ�CnUxu;f��P�6�$��;�*�E����ګۜU�����j���"
*����P�eMe�2by�p)�F��p0��Fq�
�"$�g�$)]q�pT5r��b**3��0��q5�D�q����4�1��Xg�}شmE����r)nW���?���?RTVNB����j���	��D�����ӧX�~+�Q1��׬#���E���z�7l���<��`�����v��ݻ���ª�?����k�[�
x����]��䬖��1Z4���߇�ܩ#�Z�e��}T��x&�8%%�x�γd�[<��S<гi�ɴhP����͉3�Պo�r��qS^g��Shڪ�����~-O�C�EKۦ�4��PD���TA)���-o��_������@U1�|�)w�s;񈛖MsHMJ��}�)(�$�~SF�σ�����A4b��	̝5��om���&M�@n�l6o��m;~��ߧ�TP�흻���V��6ױ~�r*�
x�L�����L��.k~�{v���%b�<��J.�v��%�Y��������X���Jj����Gw%s,/. �abλ3��￉`dч�,$:���_aʛ��XRU�4��st� 9i��&%c��!�N��T��1c�0m�4fϞ��� ={>��q!�	�.q��B�dZ�ን�S\\c�W]��(�,(,w��IAR��`R��d'
K��Nq���{�	�'ԁ#��%^����=0nڂ�Ϟ�[�A�~%j|������<eD�	[U�é��QVd>ژ���R�� &�u�����֠�;$�M�v�Q{�6���0�Eh��(��Q�P�g,V�NZ�N��� C�ҥ���-&��팵{8�=9���z�#q�<陊�p{�[�H� �����^o����h�ϯ4�&-TՔb�S�Ή"΀Ř�P���H�}�jLL�(�p�-C�^W>��5S�D��79��9IQ�q��Ju�[��"��Z�H,���)&����L<C�`�U���Ky�����QZMD��$/>���Dl����"A��ъ�|q_�]:2r�`��v+��8��nf���,^��M����!�I�k���gX��2Ǝ���1b�4�J������<��o�c���jB�t���O�"�,�����<���6�5HS�Ņ�����(U� �ƿ�Ӄ�����A�c�Kc���<��!�^߂��{+HZ$^?l������y�N�4�� ���=�3��W!�V}M�6�Q�V<��p�8|���ȯ����pZ�ث�IJ�y�Q��љ�W,�~�\:u��7�6�Μ�Ì��2����v�i�,��n��Fl�il���Jts8�yi�Tƽ�iZ�������G��Kw*�>U��D"��e/��^�\/Y���y���W�V]��"[K�Q:)��^�Д���U���mEW
�'�1'%6��*����S���P]�y��������e��k;��{�_����s���_�p�܂�X����c�3����ƙ��#��*O��-U:�/��t�˖j�v��t�	
3�R�)]ZZ��a"--�Ѧv�z����4�+ܪ@;�m
2ٚ��|^���iOb���d�婠��l֤)&���e�!�:u
�3���\.�_&%+�3���*eV�0�	�ϫ���*���%/<5�;B�%#Iv�q\�%$';�&Y�T���b�aO����3����~"� 1�O@��1�;ވA��䦛{���Ji嵺�B."�R�H(G1��D��å�W� �GJ�b�G\5U؜��ב�(��r�|/�)D0���[R09)
�Ռ.��r���Q�9���^9��$3�H�8	���3g��I���U�K<e�����]�mހ'{�GV����pB���������,��kv8��^�u��.��Cta��g0�'9-��E,�vǎ�f�˯�҄WT�&&4/�Ô)�x�띌3R�Is'�˗_~�Ɵ��b����VbOMV��О	cGҴA^~�#G��U�W����`o|~��8�%d�k��*=�	�ܗ�7�e��?y{�,f��!߮�LqY%����B�{��w�<'��]�&��QPXĸ����}�i>_�sJ���k�Ft�t���Ms��.�xq�nH8,&9F��=��=d�`5����e�g�gѲ�u�8v�@X��Z��Uմjہ�gKW"�l���_8HRvz�]9j�2��1fd�0�����H�A�|�E��h��͝2jt�8ծ]�����ׁ�����z�`�5%���άW&�.�TS��H���A��,�6�A/*1��T-���r���V�fI�R6�f�򨾻KW6n��4�.�i��VV�N���T���hPdD����tR�M�F�KS f'I�z�D�a�4�`X�`Lt���d�����9�^!?iٙT�x�AŒ��h�(f�|�>�ћ��M�R�Lur�Rٴ�{U�qW��\�L���������0a�8�%��hMq�Z>e��G�s��E&LxYEfFcA�̛Gn^=k*!3�/_a��w	b�5㰘��ig�;o(ƶ0��8;��c���Č������㠷���Q��)�t��$׷h��74��Щ�u�����s�;$�͆V�ǪOp��~:�nB�U�&�S;��g�SP^ŹK�X�hm��
q�������*+�N��}�N"Ҥ�u�c2%����1L$��`�����<v��<ξ}���x�&��:�OĜ�?�%řL��Ms�<n8Vk�޽�����v���&��>�1�!�zG*�P [M��8v�Ȅ�#شa=��;3g�֌�l޺�ʊjzv���"��C���̞<�����U���X��;1O<7���#��`T��8�D��4vSBy��B
�.�����7�&7--���2��H\幇꽐@e� ���5ٜ*_>�q+NT(��]������ɨ�����x1�$Р�os#��lKe%>��rhW3��=�Ϝ4�l�����K�V����?s��ѫ��~_���e�qU֨=^8'!@�u\
v�X
��4���YX���MyPkuj'��9w)��E���HL�x�_$��hR6�Z�^hٍk�h�ŕ\Mc0��D+�;��=�ڣ���&�P�v�5�&�bJ�6���X    IDAT&!�:f2�_�pt�j �!I��x,����谘��j�#�Wi3��%Ӻq=���XX�g	�9�)΀��ʮ�Ŕي��Y�Dc1�^ai��{��A�s�N,Y�1ZC���~�.]�p��	��T�˪x���Lw.�~�nܯ$Q�6��fLPQ^���#�1����R�%���[	��f6)u�ـ��
���&L�&yt���jZ��c-�o�w��#�w`Ϲ���F\���{<@�T���;;�¥q��i
˪1;Rpf7��qb����O9��i�)�����/�c���(��"�b0ڕ�@��f3����.�٢�avy��������3e��Ty�DE���4�L��[�p�.�ж	�=�,��6[R6o�����X�$�ᒤ7ȧ<�����.��<�_����{ye�$f�[����RU�&�i�Z�l�
�1������`a�כ)q�1$gS��b��%�Ѣ� �����P='7�@ ���H�KB����2�X\�¡�Z1ɛ�Ǫ	g9ijmfu��<j<a�����B	����&d4cNr`7[��"#��NX���k�J��5�UAwD\�qϼw&}�i�.�����o�]0n����W3������%uC�|���D�����d�b#5,�ZY*��X�o�	�o8F�_�2���(S	���рQ�hm"�U&�V#�2��UX��G	t)�R~���Ҁ���W?���Xm�C�������y��sÉ�j�8���T+]~:�b�41l�(ao��Sh���a�	x<�*r�4.B̓ݾ�>_��λ�R�㒍-�貏��������	�ԫ��������e<��A:r����`�'ѰqN�:�ݤa�7x��^��o6���7�-��d"Z3�b��7)����4�0��M�K�����DV�]��j0���ͧ_~NPc!a�O0��h3�z\4�r`҅��}��˥�m�v��\>�\��5ǣKV�L��"v*��e�*4Gv�6m�����K�ĴF�z!>��"EY�jqno��L�0�gOs���<p�/�''9-�ތM��������}h�4�=���Ң��<�Rw�ـ��$7`�jщ[����t�/Y��}����̜7��s�Ǯ㔗U�b6�_pC��D��;/�B���Gu|��.V#��	�sz�`m\�Y�UMS�MGf��#/���������T�o)�B��n6׆��cQu�HA��Y��J�Rs(��2�㥸}!U�.B�
�KR]Mq��IF=E��f�>�*m����nw-�5������X�u�e��q�.��g������|0�5�n��������QX2���be�i4����������֘p��r�[nc�[j�qƵ��T��dB��t
��B�M�|S��-�{Bb"�'���O5	y��ZT!���Z�٘"ę����<k�$�E�
�W�;�3���p��I�!�#�i�yn�2qHR��oո�.��bz"�����AL���v�x����EU�o�|��g���*^��o�Q�4�ٿ� �3��I�˭ ��t'��z�NzY5�Y�)����g�XTE\k�l%�V=�B�34<�p7~X�-���4��$�`��C�:�u<5�y.��������&eன������ן��i=�	/�;ݢ���U?l����AC���(i��6��9���;y��;()�H��9���{(*.'I��~|��*b	�*L�;�租��{���I�<�W�OYU%{��Ee���O?�7߮�`�)�N7�f���XF�I�^���0�~jE5��R�[��rUa3B� b@��zN>Y4��kV)�������i�_�;u���pć'�&5����Ԩd�h�ė�7P\�����NH�O5��$"�	{h���E�o�^*�U�&Y�����}m�J-�a�{C�y���+�TH#�Rqa�G)��ܻK>�`ub��)/� �Б�[�^���#A1�S�*�1����l6�	`�WЧkǏ����:q�]����#pr�7��sǭ?q�=�pmX4�y�O���\A�n��Ք��}�jWEU&������+�[>Q|���y��k�p���-�LD'y�0�Mz%͑���� �1�P.\R�#* CHB2I�'��b1G��V �h���8�D�쯥��n_#�/r�
��tL�k���zq�����J"�-�3�p�.N�_C�QC��Lۦ�	Ք�`M���,�W Vӿ���q !Li��бcg���Jrw��Q�0�y�f��{T��;�Y&��/M`��e���� �i2Y�Ѫy3�8�h�'h�V�<�4/�:�]{���'���F���J�����|�t1��M��qc����=U�ף����_}ʹ����WH���SS��߷�D�Ghۺ%%g��,"=9�6:�d����̘=��O���e����B6�\N���Pt�j��� u&�����ǌc��qL�� ��x�צN���]�t�8�P����Z�l�q��QΜ9K��j�4ڢa#G�����?�������1x�Pʫjx♧ٽ� ��^��H�������	�>��w�}�v�o�x���}ˆ��	�⤉ul�K�����Z���[�Ք�h���<|����Ӵ%�K�	�M�T�l���C#�a��(�jj:��/)[�^�je��ו�T�Y
{�U�ɼv����LQ�����p	�S\r�C#`����K L$�#��c�m�Fo��
�1$9Մn���ۖ,��Ұ:p�]��k�{ݽ��[4b��S��w�{3�d�4�U�Z�n$��߽y����.���f�ګ{u)b�'�Z0ڒ8y���ށ?nU��l#)-]�ϒ�%�m)Вb%�B��M����G��,�����贄bq4&�h��h�uZ��*��a��!	���'�F\�섀�
DH����"Q1����#!������ �#	ɺ6hH�h�(����NR�Db�o�)�`$���\�"���ڑz$��JFz*_��H4D�&�2d��k��M7�¾���:B�,!�ɵ4oޜ�n�|�e*�AR�p&�O�"VXZ�t�V�h�c��˙9y<3�x��������0�*C��q��9�|�˾Yó�'���IyI>߭X�ȡ��(/�1c�(׀��`��'K����Y�z�|��ߎ�g�c��|�o>�����#�'���\���g�:}&OEfv=4�0s�}���@�^=��a���j�*����V�l�����<7�|a�qG�v�9�'9z�z���MZ�ႏ�"��iV���~��~}e���|��cƎy��{wg���9u�47�����ΰz��a#�����?�f�S����FX�Z*|~R3�������i�L��K���%#D��=>̱�3���1z���̜l�ѐ����j��>X���L�*]M����"�e��Ңr�V�S;�ǏW���f)�j���C4�܆�L6���BjԢ�a	T���^+�u��WW~mB�7��w�<��|�gR�d��d�tU�ej����}��suW}u"�)��.��C��r��D�A�ՙ��3��j�h-��?7���hBT�jծ\����4��+�VX�t����-v��)n��qG�j�F�A�A��ъ�5qܞJ�;��uxF5:�c�@HeB��i�h�>�a�j�q�3���d����!;�J��t��*�g��M�%3I1W�r�[���Z΁VoTY�����e�*����CJ�&^�!�������ŋ��/�<)�6"S�X�*��ʕ
�I#KFoM&�������ύ>fʋØ5mY��]�{?��2����f-�g������&�:K��|��s�:�وͬ��mmi׶[~���_#��2�V�a����z���%�b���4o�G�F�U���+WX�f����՚Ƙ�Sx~�x22����_0��c����.�\8ǫ�'q��%�v��Q�ʪرc7��{RI����%Kr��1�ӋV�@vF6_|�%��cŚ�H��ą�,Y��G��?��>��"�a#Z���?m�^^�����d���q��?l޹�;:�B�>ʝo#b�s!��];����|�1����J1Ʌ ���N�;͐�l��Cݔ}�˥�B��b.�KZrZm4�٬P)�'���T�����Ev������2�}�}��$�����0ڝJ�y����1`��#.,�D-jd0[�����t��fLQ��k�xmB����[s�����	�����bь��./��e��Ϯ��e��}�2���T!�79��k$>T�������3�"ZlI��ufB�	�� Q�Z�C�$��M�jJ�� e?Qr8)�1���N왙T�z\��2�G<n��.�����^����Q@JNn�X
��'� �F��)I�NoTs��Q�����ɱU�<|�U�8�����+�>9�����o�%��,:�4���.?SUU�&{�~��'r&�>��߽�������}$%%)��/ Zc�Ҵ�u<?j��Ƒg�&�)�F�Sρ�qU�Ӻt��r4�����G�c��׸�i����}'N�������d7mN�œ9|���P^Z�#�O�&8�o77���M�6q��9�þ��ݜ(t�XX�E�~���~}z�)�����&���ѨA+���SCG�p�tyy���,���5m@����
����o���Sg.p��9���n�A��$�z����]:�m�V���kd呙����3hu�uL?�%-�g�^��pKR]8̼>!�QD��m��&��e��<������뚱�m82�hѪ-G����gx~��O}S�wv�Ӛ�:��dF���r����~�f�j�)h]�1cR���c�"����ZU�����ua6Y���RZ�f��Mx�~Om�թ"\%�@���F�iل$�H�_Ebj�`����[��K�̞2��t׮�ڄ^�,|b�ѳ�
���G�l��J��x��+�����+��8��d!ӸF2�K������']�l�Vϥ˅<1pk6l��܅9%���%�%7u�I�Fh=	�e��}�8���S��]���Z}��Rq�c$,V24"a���JBn�` ]<���6�S�Wk֮�dMR>�I�T�D�T��UcHD�ܴj�Bi��_��ACLi���fR/'S��z���堖�M�m�A\�"�� '��f3�9����˼>��*�N���s�1���l�m�vU�9�T��J+/�2)�2�_��YmI���."q�~܊��Dg4"U$�&�P��Es_c���d�6�U˦thی���F�9|�|�����;���c���J���zV�tv�r'>O%fX-��߿�5k�0w�R�T3`�S�\E|��<�2�x��t��N�I.f�?o�F<f`�����?���L�,6�c'��Q��]��APYU�r��u������0=��ڗPDJY��	��ކysޑ]!��4�M��y���4^>�U+����8�R�RD-k�	����};�h�D�:�/ĥ����}����·�d���6ΥA�f,Y��߮孙�ya�$,ii�DވY0�� NS��:�v�jJć?!�K!g���5#ϫ _�G��vI1�Zm�q���m�Fב�������_�z}�L&ek�̩GT#tN�Z�ăAL�t4�����ӊE��R}��I�
z8��_�x��ׁ'_
��#g�kW)�/��
�uD���@@�����yT���Uor@Ɂuu�]v�M�6e�K�HNϠ��K�'�h������tǐa�ƨ.)P�(�x�Z4�[n���������c���:u����əLfvϟ�T1�d0�d�~�\V�qѸ7jҌ�W|GT�_0������|�j�� �\ߊ&������LMYw5��]]gN^M�6F�/iI���J�����DB���Oh�M��ޠS|��d�/*��&G�Д�����Z�sr���NqI)1����T�JI���HD��j7Æ�a�����s?K�8�Y�ؓ�A_^t��>z�ǌ��HS(@�]�Y%�l��Y��G���ٸ���������j
**J���Jk-{t1��ݼ��9r�k~�ǃ��Q��鯾����n�	��Kzf/����Ezf#{r0�����h%;5�wߙ΋�F��b%� �3���>5m�����6n�������=��+Gc!lv=N�����ۅ��
v��)��%3������g�~��̹�bZ�hC�'B�e\Xr�߇�b'��?}{��V����y�����$)6�����gK��Ͻyq�Df-���4n:�h�ம��K`ք�I�ѲY}��R��(%/'�d�T��>����;Yq�kE���W$mM��닊����1&eR$!2{*���v{
e��'&S�l�,Y��(9wr���тIU����nY�጗������~����'�����?vn�@�>~OA�W.��Sv��C]yj�0
R�hT*//�ez��[�Q���b���I��L�2EA�Rpz?6�2o�����с/�b!��	V��p�X�>ޏ_��mV�6i��-?)�+���|'.]NL��T�JS�����&������i�F2R�k���#�z�zJk���Fv�F=<x�=^:��K�վ:5#�K�.)��֭[s��u w��3��H��
�DB�[�TMT�B�D;�V�lN3�Y� j� MSQ��8JL�����Kr΅Y/��z9j��r�k�y��P@5R"��f�a�_���1l���ik�ubA7o�{��߅ޒLfV��¾�e�p����z���\�n@�@�ʯ0c��t&�8����L�a$����II
�֩�fQ�M��u�y�ow�����RּW	��<��T@n�V�:x���Ӥu�:3�{v#;=�^��/qC�fW��xhٲ%W**��$X�n+��O@Cff�"F~%74�ǿ��`i!]��s������������Lxc&GO]"3`M�%�O��(�&�Q�AЮy���g��))*#\^CVJ2�嗔2�jI�^�&��1��W0��(�FcA/��ϥt�ե�l޴�AO�d�Ѿ�u\ߺ�j�T�O\�P����� ^>o@5ξ`�ŋ3o�{Ly�MjB�I\���rr��(_�Un�U\��n�b���ND!Q�F�������{:|4��G�ᣮ�_��	�������ą�R��)n��S(̿��]�Е�ڿ{?����g�`��]����N���|�`��JX�EW���0V���o{c�iDe0NXgEk�)HZO������H���ts+�mF�nT?�����{���s�<��f��	L}s:i�j
��H�^�9��^��҉��Kqa�Tv��E̘3�Q�&a��,�c�[��<�]�yㆤ���DI���C
>����ҕ+�p�͔��au&)�lir�xٌV�K(��(:U�c�p�cXZZ���m�2��vq���Z}�N�|���.�s�/���Ap2���*��<�r���{̋/�g�6��+n_�ف�`!$��	�.J�d-oO����P�to�6���Ñ}�E¬ݴ��CG0��9�e�b���
��ý�0~���e������+��mԨQ*=�w���sU�1����MY0�
.�z�{�1=�/O~�7g-���AN��q�C��aFW.�Ep3�����Ճ�l$-7�%˖Ѭ͍T"�=~��>�9U���<0�a�%p�!\V��UA^����e��-�?yB5B#ƿ£�%�^S�I��a'�7ӈB!�Q� ޢ�DB~R4$=-�`iM��Hy�7�kNYyU^7Z���������PG���_]J�_��72���}�|}s�3N�8Iχz(v��l���+��xB���v���=]����+���ULz�N\($n�әH�Ȑ�Z��*J<b��������4*9f4&���dl�[l����w~<�Ց�t�u�L�6���'�͹�Y��:	�R���KKԄ��k��]FU�x]��򹫅^>/EG��W?'r�hB��h��`�%��ۘ
_� &�z�"�u���W]:K�]�]ap��)+:K�[o���7�{��U��5�7q���,\�)C�A-����+9|�~}{�����N��u�\.5l��'hд%��l���j<�?�,����n�ޣ~�@�m��đÇC�I�F�	8H    IDAT�N��:���j����N����7!:�eB���I&�$�J;{�.WF��V�o0q��1��.V�Y��ɱ���&"� ��Y4!a��O>��Od��M�ڽ8LY��#��ቁOs�rz��٪v��Љ[X��C�ۖ���֠�k))-��+�ۻ,ZH�N����e�;Hɬ�3٦u>�=���|]ɻ����1i�K4����׆���������b<;�)6�R�^����
���)xt&e!��І���A\E��ph?�<؍F�5!��K�����{���AR&,D�QV+q}H��Y�x�}�\8�Ô`�/k��th�a��?n��[3��L�ŔT��>	<ABx���*&�����kf��)�+]�ں����f��M�;���|���h�N,�T���k<�*�q5x��X��;�>;D,��խ+F���/a0�(-)�i�&
b�]Y�0����^Z�h���
��/O��$��b�CH����ʈ�������f!f�(�f����C��a̎$Q߿Nq]>������QW�/�ڄ^n�i�>��d�bֲn�L>z�M�.ֲ�C1e�q�,��q+�S&[岦��F��(ӫ�2�����"�3�w�b���5؈���*�B��i1��RLa�x��3^'��g�{�%j4�\�F�MEE5>_�^�� ?�
�wZ/�*���ߣ�����*��Pr����7ȿp�*q^�[ɨ߄�W�R����ᑞ�����4q��%Ξ>M�f�X��J2��QZQ�՞DeM-�\&�Zc�ZG8�#�"����Dsl�XTQ�H�@Ч�&iH�?z�������f�2n�h�S�#�����iX-��{Oy�ҪF���=%��۶���)�R����uFz�A1��>c�<�ͭ[Һek���{�<�G�s�!6n��'�c��Wy���4��F5���5�~n�7b����rs[�zm
C��xo�=�#F��w�4�ue��+��}�oę��2�-[���[Oł���g���i:ҲK?�RSZ�Ӧ��s`������B�[3f�X�ӟ#�Y����Z���߈]�$�E���1�Sx�&J�^���wU����8p���������)D�)0�A�M(U�]�u�d-��T<�/�g/d�;�����'�������G9GZ���tf��1��n��O?�eʤɜ:��6�X-�%���V*��j}�M"Y��7Uj�4�>����t�,YJ��}	h�$��b4ەIRyeI��+�Ù���hAc2�HTk�ւ�lQѺ�p����r��]�Κ4��:p�]����#p��ׁ[�������ϥ��S�·_U;t)��X�K�L�Rȯ��%P�U_w���?���jQ�����qv�;�+�P����LPcT)�tڭD}n-�������ؽ������������4��^�J�����־#~��w5�l���#*�2|��s6h@���)6��ɓ9w����<��şb0�p�|��.����p��A>[�s��ɓ'�5k��yjw�י��xqڜ�R#���j�`b��P��������F�z3&���x��,�C~����vl�y+i��*�M�˗/QVZ��b ����A{v0n��S�/���e�������/,U+�S'�*�xI<��!��y1�A�>�f����冶*o��;;�v�X,v��^�d!�>9��w?�M������]U���c(�|�[nlK��|Z�hFiI����R&�ɯ�ذ��WTa�x�;���N�0{��宻��a�O5���CcK"l�Mh(:y�S�b!rS��b_|�!�����
�k�iԊM��˕[��RԤ��"8������TԨf/=/��I8I0�!�R�nU� ��[48���A0�ѠG}�K���pЃ�nV�sM�e��_Ū�?�y��̞1�-����e��=9{KJ���HY�e�,:t	/��O�,��g����`��U'��*�HB�Ĵ)*ϓ�0��!�i ���Μ5�3����*E�(�J��B��Y,Ne�d����AkQ�B\/�A���!U��w���;���C�g�5Ƚ?���{����6x�~~\<���(�{Tda��E����:e\ݕ_5������QX�f���*4�Z�$4������-� f�ډ�X�8z���ط_~� �&F��<~\��CCeY1^��3gO��0O�{~������ҢJ�5m�o���v�kXM�6-�t异3�a<I<�a^}~�u;�F�f�s��j�w��X��|�=�u��
(������T:��3�����P����KN��F4V��8ĉ]���[��`BӐ����b����&Fii)��׬�Jq&���C�mf�oӒ�o�AFz�j��_��Wߜ��զ�t�B1�p\�K:�N��e<�_�&�Q׵h@�zل�^v��IF�Z�j��_W��ojI0�LA%[
	��X8��l��LΞ<ũ�O���[Tðsϟ4n�D����{7)��{�twu��g�II�ADAQ���Y׸~֜�,F@\ATL�� Q� "*Y����9Uw�<�����ݿ`��g����ꮷj�{��s�8��h	]s:�D���!�?n݆�����=�c���8| F=��68x���x����8�0�q�}fo��%�V�3�1Z�e��R&���͖,�j^��H�X��:�vxKJ�&��pB���*V�J�!fq#�Rf�dh5*�#�X�q�a�|N���`�'ЫS;�6�j8�L̜�$N�s�y�]�8�;����p	���DaL�Q��ѐ��d����b��_����P�Qt8�PS[%U�7'�`��2�9p𹘿�+#�� a�����T�-��H:��E�@3O"�C�U��,b˚V���#ݚMaܥC���C���Л�^�R�7�����o_�t�o�{]��K�ro�l`��,��2�;��T5-D7�۫�M�|M>�4����YX�t��X��CB~ܾaՎ�)G,1#i����L6!��P}9�Nz	����
�6�+�|�8Tz k֭F8��{0~��عs��o�v�{�^Q.#���ҥ�ڵ��t���kR�U�(�U�^�[��w,^�5��蓸��;E���y���ޥ��āC�����&׻wol޴V$W��\.��^
��&0D,�V���X3�Ӛ�����A`jꓓ�JFq��a���,�~~;R�	�P���`V3Ǝ�RF�"�:��ݾ���kϤ���l�ɬ�d��z(^&
�S�0��,� �$Ie��rf����	���܅p������EAM�	�f�HB1Y�p��]*���bDc�Q���"�x1d3	�T�K�j��_%h�f#��x�K��HI�@BW~Ik�h�cP4�4}eR�u�U��5Ҹp[l��n�M�L���8j����儧�I�3�z*���I$�h���^���=�^JVE��	�{��ͅ!��>��g��䖭[��#G���(~��Uoqb"dBce�������j�����<�����f��:c�uc��va��_c���r�WT���g�������K�dI�dD�1�lH�p�h�jb����$�m�����4RH��{�nvH�bO��ڑ�gMz��ۚ���r�-�{��{���=��p1��ｍ�ߏ�T�=N����t� ����n"�i�3�r�� �\��L��̶�,E0� c�G4c�#��$�>�0U�8��#�@�	�	x3V,^��m\���9P~���
\u�U�={F��իW� �Mt����ܹ��?��cGPU[���*th�
o��_}���y7��vLzk2�(~ܲ��
Pv䠌��سW<�����nC4�^��j0*�!8�4Ơ�mV�߬8	y��Ng7�1(��/��2`���9�/�Y�=WD��Ր���J�	����G��ӧ���PQ���[�D6���h�D�j(ٔtZǊ�M�(��T	����b6�@N1�ߤLf�#���&���78���DF��#��F�T:��,P,��aȘ4��tB�ߩ�@�L*Ҳ�[�$c�&�h���9}Q�� ނbd�	�q��X���#�hD���B<�M��e`HdD�'�n5	��i�#���ӶB���C�܆J�*�yPԦ�դ��Ռ�*x���W~�Y���x��.Uo�#�CB�#�s;!��Lv�UT��rBqؐ�zƤ���ٝYT��1��[R� �ꆻn�7��V��9���sϣo�A���e��#Oc͆-���a���,��Y�ɌblV$�Id�u`"������ב����Q1�����@��{�_w�@��w�o�ro����_�l�o���!,��&�zG��!�d6I@ߵs�T����!3@rTL����V�k�kB�C�5���u��U3��<�26(�<��L�z�����0����o�.X�ͧ�����-�ܹsO�ݿ?�;�A��W_-BuM�/_)sÆ�(.,�*x��E�������e�_�������sp����)�
�����yF'���Wy�o��I�ܭ[7��m+�IMv�aXlNC��Uz���Ui�b�@�o��J=��i���g��-p*�ڡf�����w�CYM�[����n��Уk�9�u����]��OT ��->mڵEy8����A8��9G�����*<[:�eaRi/k@�i�� KS����kxN+'�,�JJ$�3�&Cp*��ّ��Ӻ��.�td��~r|�UU��D�b)�3�p�ߘV��	�ΘUaS8�h���;�'�)�|y��ZOi������T��3Y
.ŎL*	�����
��E��'y�:��z$��)�����f�����Q\��pv�"Hi�ba��j������2�8�5p��p��}�n@�1(����Kz�! 5��0
G7��`0+��fеC<��=��%�A,^8L��e+V��y�KFն���܆�)�ؠ�]p��d��y��#�ȩ��9>���t�)%�L#�AL���_���4�=����
�@�������o��z��e�h_��V����j�g&lv~��Ȕ^�F�11*�q܆�X1>ib{�""�B�����u?��>����u�#cu �1�HUCNc���kT�g7b�E��U������	մn��&��� �8�V�¶_vয়YIG���E�ؾ-<�}�v�[v�={t�Uc��/[Ƅ�o�]�>��|0K��6�C��|�ݵ�'����1	�E�سg
�
�󼦦&z��pe4"�	��`FX��m?���	C6-?4F�� 	�~�T�LF��A<��k8R���Jg.5��^L��n��V	���}�[n������sυ�n���"��i���"�7��bҠmt�e��V�HHԢ��f��j�#���5D1�6�����*8�~�
����F�`��aG���2:h�i�ݺ��&kjE"�Yь|���Ȣ��	���V��;t�"�g�yrQ��5��q��x�ʦ����������i���D<�d85�K���=����3��`=�t���M�`��M������&�Fu��K�ӊ�Vm`J��hR<��Ƃ\Y�L(�pc@Z�m[��Z�6�+��eb�,<9>4pج���qZ$i�8n���P������|���>Z�n���VX��\q��x�9��0���p+���᭼���H&���9+�,�.�N'/E��rv'2�􉣇���?om	��`Oo!�5���ԩ���R���P�=y/6-]�[w����f��aŦ�?4�Ci��R͋�8�tyK~�!rcuu�l��X�a6��p�B��d=D�p�n�	G�Ò��φ��F^��p �W-C�v�DXf��a�!(;Q�/.Ɩm��Dy�H�N�6��j"�ێ���0��ѳg9v�_8
#F_����H0��7p����mmղ%ؿ�ؖ���	��J�hw:����ѽg/��b	��
�-�������#//�S���A�ng���	����׍��s>ȝ�{D#���Q��Y���m��}8xX���>X�
�i���A�R�� �50�qn��e���;�lƀ�t#̬�Ʌ6�Eq��ʏZ���_���,�o���
��*3�4����ĉCȦb04���2;�����Җ�M��X
�A8cN[\Ή[-�X�����	�J%tw�n�X�FbQy=���\t
��Y����3���Edޝ$BV��wQlvt��PT�`�d��"�P��(L�6-V������A�ϋ�ʒI�p�ʞF$#q����eQ�v����O�l3���
��e`s8���Ĵ���łPc=���	��z��!~۷[�.]O�?�"�t�3�FUC'j됆i��,��&8�.�^��}d6�o3�I���Љ<�8^���$���",3q��I/=|ǣ�x�k���R�7�[��7;ʗq�j������8��h���i��77?�yqk��|F55V�J�>�͟sL���?�0�9>a�^:�4&�F��$�dB`7e��?C��p5>�1�'��IE'�FY�a�w�P�Lvl��J�Ua�{3�ڌ���v��Q8� 清ݧOo�ao�w�3����x葧U-8x�\�k����+A�%�}zg!�Q ����}�@�_H�c_���۟I���5���l����m/��2�Cg�w��8��~H$� �"�������p#^���Ci��fM��!.@�6Ep�������:׻�Y(=R�P$,ۚ_�������D��
q!��(/V�Y�j�0I5΀N�@5d�1d�����#�ϟJ#�!"�u	,��Nu�ǡdcb�ѯgO;|��Y|��u���d�v�M1��HI�G�oG���x<B�N�P\T�-[~��{�	��H4��alذA֬sǎ5�BTVVbɷ�`��`�1|�j����v�BU����>/v���d�V���h�J%|�t��H��1���s;j���Q/ߗ��n����_��l�����'1�/����ǋ�� |���ظ~�8���{&n��N,X� ��o D��}����P���K���*?��_�h�[���֭KPUU��'�K�x�W�����\px���f�kc�[��a19�&��H��<�%�F�o�,�&Al5���BX��4	��p�y�^{�EX�l���[z3��OM�t鷻�����ݜ�����h��#樌*f![~�*���bo�r�x|'�N�ӡXڃ2�=����}�h�q帉�	g�4:�:�X=�:�
��z�#�iD�ǌ�_��C�q�U�aȤ����ƍ�e6w��Q�]0�<Bd�y���Ubڛ�bղE�p���{��U�Va�[q���y����P�Ђ_&���y��^}�Y�<	�+�[���}�.�uCMm��ۻ��S�T�i���'U�E�3]\�}��&������/@0ĞzN�"��w݋��:���B��H�>=0�oĂ��W;]v������0Y̢ڶd�f�[u�v%A��J:	^b#k҂���D����S�)@��S>6���-*��}�t!�sh �I1��d��F6Q�;o�͂3:w�;o����r\z�e�hӮ#JK˰z�j�޹=�x�>��q�>|0srs��a�X��AAvy�Q��;K$ѭ{���"��nD�~g���
��/�/�w�ʫ�b��i��?�������ħ��� ���I�a��7b��h�`�|n�O4�W/�m۶�9��B�j��}�D$�vm���G��M�ϧǐ�C�˖�����ǳ>��^�w��~��7�ɿ���ɃE�|�k�]�7�x#/�׍��B�Z�j�g�zƌ	O>�8���
�\y��Ӹt�hL{�L<���?�SD��r��x%ePNh�7��mf72���7dA�#�B�`��i�� +��&A��"K�BI�tX�֮�x�{o<~w)���-�{3�ȯO�~ٜ�{�%Kh����w>E��m-�&��瓀N�5+Ɯ����[�n+A��K�VO:��L%��x�q�|�m���E���8�� �a�B:k��Mä���5 �P�Vnxm�=�H�    IDAT���!��i,�v9~����QfۏT�!����,�ِ��~g�٧��-n~�m\��gc��C�ڼ����l2K��w�p����)�Y5r����Q���{
#/�T*tYB�o��r�Q��d��x�sM8�׫ϙ��U�"�Re/}�c�`�
���(�v���G�����
��Ϳ���۷G2���=��ҵ+^x���7�"���B�A��a2PD�(]��c$8s��Lt�r;��n���SF#|��H�x�5!��>Q���ө��r�#UX��<��m(����ߏ5k�Ⱨ�����B������<p�]x��[E���:\y�58�O/t�������_/���F���{�������C=$B>_���9��������������`̘1�-��޽{���O�6�}�ރ@]�@�w�s7^x�|�t)�>�N�:ʚ�ڱ�[�����E�xӍb�tɷ0e32��|�J���$|��l����H5UU��;E���;�����e�]��}�b��������k?|��r_0q����}�=��~�+��B�.]��'�qƌx�71v��%�ع�#.���6p� O�h�.{cF�:^G�����i2���D�c
����=����4�yоؚ����u#O��Ռ��f�-z3��{��K�z|)Il+?|s�����I�!���(��m�+tJ�rf���EE%�ۘ�,�����1�N�~�G+k��ˇ��5⪂x��B�T2����L�����nL"�Ƣ/�``����8g��g�GiY�׊�u�?���;��6z4P��'��3O>���rڏ?l��^�u�ݹ�������t2�d,�d�cF]��S�t�r�F6b���ܥ�$+<GZ�R!Nw�� aw����سs�T��zg��C��B �ۚMQ��ܽGo|��b�F9Sf��h���oa���9,� O���1 ��Fc0$��WN���ӑ6ؐ���٨�~��K&�Y	���өꀛH�c"�C��T2	M\rr�1[œ���i5O��̈Ǔ���x�,]�ل�EE���$̜=_���֣ϙH$�]��b����3O��k/E4�?���c�C��]1s�����w�)��o��@�{��{���M���O[%yRL&L�23f~�w�N���_�D(���:~��;�/�PZ*Jր����ߞ�>����v�D�.]������ǟ`����Q\\��/�cǏ�c�v�UW���ɘ<m*ޛ���ф�K�����'N�?z G���5v�X�~zWq���N۶mqN�r��;~��s�=׏��[6��o
�_RR��o������c���O=�h<�/}���RP�U�:��̈���'� �"]y�Ŧ�ߢ&�0��K$�͉��kN2b��>��L�h��d������>���-z3��o̘1����	�,��~UG�a5[Pﯗ*���Z{�Hc�Q\�JS�k��˨��*"mW��~�F��=@#�Pm�:|�{V2��%�S�b@:�@2� AC�^l\���8�بΞ�	�m��k�8�`������p8�@]%�z�q�x�}fQQ�L-�O����է���Z�}*�g{b@�m�8�=
���"�����m"��M�C��h�%2~Ơ�D��j�JI1�=�$�3��B���XgD8�����Ed_y����TT�	����ǰf�:�ti�
�N��O?}��̚�9��^��-�Un������T��*	�|tѐ�8D��l�hK
�}7��p�QSS�ݎ���ڽ]�w��j����Х]'����pyܰY=8Vv ˿�W_6/<�$6�Y��a������q��kp��_|1�V|�A����/<���:,_�_|�@��'�|��
j��OJ�p�"��\�S�.J��۶m۶m۶m۶m������m��s��g"&�n�22����V&�粹T�����n�ȥ[�}#Wm֍O(��3�`DC��n3
&�����eq����T�~x�S>���o�*į��`��3�v�ݑݼ�@��Z���p�h&���RjY ���v�HA �H��h7����s�����3)�h����h�������e~��������Tϝ�ޛ��w+�!�l^�V A����E\�Ñg����cx>��_7�d*4�����-n]�Xu������sa{z�T��Q��NH� ����4|�
�k��h�b��^��PUߗY�/uu���a�B x������T���o����}O����9q�O�*a��H�Jj�:����	~��6�|�>��R#�[h�۶)�-/�����Z*6m3�v���m&�ģ�Dov�k̤��@Y�8��Ⱥ�R�)��%T�o8��jqԤU.j0@�ɨO�2n�����5��¥h"���zԞCn8&2F������vT���K�n�&��F�$�9r$er�D�2�A���h���,�9��s,)(}��"�8�g�oy(���q6�G~_i�Ԩ�yP��v;�RȎe�y���kÓ	ý&�RX�߭��	��b���b�+���F�|٣l'(ہ��o�ۥ��azI�ZEҐ8�a̌���#��rU&�(	����xσ�
�����	�>2 �ҟ� Q]1�|A����1d�O��ʮ�R+��c��3������4�-[��n��{JXt0��[��x=��$z�!A>�iK�hv����Y11�0R���F=���»"-�l2���ǐ%������|y��>�V��&|T�T���e(���D<q��Х{ɑ��7����w�c伱H�`���N�r��@@)�>OA$0����RQUG��Ī��~� y$U�4��"�h�t�.&�1[���r��r����,��%���&YE(����4r�(]<�\�.D\�7�ԉ��S�;4��?B��Rrfh��qdFz�S���?Y��3t~T ���'�v:�:��?']�����&���u���~�,��f���7���̦��)�{�I����󼚇�����̮��׼�cQ�l�������DMCE�����ٳ�6:a������aGB��*�!�MjOy��-�Ù��K0��HIp�8� �A"f��3��ɖ��!��aVwƓ�FLEjF�����Yd(���Qeu5zS� +�ZS�!T
Tt_�,be��q#�bh�b��t�.&41B��(0L�#��,�>���_wk?ܮh�2��OD�	S3Se޼q������S�FN������Lvu�/x��@�� ����0�.�G��l?�`���d�)(_t3��B��ES�g#��Ř��YG�@��f�"���tE$��z�u��E���z�1za����!sF�#����K�C/�(���;���W�s)y����{=�\s�'�N���?3�s�NrU�6���5�Q��}�d������	��q�j��o߽D!b��'8���g���]^b8>�lg�W�M0x�����FRL�T��}=���p�M��T�r١d!��1^t��m�w?�T/#�X*0��og�
N�u����5���z���^ȎǷ������_ݎp�}��k�z1�y[G-^�gE#�'�
�n�I���V�i�zD�cFb��!c7�S��b$΀EZ�:�'�s?¨�����S������
�����K��|)X���V)��X5HV�xt�����Nqw�W��&�Wɋ�_����Ϟ[FK=.����`��R��D���r�� a?:���`���]]<O7��j���!2�\��zǔ
SL�6�D$@�^8r�����2��mI�Y�r�����2ǌ�QM�Y�Y7EJB�ɐ5�K��Ы'�˝��J��9��ǫ�����@K=O��t��VOd��}�"^DҎ;�j���K�`�J�
3VCZT}�7b���p�j����J���|����]j�h��+Enw�T����\h���	
�e��dD�G�>���"
��	[�~;.�b ��$����a,e�d�R�i�|V�p�C@P�'�h�� F�B/�{���e$��φ+z�4�4:ʄa,�E��裱���逖sB��	'�{˛�W_�L#'x��9�ؤ�x<:c,|*�9�S;�贀b=�.����6ˢ�w�S�]v�ml*��V�G-���n�F�v0A�;T��=B�{Q7���v=�O��
��Z�y���y�
y�����+��}��h���t������A������Ku{��y��Ͷ�g�`�s;!g�J@#a'�&�n4/` )�o�j$�M���Y�q��Q�^���2R��c�󻵾�}����w�0�9����y/��J���e���RO�0�8�L�ub#�y�-E|�8a�� ��p��-5T.���>�R�b���c?��`���>1/���drOwR3�\��PZ&YΖ��i�T�x�����	zݝ:R��������Mb��ɵ	�r�u|�Q�ߏekEW��\ı糿����|���������0K�\�*,޸!rJ>�Ė5A�C�rv��������̚BS� .lw�}eeU�Z��Gl�58E��>�q�?�X����ES-¶R�')a�l�Dyq�W4��y��v����[�����6 �!�o;^{��	�d���?~�5�)NH�9�dТ�o=r��E�я���?���x��Rٿ]�"��Q�>��{x��Ǌ��@�A<t�b;��DA؍j�c�X5E5�]w\>���Zb]ae���|{_O��&�vZ3�K�0DO��L���v�\[9v�4�:Q�w%�ǥ�D���k�Y�a�=�C͌"K!nFN�-<v'�G�
O4񐺳@�����>�\�N����&�e>��(5%���I�'#Y��7�F�;�9�܅PQK�%�O;+u�	��Ys�Ꮺ@a�p�+*+K���5�	����7�J#��d�eHW#���*�j��C�2J��6��K�|n�����9ՃD��\��}�����8͙o܉�H4o#&vH�M������H�I��D��q��3���!�5q�2.~�-����:���ׁ̣[s,�kN:��Z��U2�!��d���ZVZ�T
��[�!
ڙ�zܱ��2�9l"��`B��LVO���}�d5�y�<�=מ�-v lq�c{�!��:9ٿ����`)6y��'oC2���J�n���f��^���)��s;�;)�*Y~��宁���� .*TmP^Eo���*�&4W���B-M�ڰ�W�!�������]��IK��B�!�R�� �I&)L������gz3!��$��9i�VjLIE-j�2�N�ڃ��ڶ�`�W��'i��H<��@��i�zߣ9��}��p����ZXzT�0)�1����V?��lU��g&�M�[5�V�7��"Bᰕ^���ӡ�u�����4~�M�i+�%$Y"�{Rx���T�_"�=�	sįM�������Z.�A�W�g���AS�a��S( w�\��\]M�;kY���j'.��͟tU:�oac?b�0t>%�1�J��\42�2:>쫭~�I����Em�'�������-n�82�8�PS+���Мx�O�49�F�\�r�#o|���g/�����5�w@�
�*
pSe�O�z�*��_M�L�9�<+�+z�ja#���\S�!�6�|e$�HV�D�ViJ+�v#�f<��J:�p�
7q)�Zsw�=";�bIUs���O	Ȳ����V��lB���o����y}�
f,M���AS�h��M�U_0`���e�7�ߏ�ɡr� �g���IMg�'tE�~YL�\&�q���K���*�U9�|w;����;��]�ֲ~�V�z`J�CE�ϑ61��Z"�%�ת`ϼ���)����H��r4�2����9����n�Q"d��A��w���tl����HJgj��#Q35c�Z#r٩�_�&#Nʿ+C��w�޸^��Q�4j[�
 �����?�{�b�'��Y�Ê�����5���0B����RE+3W3w2���|DosW;U5�!��c�P'�)�'�<��+�>R�%�P�+p�=1�]a�¥k��1���߾�'������<�懮iB�#Q��`}�D٬��>K1��@�DT/eO(���	�����x[!�bb��'8��۷��1��D��O����_��q���8��"~"q���1�`��ȖHe��o���5gh�|�o8�HѠ�g�*��o���؊J�a�y=����cu:PB]ۊ�� ����f��S�%���^ݵ�(sN|4;��eȈ
*.��F����ڴf!�D�$�6�O�:�6�P�H#��.$��<�����D5�e�$��̲lqZ�ԗ���$i#{g*�v[f�y#Y+`��`]����v!?;������#q�D��d]-==� ��Oܻ$_8�L�I�g�)LP/����ּ��=3.�JG�ۈ�S.M\x�<�94��Ѥ�܄EC~Bč�z&�bJg��be������J8����gt���z�>G�:?5���o�R
���p7��&�dUP[@�)��ՉiK �~�2D�tؼT�H�Ԫ�kj�MK�O&�,�b ��Z��B��𾧞!�&��ӫ�(+��rk-������`�K*9�ꔜ��,ʙ1,��k���F�T͌�OqY��|]�.�֓�US�r�[��N�ߢ�4eZz�qM�3��y����v�|\ޟ�mh������ŉ���ٌ6����]|�M�	��8v�B��HT5����h�]�=��I&����A��DR�8r�tZj�^$F�m���L�<~�Y�w�=DG7�D<y'ɡ��na�u��IrB���3Q�=�(��*2G���(ŕH$�h$�;OT?Zn�|B��%�VBV%GS��1�$�Z��ϫ&��@�M���R&�w�`]�']
g���<��-��֥��JeH*FɅ�HH'(�s����aɆiJL�� p#T�Rf=�B�-l��,����g�6�}b�b��'+q���'/X7/�視���o��?��G�V�E��qOu��B�!�L��B����A	(��$�OP��¤�q���͊��;���ѭ�8����9�r�3آÌ�D���~����	F�� ��	;�x� [�;Mo�{?l��B����+���V+�����C���
��XE��T�"���K���4������W��f4y�u�U��G��[��0�:�Ν&���o��&L�,���Y�G�n��:�g1������XGZ���{��:�C��X
`����S�s��S^w}�~�@��.�
V[AO�Z2w��q.�����(	���"k����^�M/^̀N��"���Tu���؛���ݪř��Ϭ:;��A�Y��O"@�n�$�d���CK4q<w�PW/N�/.񌙝��39��f�]T��1;����� �d����^�,�N�֊p1`�x�ʔK'e��<	��!������Q��Ȍ�u���V�-eԬ�ǐ9�n��)�kw`��UHm*�T��V�T�y��
��!5�_Zc����|'F&��]zjO�E����T1�8U��dc�%T��J�vLVKD�\��V�
է�=��_�}�%5%Ve�b���>~��$�BA������;^���ӡ ��ff�b%"������A�d�z�����&%,O1�����x�^��U��f�ߚ�7|�}��p�6TN���j���A�L����A���~�Jg�[�|�Ӫ~����r�~�<O�)�򢭭�<%y��И���7���\L�Zz��n�p`�m��g*���8��]R��g�t[LV1`�O*!���Ow¸�T�.�l�#�Da��7��7y�AC>և����S�����^�;8�;l�]k��E�l����O�^/�@
&�cne�ܯqY��^��kXw&���c���c�N�}��qp��2?U���F����C ^��L��:� C�l�B{n�Lꇚ��4�;0=������ސ�K���LUc��Q��p"0�C��zC�]A�c�=l���M�J&�ÐM	��@�."*��'�f�����t�}w����l��������ӣ�rV��Ҥ�_"��щ J�����Ճ�hi����R���C�mQ�� �Z�W�,�0���
��;�P$�����`�::$p�^�&<�2!E�´?��\N��c�ۚ�!�L
���L60N
\>	ӭ�K�&QAHݭ� �o"���4�3�VٶRJ�1m���ԝ��W���P$B0l�(��]O)�9�"#�d'#j=}s�7���El�ltZ��7<���_��F�!�f>F�l��? 	K�~&wvJC�ht?���nI�����������?v�֍`��䝵Y��>�@i�]�E7n*
v�j�!�p�*�#�����AN�'�t#� ��q�ڷB��w��,���|�;Uy��+l�	|�`�M�mJx�US�ˠ�$���.�k��Vy��Z��6��%�#c+��23s�IIex4fi�d�_<��%H�2�ΦF��j�e�خ�`������s��nC_���a�1YW[ߏ�G���8�F&��5���ty0��X�@�Yo9��>����LY���K��Ǌ�������ʾ(�t�2�岈�(���8/��nù�����m�-kk'��a���K;��1ML���G�q���ai{"SS0� �Y������3Hg���k�U1�_̮�҇A*��挡"���5Fm��5M��JLS��W��b"�"%1���:�C�M~�lY*M��+r��a���A
���%z�O�C�J�2ۛ���S([�
,Z�Y�HJ:A)���g�";.@A�}�X]�Wp:��޿���W��IŦ:�*U�+��qh���'@�ٱ6v���T��y��CE��-������[���� G�x��O���E���v֣�1�kd^!��#Gf��'��D0���B�M*4_y�6%ZDu�=lh��8i��j+��;.8o|�T�N�P�� Z���w�Z��}$�R�Z��:H/�Ƴa������o�̳�K`t�2�3��L*R���������y�=W5Z��*���`������bgP��:̓sM��<I��Lؠ�(�Iy	����j���*�zKZ��N����ݜI?�	}*>��R������.!�h"a��C��˓��K�߂�P����� �����i���h��/� q������=���Hy��5x�0�)#�ԓ8Enhܒ}�SU��\1"T�U�P��l�,̡�bjT�OT��V����o�yA
E4��I]��W�Tt�S��+�Ҫ�̤����6�(�e�:0-xH�:?��hA������A4�!�P����_tx��`��:{�K��Ed_D�	�M�w^��&G4%��QH6�)b��ğ7��:�lq6~ޢl�G����6��V�p�-iD1����2pMh43e&Z�F��5d!2d�]�"�/x�M�i�_�
����.���L�A 2{�q���3�W��b��a(#� ����=��K�S�\���lCE�z��0�����qo	�b~!t�|��%$8�-FU�R1�,\1|��'�ezK|/U祐>�xwV|��t=�.��n�KA�
K �����i�1ӓ;w��dP>噐VD�[�����d)����ҞH�T�eT���;s>/%N��Du4xa{�x��d���J(���C���ȗ?��L����(*���r���;θ���'=�'W�MM�q�����q�,�D�W�S[�g,z�����P
� ��f�!��+PI8°���AՄMC_0�� �*zO��X�#��s��Y��"&`Wn��Pz�&q��HHE��7��A*��+l�{��oaҮ��";�_~��x�;�EIQ�4�v��Oj�P�s�	cI`�Ͷ�SA�z� _rD�s:�Y���(�ZTeFj𷭎�[� ��je;)�l4$:d�^KU~�8�佡~���B���:0�8��"�/��T�U�2Bn���g�["�:�b(T���'U
7����hmZb:�w��Ѥ����qmP\�a<�����Z���u9�.��;4X-��螣��#����`cɑ�9����c��>�����5�?�6�<v��S���G���H�?X�=���>+e�ż���'�v�:���z�9�����vr�]9�R}��՚]�U;��K>۾h�gd�|��b��U�������S��ݜu�߾��8}	�'�~�����/��lI�ϻg�������F�VC��<�] t��ٺ^ �	�~�ȳT钸g����?XB[w�h���>�b�}ͧYdV�q$hV��買��1�>�Q5��1�Ph˂�����HƁsn�Q/LoΏg4��L6�n׫X`���0_{pw��g%��F�!��5xP��4J/Km/�RN�C.��WK�H�&*6�
ѮΘ�\y#�A�Q{�6�(S���6b�`��c�͒c(��G~i�c�`�:l̄5�!�Q���OJL��eQ�XFsE��-z(�Qc�iBSP*��儬�9�[w{����	��}�]�TJG���~c����|��������w%��!���G�׬�#F��+��oY���Nʁ��G���%�3�@�94��r�I�n�2C�l�^�d3{��{v�z+�`O��T-�#Y��ѳ�-D :�!1௹\�e����@�N|z��>֯�P�fT�n�-�l�jZ����e��h88У��pA��{��W�܄+����v?ܰu;�d��IO��'n����z��M�|P���1G�,uBe6�55Rj�C�-�Ɩ�����O�QRgC��5���^Pa���O�Ļ��t�E[l���+�	�-<IS������� �}��c�>��b~�&/%z�Ƞ$�N��ǎ��4�N����%{����n���"vfh�C�]���Ҿ⥇qg�;�p�Zϟ�3?������#�
�K�����	*�C{_iP�@��d�B+��@�y�)_7[�ʜ�!J�ǒ�$i�ZkRp%�F�S��_R�,�3��]�C���WH.g/��5II�҅i�)&�fȕz� 2�$5�(T�6b�;*��|UaƢ��������Ǘ{n��-ܢ��/w���1�,}s�Q0���� �� �v��&H�/ߚ͵�'��րqu�j�B�'ڂ�s�K��l��NX7揚B�>�L;*���a1��C�����}���u4{,p�鿥W���1��o�"��ì�;���_\e�/����!���`���vw�8�j���"���\��*�����Pg�Y8��lι�{b=����Nu��r�*�/�e�\�y�QӝPL���ɋ"sxB.�{��SNY�R�a�Bl���kՅ���H�s3�ꐲ�`�Թ��z�Ϸ��C�ބ�>Oޫ�N	C�9k�ਙR$t@~�7�����1 Q[Ծϛ��?����Y��%^��+�����n�GE��c�!��JТL����Wh�$8����G�FWK�k�qMg�x�$}7 QOQ�o����;_	�܏��6�x����'��6J[��vhmhaڥ(F���܀@Y_�NN����Z%v�����k������{+�p W��D����΁��e2k��RƁ�-`s�m	7m���(��w�
�~�6��9�% �)J�R�?��n^&v�cC&�`�T��[7[�<�Oƶ�I'��JwL�WG�a�wJf��/���u��
�$SU�*�A(��c��Y�E�k4�8�F���O�p�$#Ǜ2��p����� �w*L6�(���?������{��Tc��l��l6h�#áy�~�gB?:q��1F6J�	IEu�{	��ޗ��z�Y����'����[.J_�u���(U�\�WE����NfF/9"�ސ�4m�)�¹[�t���w���� �WZ�G��|kox�.%�*(A���` �꩛� oibo*��|�}KK���'�rqdy�_�uk<�蒔��w��tE�}z|������I�V�q���Ë�SL�/�l'��@��sg29Ռ��NQn�F��9i��f����!�ǃ�#��]��Ѷף��X�ѩ��qa�u
�g3��t�v9Q�K����c��O������G>��nE��#��&V�p!R�]�\vĳ�ru0c WLfD����g�C
��j�G�v�P��'����[�p��_�ЃӠ��$`@�>�T�lʻ���=\��.]0�������U�4a��\AV�{�
AE=�{��,>C^�cuM��w_�Դ:�Hv����3�5��۪����?����!�ş/ ��y�������f�����8Ȗ�m���~i�M��3�qjY192^�1�@����<G������}q�n�v�w�c#�q�/��ba!��@��9����O!����8��j:��������EA��g�.&V'v�x� ���*���󔫞j�v���$�'\�>"���;�&`�B��t��w��NO��mD�������q�A;�py�����^wbT퉾����YAc�MX�m����G�,�&2���3
{��z���,(���4;\��q9'4���	�ƛ��7(8�aY�+�셓�++T��&��)Z���+���U�� �~����#V�u~ɪ,��ޜY�{F�wB�G/9�J��4в�6� �r�U�@c�53��6{�o^lnC�,�35^��a��2�aw����`��R=��7q���r��d!#̯.�����H�vjW�М�d�0J�YD���zJ��׽��ݼ`�it����Wi���&�e��:�`bjr�8������}�`��kP����34`����q�Un�.a�ݏUD��?@pܱ��)?=H%��]�>}g��"#�d��٩�"kIR�b8? ����!2 �{��"I,XuY��R�Ĵ�@�7�����>��W��BH;���"g��xx�9ϰ�Z2���*P~�`"�g/	dxl�-�^�}<2�axM��]��J������ç��A���i����c�%����G����F������rY�Ѵ�ʱ���`M/0ZT-%5M�N�0TaL&_Hry��:E%��,��a.�9�"�����S���ս�����pJ^+�X�̘�� F�(}r-b����80i>�������_�@-Ӏo�Q�y� ʰP *2�/�dRC�eSIVR��35\��p���ڒ.�v���ww&]]}�-EbmD�9�?�|ȟ���C�9ZN�jl5��Y�Ò����bY
}������J8��������OAπ��*ׇ���h{�_�;_����؉���^�Q7�[n�</����;���`�L�t�0k����YО�����/ �����_?���� 2cO*~����A{��)��z�,`\i?
r�C�jСm,�����ɏ5��e�\hʫ�+ �m/EfG6اH�n�^�U>�M�![��}��"d�����}?,~W��܅l
A8/UBR�_��O�u(Pf��d����r�w�B���,�*�������c����h��`�r"�z��&�]��������2��0*B:�3��j��������5�̛�H-�QA�O�jwO.��?"e"�ڽ�%�Q+7yg�L��֡����'j)�5�I�����ZS�A�X�
�~6}�u?�'��m��u����}b�&�<�%���OY3���g���H����j��������HJ���h��ҷ����`B���b�K<����߿}{��"�_Ok
�3�;8��3��.k=��6vc?��.���Un�ܹ�֬�LH�3��E���Ӧ��;���z���6Gz�q�4v2z	��C�1�ð
�@aJZ�S�9��t��(��ܝ�_�����a�ˠB� T��p.]OUWM42D�eW�lF�Ծ�[����@���o���w�������@d��b���Ֆ,X�v%����9!9-.�^N��8��7\�z���=�|��S��~�ͱD��ϓT$c����;�B��:d�)qf#�g3u� 7�)���Pc��R}C�t
� �ne4��C���u���j_���� ���_:���Az�V�ozBOP꽨���U�U =ZS��I�t�k��u��������-��y���*��U�Q��7�1����h���}_WV�1�o�#���F��'<F�cm�a���ܓp����xL��VU#q������C-N r��Q>=�:������^q�xB�1D��

:�[Ϛ�W���	�`��V�12
l�,��,P��٩����X1�̲0~~dM*���.���t���~ada71
9�&h �;s�R9怃4�YCD���5 Mg�v��SH�=_���L(��� >�HM�k��Ĳ�`W������,�Kz�,^��*B�ǚ�3���b�cv�Φ�#F�Q�5�]t���AD�r)�ϥ���D� jǮ�����`3�A��Wx&�3��C�|��n�my{�m���0�[�Z�r�(sJI�(��F"����(H2:)��5�0�A��3e7z*��8���fRj`������c��{�Wf2>�M�'r�)�;~i���s�0��,J�=C��R�yj��Z�s�D�9yk_���k�J#�M�e����I��?~�X|f�ա|<�`t�Brb��%�� ���<Ѿ�6E��,	�42�@���ۜ�S�-~������a�\�]t���CR�<ƃ���ԎӺ��0w�1�7�݁?�*>�щ��8ذ&$��L�'N��9�{4Æf�����]g���YX#0���� s	���@PVΈ)���N�r	�����H�R���#f!P5�?�p1zLC�Ԅ��y2���x�Ər����ҩׯV�~����#e=v���*JgTH�.�TX�B:h�ii���>=aT�ݛV��Z:"k��q0w�I��DC��i���4V/�!�5�p�r�q|�[2�[U����ņ���x�x�Z��7�͝X����M��b�0%U|y�9qG6	mZOs�ԝ)ME���âE���@�r��6�Y��~��2�O��O����C��EM �x��w��ϒ�mP2�{��;�S�nf��Ե�"��X��~a�J}�W��ikznR6ԪVq��~}@	E��#��(��+���'� 'X�,��S���ݎ��x�����n~�]�X����>�ڛ;����B�c1�_��~���~?�B�5r��$��2y�G�ď�D��ӎ�)Y�a���UI�Q�K��2a�d���e܂���`y�wZSK�S��<U�7�P����R=y����z`4i������)]�u/�F�H`���G �{�Ƥg�����u�S�HI��˦Thy���j+P�L
[�Z6!P��!����;�[7p#��Y!�\���lmLG�\�Q�4��?�8b��Q�˯�@ꚏY*P�d���xW�t�d���:�Jew�F/��xQ����DRAAd��N�I�.j"*���w���Zg�}�z�!�R/����g�����yQ�:ݞ�p���:l(���w��x$�ND�N���CQ9-���p2 �J��H^Kݧ�N.%����.F#���F�sD"��P=�(:=k�R�; �f��>��-���P�|�Ӫ��w+y0�a���ߋ�u������tI_ ��j%����p&�"�E+��>>���&ˮ�B�fi�����dΧ�C]��!����t����c��]��c�6���FM2
J»D5�U�<o�:��j��4�o���{�����p�y�ңx7�mZ'���X�D�N"�Z�m܌�Δ5Mک�[��Z�)��j���0Z�7,��P�� �s�yn�s�~�Y���鄐�:05�\�բ�e��[7:� ���EC�2f
�<��G�'4�����E`��K��@�=�A��%k;۟c(4:24�-��S��<6����j�G'�mt˔Mh����c�ʔ�\h�fjCp��6���ߓ�|j���o���䀿,��O7m�כ�^�[_��cfe�V$��y���l�Z�ۥ�G9��k�S�Ш���ܪ�tC|��gķ��y:�|�u�h�������i��G�iȄQ^Ri�m�8��Y=����:9�V7u�{�{ɯ
�]�An~ �dX���]��T���ƥaKT�-w4�s�s7�M�Z�F�-"|^g s\z�d)[eH)������	�:��
jb����9H�lt��Ƶ�q��k�^�s|_mTz�A�.Y�B*/��0S��f�a���r���s�Xq�Uըz�|n�IJ����m�CIA�zCe.�]�l˷�e���r�>�>�P��3���A+'l���` �Wt�����IM�n��g���
�|���Ǿ⥒:�z,�D�(����-O+�9o��\��_��J���~��oet,~2� ���[��{	��8�&�	�Z�.L�8@[�Q��A�,Da�l 93�{�I%(�B̀�]�F����П��� �����!f���Mอ��I!L�+�9g����(�4�UPU��A̅j�:j�x����:h���_�pR+[*G�4��j�c�>�F����0gP����9H�<�.�9�
�]g��C����2�ndy�4n���	�V�3
&������9D�(��?1`q��#HGEa��lx������<����c�}���[�J���E6����m�z���|s����WB�	����&�O�L�TD�b^\g�~>��\��x<߁~=�<����k�clv<E��?¨7� ��`�2x�H��s�Q�j5bKZd�.c�w^Y�Nb��j5�\(b�<�sPf>��JK�_�����UF��г	�MS�9�����Ȃ=�DM�1S!������~�VF��s�y��� .$��+��M>�쵚��$!Vd�uz���V��c���Y�{o��xW�|���'[���w� ���:���3t�����L٩E0���"�=��'b�b�V�� ��d��ֶ�/�9�4�X{A�)"5|�2G%l���;jM��'��b_���^T*��T�?4�T.�tޱ�(�9D���8XJ2�R�AyW���Ū�K8��|��fS�w��Ԑ����)�bxw�]%��Efۗ�f���� �k������P-쁀�	b�М�p8l��N����v�8���-��}�j����}w�@+�
é�uH��qK������$p�Ԕ���ŷ#!���|��"g��N9\�V��c�`�T� @�?�+����~��l�p5���Y{�&ԯbf.�fm��c>�nE�F�%�h��,�"�1�Ce�t�HW���ap�.)��|�(G�FLF7�L�_��<�u[���v�:�h�ZB�q����˃<�}�Ι���O7P�z������0�)�	�_�do?��t���)�5U��[�7b,d�� U�f�8J��h�j�߭y�����Q�TC�i�)�����'�\�yb�<1�3k�h�?Tz3��E��s)��^�K�����R$^��@��;�������s]ɚ��&�\յe�$�|�i_�v!�g��ϗ��M�wL��ީ�p6N�rx���U)�)1_�)^}�"��1%�� �oS�p?t�����8/����VX�}�������J�:�������P���(��F�S���6���m�rٰ�1W�В(��;fcVVLQ���D� � e���k�k|سb�Z��0���Qz��B�>Jk��r"�.���Lǝ��#G�*X �&��[�g�/xf�o膅��9y�1i��|\4vYO7Zr���U�`2������᪖
F��e�33{�E��*}a{%0n=����M��	���L����u�\���C9	vtT�=�L�3��{�xV3��X`2!>��L�haÉ?�i!�}��tB%H������w��.�����z�Q��<t�թ�jO�c&ѯ���!un�����I��I���ct5^P��4X�e/<�]��P�A� ��*�@(���*$\]I�d����=F7�pmw�a���k�h��:z$�U9�F��Z�,���cs��w{���0�^r�*��bq��O�Fk���6~.�a�@[�A~�����e
!���5�����A�q�oc;v�aW�p����шip#�S�d���(!F#�h��T�^��2O��=�˝5a*�՜�����Y����g�a�d�uy�]�,�(Z/��MБ��!�
͛���]K7,�a�_)��Q�� �@k���ťxu�hL�:+W,5��S����Fl޲�ϕ�Y�8]X�������3�_5��.�P���/�!@����?���_No�!����#���,T�S��!!��2�@'Ee��!*JH��V�MY�B	����R'n���gKZ\3������B��������r��Y���Iuοӈ���1��N,�T��Ŏ��Ź"�������N�f��b���8q.N�.�Ӧ���=�p���3xt�������u��8y�4��\�Ą$��0�.[�>>���(tZ�8�-�
��n�-G�.�a����v�]���]놗_~����+*�+�2�4�n(1�~�lP���Q��JpWz���o���z��"�T��w�E�������t>��vF������F�>ZxplLe�� \#%�W��K��r�
x}N�c���ʸq�y�|��ǈ�&VM��&����Y⠋M���$�ez�MSG<�%%%�^nk�C��z�XPR���G79�.�/>�Ic�Q��C�D2�]l�X*}����A�sY�ʑ�ҷ.���t���ɹ�T���[�ݴ+�v��W��T��ˊY.��΀� �`��u�40���U��4��J����%[���1�/�r�</l�SS��_�`4#�e�������5���st���>�ݻ�ô��_���Bx�,_��<���*����r>g^����P7%��t=R�q��=(+���#�x�Idt":];n���~�mD[�l�D�O��r':M[D;�q��?��Ն���t�Oĩ�����QkA������z�}pSX��t*���)��x�mK1��˃+�[L�IV������Dqa^5ƏǮ[�h�,�7m�ׅo�Z�Z�aǑ�X�u�>�о��#��+���/�x���S���w,�v�����
����^���P��65%����W*�9@�'�Xdu*�������ʞ\��\��e�]
�Xn4�^�2Ō��^�������.+~sz^��\ ��k
�_ 3eb����3:���N�:�Ri�t8��w)��k��*� ����i:�
dB� ��7[�x�
'�9��N���_�Dlb"|n/\��gO#1.���?v		I���BNv4j��Zu�P��p{8r�_#��1<7�I�ҩj%Ǣ��"f�x	�Q8r�$�л�ۛ���/W�RR���"�Ȋh��z�����@�"G�2�G���!=��V�*]nD�3N�65:R�/�Xi����P~n�>���4�D����`�7��N��^/�L����*@�Q�o�|@���L6QW�9Y�5r8S��~��+��kZ�I�4t��.��n�.Yv�_�+A�i�'{�������J�=�O����'��_�5�r_�Ӊ�d[�9���� �'��1�A?uz1eJ��S��Y܂+0��.��pJ�]���(��_�����	�QI�+�Ye�ץ�%�/^_��=^�H��O:M�#প�Gz� 4�~'	�D�-=d�����v'�z9�U28����t*�vRgkаQ:���k��]�=~޺ǎA��)���^^�f͚����݉���������Y��w�M7wf_�Z#�yI��<�Qx�4����]�h��&�.���ȱ3���Mf@���k|-�T����Acw��p�u�b=��E��^	�Je,Ǣʤ8�*���t�sz���|j@k2���:�!�����t�
�i��xi�襀N����=�K��
���(���!�S� '�F��{S�a�/Y׵�]hsMk�m�	%E>�Ť�o�Đ/���S��]����x�nݺ%W��v��zB��o=��{��;,��$%���O��NY��ᑕU��؃C_d�\�I/Q;+�$	�eL,�^V�.���S��8�]E�*�p��`�Ub�����6G����w��%N�[� He�V��ų�-�a�UXٛ��5�\lp���qI "�V��k{# -V���rZ�j��'O��3�3��v$&&��(a=�4�\��6"Eee�X�a6@�/v[֯[��ݻa֬9�h��O��s#�G�F1t�P���`��8��{�J���G�r�~o��Ѱqz١��R�4a��:�u�����I�
��<��9��8u�d�CgA��'R��|o�j����Ru���i$�p+ha����u�܆�A=Q�uB����Pr �G@�
�^��J �#x���}F	�s�Ч�5	{�mg@���^��l�s���u��V�l?|���E�N�o��aҳ�=���}���W!@�o������2kV�%[�m**-�/x�y�I�Nd�;�����U��	�	(e�X�[��dUK�.����X9�E.dP����.f?�N���( )�j��N@J@K���j�EշZQ��&hw���*�E��r��$5��-����4�JS�V��>�dd���-77��hf/�w�R�B%..�3㋊K��y���[p��I��m'�~��v�G���^JI�)`u�í3#���)u��aZW��M��g�=���$�"a�e��;y�[$����݄��9�%p8����Pk��駟!�܎�u��#��
�����m5<��P��Ti��7@�s����M%*t�*��"�f����?2�������Bu}sd��0"�ݠ�PEɎ���S�(�z���U�WA�� :��$�垟��F��9s�e�z���X��F��b�ӖЅ�#�!c��l�6�!@�?����}��O��ߜ5����G7:�.ÜW����c�V2�=�r��	)`�$���xddd(�� p�B8a�"`�A,��N �]����r�xi���b2�����F�,{�t�8&�C�se�*'l�y������!t!˓hP���0���"̨��ƞq��Y9�-x!!�u�z::Od��ɹ\�111�*U��pyС�(��b����𣙸����|��D�}�����ANN��p�uͿ�=sW��oX��z2S-]�Sv��q�U�N�;������ѽp���D<��SШM��h���д9��Bm�
�Ȕ�N#��=��~�)bU�踨B'Ю�}3U_5���t���̺�ѿ/7�Q����_[��&�#�i�) 9�]\��iiʣ��Ae��E<7�,�;�lۈe���h�E+p�Mw��2Ae���Sg���1��
��q���OMM-�o�[B���:!@�k]����P��hӑɶF=������M�l0z�{�쩜jF�E����X4m�T�Q5�,؞��1�P��%�NB �}Z�fW�ryه'@w;�eN�a�Q�T�[�\(H����PƷ��T=Q�d�D*�wr��`�p_�E!9:������`��]��H��MR�J�����h�w��)�腸Πײ�-!!.Z� �}�6��QVV�����>C�v퐜����$��E�ԉ��v�=HNL��߬FA~<>_���\�g_�F�޽ѻ��X��f"5���_�v��I����l���x=�+-���Y\��D'���+a**ƣMZ!����*��)Ɏ�_!�}�zßt�
&�]�\@W|��L�����C�º����Y�A��⚧G������S��� ��𛊟\�ӸT�X(�c���Z��c@��D��Y��cسOa��Yطw;.���v-Q�v
�ed��[{"`����"�7���ڵ��~nܸq��Fzѿ��_���;8}��s������2��4^�$���a@�|طo���0��$%x˖-�[测���!*WY�J*U*�e6���d5�7d�Y����td�����&K�T�S��1��ɢ��C��"��}2rT�S˶��a��ztЍ�fw�n6$��R�G�,� ��޽{����A Z� ������=��~d�h���:t�}���>cM�����S����׷�*�Eaa>���~M�Ӏ-k�'���F���?l���c�/Ƚx��wb��`�i`Һ���א���{��Bv!z�ꇸ��_�1v�H@K��tv7{��0�E%MC]�W����Wtq�ʠ�� ���j_j �]�+��"�.�� ��s�M(�i� �J��G3�hj�R�S� t�܉~�jT��6 EP����s�"�{�f���[0g���qW�l���w��e�+`��
;�M����r�m�t�kC����~ϼR_!�W���{���f������5�|�i���0�-�S��p�]8z�([�DE,�kd�!z��k^��$�I���;�,Q�r��̂'�$�����{�s����V�A��!:�́)D��j�^Z���BLT{t�uK��Pn-�^�A�ŀبp�*�]^Xm.�Z�px�9S�Z����eC��#L�AJb��C�5�q:�n����4���TQ �·����.{�F��{�qq1H�[��	�˃��� �~؈�˗�[��������-�܂7&N��^��n��0m�س� r�p��i�3�}<;�9N�ۺu+�L�l��]���Of����G�h��qgg|�nΞ�A�^}��Xg�C�ݍ��-_X��r'"Ic@qȊ��v����A,�Q�~��M�p~^@���h�4R�N�Oº�ﹸV���{�6�`O�E����A�"�ưN��Q,/���S�L�+�vZhqBݕ�A�Z���Г���DyY1b�0|4����̟���w7��E�1��o9p�|��%V�h\o��
�?ps��6�UvA/w8�:gݞ5И��>�����p��e�ruj;v�2��o�~"#�дYse>:��E� m!F��6)$����6Υ��T!;]v�ѿ�b���Z�Iij�w��׵��=P±l��ɲ�f >2I)��5�/+Dv~.�j7nm߂G����"))k�ߊu?l���%q��x!PZZ���'�wW�e��Կ4~´?����|�r�h����tj5DE��~R��l1�p��ol/�Y�#P���HLN��d����Bz��[�طw?-Z��n���x���p�M��͉��F���e�Ͽĉӧ��U(�V`��ߠG��ӧ�����`Ѣ��ʺ�VBnqx�x����=8r�.��G��h�� �}��]�5E|��Z����z(���Ao@�H�C΅�>1��ǠzEe�vF�b��8�*��8ZJr�	F�����re�:M���8�2�����(T�}(�9���B�^=���#�M��+ѱ����vEG�T��*m��V�3p9��i�(����!�0�\l޲<�	QhӲrrJ���Yhͱ�E�̧B�K��[����4NQ�5�~�Cz����k�|�o�J

M�'���g������5ɲ���Ç���d��	�jݦ��q�,meģ���	e"�Dzשb�	�x���J���/"''�OU��i�Y��]?"JW�ݻ~�5�݃7&��w�|�&QF3�7o�
�Yy8u�|�b���ܐ����W�{����gp���І!��D�������3Ⱦpz�O|o��
����f�΂7�����F=���h�?�' �L{! -��~;���"^��F-Z5��D�qdAJKKǉS�p��)�Y��w��Q�f��`wT����A�V���Q��G���0`�`�]� y�X��w�ׯ�rrAʸ1�_�ƍ?�ȑ#HJJ���W↶�`�~ &)	��wR��弥ЕXqK��{}I�(p'�瑧����AQ(*�����>?�ڣ��ʿ�BכF�ċ��Q���D7A�k|�^���e��f�[��ՠAr�Fh�.Qw���+�=��m��񹺊nY*?���l����	�
(���3�<���NǮ_��E3��݆��oĖm��sy��EšԧAf���'�0�o���P���/w�Wѷ��^�?qؓ��o��ǃ[���M_�1C�h��Ơ�Z���D7V���AIl"����>���j���t:��s�[ο���8y�d�qz��Cpb��ϑdv�ӿ/�C�=�������?Cdd2zӌf(����S�K    IDAT)���u�`�o�}�X�h6ƍ�>_�Qc&��6�����-�p9��8p��^��e�ߧF?�4��t%Z���2��%��&�&�[dD4��#"-B��dm:t,�����$t���ۃƍ����_�#V,_���0#�&�i�4l�~n���ի�M��`��}��8̘=ޜ�6Ə��/��z�kq�|@��xs����K���_.]�ӁܒR���F�� 11+�/����u��[�Nк=t��:5�[��4�h�/2�iZ�e4m�b�l�l'Ti�q����|��;��/ 5U�n�+�ԈLN�9%q�ç��6��14@��%`��G��s^�����'Q)%�6�4"~W�#G��;�E���Kg�I��HIL@�VעC��a�#@/�p�؊��z�w#>зe(X�O���MB�~u^�K�jڒ�mg��x}�Cꁘ���tT��\�K1�t����h�T��/�\Z��0��.+8ie3^�=�ji���ٳ�DeSeH��Ť������������sx����y�i��KLAZZT�=�s{)�<�w�r�|�>>�|�/�*]4�~Zg^��pΞ=���C;n���{z��v5��5���R�3{>;�Uᑑ�H�O�+�p<C�N�Y�����h^��b�jw �n=X"b�e�6,^���vzrJ<ꤦ@�g����q����cMaزmΜ;����aȐ!������?���~��?o��snC�F�Q�uK>z����
�˯{���G��\K-��������aρ�б�<�*u/����j�X��t�PG+�?��)'�P��JPU�C�i6-m/>C��gC5��ˁ�$=����v+�\�c �ޯ���G� ���2W�u��Q����B����BAN6F�~&N��};�B�9 ��}5jKT**<Zh̑x�ű8�U����6�>|��m�4)����!^�� �|,�Y��y��ܢ����=":n�&����ٿ�S3�5�h� ���*�T��4E�27t�S���mI^u�YYY��Ϊ�I//+�����%3ct�ZQ�FM[a¤��պ_���Q1hԨ|Z-��8���"h�ě/��\��1�	����xq��К��������iŁ;x��m������������B���{Dŧ2xS�N4;�^G�Ah|�]ɘYY����Z���ի�Cn��� 19%e6�>}+��)n��6�z�[����P<Pitp��3��B�鴃����\��Æ��%��~�w����x�١�ر#&My�=���<,��6b#�p�l�o؈G���ZX�`1�j۶m1b�H~M�I��0<[^�h'�\Z���NX�}��*�U!�E���<�$�"@��^23��&ڝ��]��d u����3�i��TЋ��8��g%�~O	���E��M�9iȶ�r�(� �����?�ӕ�p�7#�v
4h���z���}�e��-F���~y��~�[4h�w���!��3�?q���Mޚ;��O6�RRPȀN=t���"&�V��>r�7���(‖��M�3�n�r'�]gL1�̬�e�:�(6/
B��B
�S�N�v�6{�=���PQ^��-3�a�Nl�uN�ɱ����8�>�<sY�9�8�q۵��,���:��M�Pa���k�rka��G�f|�,*�Ǒ�`ҫ���[;_�#�C�U���u�����RSSY�}���S�)d�T,�#ʝ ��L=��5j�ۑ���� �v*�z֮�?lڌ^=�g@/.�ELt�6'�a���'�&���cެ��Z		�3{6��V���Kpzh�GtlΝ;��	f#p�|v���>2Q��X�p1tzڴo�Q/��
���Q�.�޸J��n
y!�Uc$tc�b�����U��x�u�*�R���'m� p��)�x�����aћF͑�_�5*��*��J������眔��4jx�.���ee3�>i�$�:}3>x-�5F�V-p��Y���0ꥵF�݅B�m��w��t�{2C>��J\=�� �깖�{$Ћ�r���,d
�)ѱǎQDobĨZ�g�w㴦��6���&�\�S!2��,A��:P' ���z�ܥ�):�T⥥��x�p{��_;)�&�.ؽ>�V�p�|tZ�"���X��>wٹ�0�԰h�h� ��o�0'�.��h"���״ez��aߞ��j|0�HI�M�2�0����F`�����OOO��t�J��\��&[��G�aʝ�V����"�nj*W�T�RPMR��HN��U��G}w�}��QZ��zuk��v����h����6�]n�j���󚗗��^{���EJB�-a���O��s�qq/<�
�qg[ڿ�f}��~�X���(��Ѿ��3v�i\.�ʩ�&@w��q������z�!5�B�<Y
�yz0�+!?��)r�y��+���.��#��F�\w��_�q����U���&A"�Tp��ύ��\<��3�p�سw�}m �q1�W/�ݫ�@e�@Y�cѸ^�-o�t�F��s:�?wB������Q������<�p�s�b��ʊ*)�E��B���E�޴9��)^��T]S�*��5�t� �*Z^&�1�U+ �/��D�zaR��7��$9h��k�Ώ4[Ă!�AqiW3��N�
��^��������s���0��8����~�l0�TP�I�M3�]p��HLNe�[Y��� H�Z��j�)��ǎ�
]gXX8�IkԘ��6��鋨�D��<���k����FРN-�ujس7v�N�GN�D�N�p��<?r���PpX+�z�w�bc"ѣk���^4n� ����O>BqQ6�e�V���#6&|�ˍ��?�G �SD�kt�ۧ����5\>�ʘZmP,�^��<�-	ңT��4�O�Z�4O��|^/W�Ԃa!�V̲��:o$gpy}�җ�z�4�7�EA^�~�I�]0�lߌU+�a=��hpם���.}p�l���7&�o��
}݄g�?��k�Is�k����x^��kl�()5�z{��w?��P�(/.��b��c��LT�B��(���lkºE�!UsUq�r��Ӎ���T�����>=8-�G}Z-�CGU/E�B�N��)24��s�ˬ�<>N9ӫ=��'0� ���r��r�{���~�W�¨)��A*��8��7�Asu��U�SR�'Mf+..����ܹ��r"@=����u�v9`4����MH����Ɵv����bl޼O���}�&
��Y����jJ�|��[<��s()-��ؿ�\���������U+�����>0t()��?x���p![�lǓOCRb*��#��������"��u�&���Hl�^r�#%y0�r(����w�?����Ѣ18���e%�׫�@��a�������g�q��)�0�y|0�#�%��h:^����[�U��Ѫ*<�X�v:����MF��G<>�i��E5�:�˜��׀���e�Z�Y�mkan���/b��g�7Ep_�|�z��>���覯�`���l�=p��	E�F�(3�	�hik�Q�r"�w@�S�^nǀ�'Ϸ�Ru��j8���PI�!�yUz�=�J�8bj����4�z��aZ��x��N��=�~���XN�=��-ft�y���D8�Ѣ��z�ȑ�(,,�Ł�sp%_/��v�>��h���y�>8=>���}�zu�*�u��P��K����j�_Z�f��G��!+7��zu���Io��U+q[�1��G�ܰg8��Ա}X8w
�5���l޲�{�A�zi�j�;q�=�0p�@q���D��"K�˛�����HPS��⌀Z ��J$�>ZD�e�2�M�ٮ�
��g^�wu+�<�����9�
���~����ѣ0��w�o�N,]<}zuǶ-�1�������V}��;wc����h\w���_��k�=��1�5��O�?��ܵ���\��_���3��U�e�B��0�.��;X�ݮ}6�I�|�^u�޽.997\����=�b��|ue^zp�;����Р�H����F+I5�@��U���$pF�%�XJ�O�Ia0����2B���g�{��:�E��V	�Җ'�+1T��ޤz�=?ː�
z�'��ƍ��s��� :1	�j�D�X�1�?��6��7t��?
��Τwv�g/fa���0~�h��Z���c���P+9	o�6?�q�QHOO�9̈�'�Ι0h�8r��8����Fxx,.\�ۇ��vŀGא WK��}��@	p��@`�����'�p�$]d�Sz�T=�Ǯ�܃��j�V���T�K@��O-\$�^�Y��b�ˣ��;o����X��#4��������ɋ(,�#2�.r�lȳ:؇�:#�ǷFz(D�_���B��ϝ�+�&͟�j���[r/fE|����@W��Q��'�k ����"��VC�L��Ѽ���(�).t��2���栙��Eī��6�y��R���ʓ���"��Nzhb��*�v�jR���x?[	�0�ЋV1�Py��b`�n<�3O��U���T7����i�B�'�8�ݯ��b�����@�LF�k29A����e�К"P�p���1"�ϝ�w�|�'DZ��H�W�M�#�"99w�s/�8�/�Y���������E@qA1�~�-ޙ4	7v�~���GX�`P�pC�FȾp>��]���t���xQr����#��3���P���6"9m�q*�-�� ]}Y�z@� _êGe&�Tk��Զ�����:/��bλ���1~�8L|�<�+�C��0Q�"��K��Uka�J�9>v���D�7���q�{��⮖O�?~!@�����o������l��Ή$@�g�'�����'U�gϞa����j�*ӎ�ߨT�"�U��9ϛ�W�HT�WF��L��_.f���6ѯf�����Ŭs7!+7�����2��Gq�"|�hy'�Q�)�[R}O�)���d����)aᴽ\���Ѿ2S�Q���D�S�;�"��h8��a���M3##�	�e刊�������s�a����xIyV|�O��0#2�7�#}��w_������S�Ga��s7i:�Z��
�~��p¬ע� Z�=�܊���%������棴8��68�t�� 2Zeb��Sa���=w�����6��(���� ��T�UJs����,��~Y��j�`�� -�g*���	�/=+������E�R;J.�|n���0�W0�q��a̞1� &2
u�6A�n�PP���c�0}�|DԪ��������C!��w����p��m���B���Ղo�n,�ɍ�d�X�}v0,�qp�U���~�����d���*>�m�vj=��v41�T(��9VU��e�KG�O'ʝ�6@]t��^�n������$����"�������>/���h�$	�4h�:�=>aâ�2JP� p�����։�dh�*o���>g��G0	���*t�ߑՎz�#"T�@����� �j#�l6��/&��U`��0e�D�ׯ��sg0t�8��n\ߩ#&�7�������左"����԰���>s��?v��F�f��+�Y�	�Ǎ��r��sz�釔�X�tR��M�6x����i�,���I� 2��,x�����\R��Nys�[2���[�7�ʝ_-%��-����z]�
=O熆��{��&U�*���*��ƌ�
}��hެ2[�F F����X��g�ݺv�E�丵�����s��j���_W��a�-|�c���!@>�/���af΍Դ��e�
ٶ�~Vn�����p��vT-!�'�$�#Pg��Z�)�����i��4��/`��������Ʃ*�_�ԫ�r<%�tb������9�A�ۈ���SO4=U�t,��ۥL����X�N�X����������(�?U���Wiu0�l-��6��V�D�åRa��C�z|�d�@�׋�hԊ���/���ۃ�}����F�W��MP���0�lv�6��%���o�:8�J�u�!>Z�/>��O�����]{ѭGv0��n.f�_�Gпo�wyJ�1"�_iO�D���>���/�(@._�ދ��F�
pW��v�|�=�U��T�ә @w��Pܼ��ɺ�q��aʝ��?[�����u��踆0D%���SP����]�ѮM���F����O�շ]Я�k�?��%K��[�{S^vN,Q�/�q�ٝ�)*T��6��"A�MT���9�p�E����a$u�`��3�gU��]9��vHGh��R,��R�B@���8V��9��Do�Ga��nPT�^���&��T�$�Sq
������1�|�	��Z�;���N��+�zAߓ�^��Ĵ0z/��t:x[
�!q=G��r8��� ��"b�WZ��v@�bdI��#\��I�B$MqSD��ɵq�|6\*�p��0D��ꀁBߝX�p�I�<xd�Cօ���bD��)س��8���Fll2/Y���{��ʠN�tb%d�+�.��� ԫ�(dU/)z�liU������xSQ��\���V0�$���.���*r/^��1c0���r_�|��GFZ:r�������'rs�u�XU$�En�2���gd�ր�Z�/sB�^>��q��kݒ���|�XL�"-�L62�J�N��B��J��=rzN���sn��aMձ�!�JVZؤ��	b���ь/�Ԥ��z�^�<E��!�@��ڜ�:��+$�xߪ�|peĕ<U�$��*Y���$D�{<b�L���؅-ͧ���9��~�`7H{�7a	3��t��4z$Ԫ��_~���~z���ԹYO	�>^PoCg0B�7����A���(�2E��v�H�l���vC�*��Q�Ê�p-n����B���tyqw��[/_|�5g�w��}���>�׮��Dh��u�}U������CQ�_򸊫���dv����?s��@m$j}h�
��eCA~.F�z'N�ɓ��`��xY�^c�Y�3�^-̉�� �)j��e��'CY��A�������C�`����?�ZV^��q���0���:UM�B]�I{�d���g�דϱ]�Ke9��)9LI�`(A�~/U�@e?].&�M���J6�H��
�"���W�喂���Uv:�#'_:��\|�~��l6��������S: �th5���C��t�x�B��Ά�8|�y'�j-��>1�/V-��t��ѣa�i���F�ƾ����d|�� v�,@�W��Z���}�"��D���!O<�ʇ����x���9��wz�xѱ	X��L����v�ߧ7���#�~b�E���?�j�j�ߋ�t��}�^��">;�7��P��H����8{���|��pb���@���!<?�;�GNBmN@�ZɿL38������2�m��/����s���a�֊
k�'S_a@�"�CM�`I)�wp�-�q(Յ��%��6�zs	zR�.��I ��:	���'�c��rAQ��.+M�/��� �h�Inv�H���F����m��c��@2��Y���n<�Ä�_�7� �_�����p��۰����~Wg�A��4|��tN�3�Yp���p�B6�-^���g��(v�Y�s��+@�ޏU+f�N�($%D���<�Ϝki�+����u덄�ZX����w������W�T�?�Q������A��[ToU\���������'�5�p�+�'���ñd�Bl��=���d6C�V-q����S4�g�b̤��X�D����S_�33==�^��!��_k�g`���Mg���¢�h��_{�iD�E��
�Ka[��[q�l+�ru�vY�K�La�^���It&�����!+wzMY��}�
	��g�}P��7�j�2D�PSv��b#�������(:��y��H� �*tJ����S��Dxt�#~�q *���?]����	�z    IDATj�G!�V-�6�UL�4	���*�v�bL�`&�}�G������p�����aj,[��-@Rble�x���Ѧu3�۰��o��Ï#6>6l�No�M7ߎ��B��Dl!@�׿���=�?t�~����a@��d��6l>z�}�9{3?���-��[oA�Z�а�58u� ��b����<���2c��^�u� �_��W�+�*�+��c;M���M�~**.�]��X�2tW��Cgz\	��WD����e�|GY�K��F`��k���T8����e����hYM�6�3.A�: �6ȃ�^����N��˛�|=*J9� �o��'!�7:�<n����++�`�B�U��	�$��^�����Dx�Fl�w���ZZ��fa��G`1 ���ѼE3�۷=�0ޘ<�r�f�F�:�#�9W/��I�`�1�[TN�h����<���l�ٹ%�'ѪEdgb��?�O�Gп��[��,���~1HGz���/Z#�H��'��n�{�O>�ϐ��J��c�k�!���)wr\8{#F���?��=ۙro׾%����V�щuq���~���hڨ��w�?ӫujjVͽ"5��C�^�?U���R^Q�t�h�4�1t1��πN�(]���s�ֳ�)[R���+Imj5��I@����TZƂ_��%8˛_p�^����b�n��+g�����Ň y9�[����r��,���-����4��yC&Q/b�8\^LF��0FK8J>8���ki)~X���F��ii2h����ѻo_�Tرh�'xg��,��G? Z���\6��X�Nd�GJB\�"t��	6[1�6/N�:����`�'�"<*=z�Fǎ+Y:�y��H�|����W�_��P(R�|j�;��(b؋�'���}Ό��u�/X�t� ��Q+�.V�����a��DsTa񨝔�����ul�$���+��}���u�ͿmϦ-��1�������Oy�+t��	йbU�\�_��Y��do[
�(�F���W�R'�kmQ z��~��T��-'�)!6r�!�^��$��kH%�t��]�FG�C .� ����K���#��rU=GO*|>g5
Jʘ���V���X������ZT�M?~�����SRРA}L�6cƽ��?����bL~�=,�z=���ч��v"J���B.>+L:+�gԅ��V�Dl�Ǐ�Vƴm�Cl\>�l5ⓒ��^h׮]�����۾V�}�?b<��?c�(*|��֑;ą�ǎ���ձ/W��R�$�g�~��8w��{�N7�ˆ>2����ư��ڷhq�?{��W������U�̿q�ȇ>kͮ�9�9q$����s�2��墡+~uэFV���t	䲚cnA]�>�|yU����~7�'�f�-N.d�\�b�}���5�A6�Ԧ������b��B��kȅ y��MVV���/�S�Ղ�}�</>U湅��f�����C�̓���C�7�VQ�����>�n�Ը�X�.7�
�`������qo"�gF��	�%��|(VV�E��!2B��C��(�,f|��

�q��)t����S���M��x��c��̬e+��V��?n��
:��r�Ο]��D�'�9�)S���W���o{�h��5����D�q��h֬#|3r�v<=��ͳ�q�:{�5ྶ�C�f���׀�>e޼��߳��rŭ�>�����b5g��T���2���FiP��"�s�%�U�kKE:�muRV�r A�^KV�<���(�<����d�x��|&�o�/��W���L���R�L�R^�����}����δ�Qh�_� �^��tk&�0��z3~�{� �����hݸ,JQ	v���0�ˋ�����C���j���`W�֪8�PjE��p\Ӻ>ڷMG�zc��wqp�F�5LEaav�ڃ>�ABb-,�xRS�k��\��c�׃����5�k�_;�`�|S�lH�}ΥДD����a�D:7r�.�X�*�wc��ȼ&��q;�Jm���q��{&9G��vb��)/<խ}�F�
��v��Zo�������ʹE�2�ݽ���4��_���"Lg�y��v%tE�%��M� �+H������7݄<���/�겲��� �@q�\������Nۈ�"���g/�ݤ
]��%8�^���%K�\��J���j|�\T_����
�lm#Cs����' �qq+��氳��-w^��c�;�����W�89rΈ�\1�%
�k�^�"�"�(�� DQQ	J�9���LOO窮���k�8����SԮ�o`��Nթ�^g��Z���e@w��>v�Y�䒥�=����hݬku��+��i>t�]�	s�~�={a��C���#d�� �r7+��I��{��ѧGw�ز�V-B׮q`�1��{ }�=���lܰ�.7y�ɟtV��֎���xӝV_Ċ!����A_��L��骀N,���z��v�ڂş��7��W涵��Zܶ�d��P�z�{�{�G��7���mk�O�>u��y��	K�������P�[����(�Z�X�F�b�E����E4���x���v-"^�"U-��HD�z��z�[D��K��SD��A[d�¢z��{�9r��U�&q��B|^��N���%��,G�J��t:9��ؓ&�A��a�7Z"X�m��݀��N��+�Z����E���S�<������[o�]wu����s�Wlȯ�"�,Ģ/(A�[|�p�����zCQHY��y���[X��X�v#�R�p˭w�}��?ʸ��)���_�EFH,iP���E��4Аy������!C����q����O�����Te֭�{l*���8W�!2�X�{Fx�W�F����������p�~Y_����&-��|��G֗9IK?��_� i���il���UD�J�N�'�r�
F���E�[oP�Y[�c.���xE˔���v0�j+�b�&�o"�->+������U'؉}�
�d��Ы���1k�j*Td�ĢF�SV����	��*%�INI���\^XLj:�/QI��~�~�6H��R�-�=m2��<��?���#�DD�	���+V��1Sq(��n��F*2r`��С��p�f+d_	���>.^<�����bG���b��Ν{`��B��{�]�+t#�S�aU���	��{sK�b�Rݻ��� /Z-����o`İ�q��I̚>	����ذAS��y0Frۚ5����JN�7f��w��e���z��7��5��GH�>}Ł���I˦����^�>D���\NN���}�PtN�N��x� ���!}Y����zU���W���q�"J�ߔ	`,�+"x�rQ� j�W�-+�~�+���bדp�p|��zU?���qȋ�JeeeU�o4 �NQ8B��**�cw6kDN\���|'Hq>:*��"���z���<Я/"�����гgOXLV�\��<�(��`*��g�A��x��e�"ޢC�n�ЯϝhZ�!�K21�Ñ(+˅�̃¢R���{b*6n��Jq�﹏IqT��Q�TX)�7?W��q�� y�!�%#�����r�>�A�1)���fϘ���R��n�+����DN�?��k(�PТQ���<�D�m��/]����a@��^�j�E�,��?�!+7'q���1z�+�<�vE=�T�]RQ��oj阘�Jt��\ >�0�����5�XAQ��5WgW���."��M�#��"�.�����"�)|U�M��Szu������E,PDJ�z/�H�Ӿ	�)B�H�)
�6�N�/Kj?��wP��'3a�F������;�=����Q+=e奰G�'�*kӲ<.z��?JQ(�BPt!=^ؼ~��3�����@'+(�=��~�Ԥ(de��+	�X�QX��$$&�WϾh��
���y|-�	������1��S٥�� ���h��7Bmk�.j��c����8v�,�?W�o�k;^�:��M�άgON�KCG��lR��9�͗�4��C���]����~�3V�ِ����r���}$,�q���6u-Z���ip�Mix�N��
v��dEd+R�"2'*"E0\E:����
���~wQ� L��/�t*�4�E�^�ht���U�₍,X�t޴����kn���M�N7�=�z���h��5:kw�_���vc�׋�H��eճd,1�5#��)w����%�0j�l�q����aAaf�^	Z��t���=	�ع�{|4{n��	��fa��}x��ǡ��g�A��{��h}E�*�~0a@��;��z��^%>
m�G��O"���i��`��]L��� ���l�($%5�>t�9u&����r�7��Gz���.͵�G	��xU~�c3wn�k�m()u$~?w<�y�yx�=0�(
w1�K0�	�(:�n04A�# �/"�.k��EE� ,R��N�%"u�":&�2���S=y��Lm]������Qە��aTb�+S�� �48[���l"��9Ku�����x���c�*�-Eb��cdd$\�
j>��� >:�K����ǁ�9j�p�a�W���?�"P��UW_�-����W`�w�q��cԻ#��X�,�:�v���F��Yb�9E@��c�`�QVZ��[w�o���oW~�ظ���>�n����%@�k.��nOۏJ�{�~���%�B��@�4m-gQE��#��E�>�UL�4	�woe�Ԅ�(�l�!�e�!X��X�T֠B6�^z��<{w�m�w�����Ow�~�O����ԕ�7�'~7g�~�9�"�4t�ʉK�ã���D[���LD�y��ω�Б)��%d�o����^?$Y�DnhT�7@�s���l4r�vQ$�c�F��l2��z�>,6|� s�,�)��'�?,f�O�ޔ� �V�ԅ��G�:��J�VT�ynH��g*U�n/�|rr*��J�b�#��.�SI�#���f\r��� 3*ʋ���Ux�gwn_KM����c�� kD$�?֟U>��s�7	�2ra�GB	a#%;) ]��wH���Nt�zΜ8Ƌ�Ob!��t���3�����>��M	ԕͭX�	�������3PEH��V	*��@���<��������#�0�]��:�$'�Y�6��e�F'ë3A�!-7�5v�K=��M�������s��n��	Ч�ش)�� q�����0��n�	S�C�1"���E5d��	�(2'`usQ�}�>���)��!��)�˩�ʐ7��0[���$�t�(����h�tCSxa ���F�F�#���d�A��1�J�	p��ˌtWE9�f���,���)�$��	��E' ���X��&���j&"�����Ҳ�>u;3���π���]Q��}�G�܃H�>o)�.��lF�>}0a�46T?a:>�49^��C/z"�0BB�v-�L��k��}۰�d_<�����G�� )��]��������ѬY>'�v�r
���ʔȯ���o�=f�T��Bz-䐖���|Ⱥpo��:&M��u�W����e����HM���FP��'Nb��y��i��{�|�g��{\�?�>��n��'���ɬ5;7�%-�p�]�zUJ���sW�N��Ѹ`�U6�f��R����H�E�{Q�Oѹ�OUk����
�#��	|B:d�۫��b�|倪�N�D�����[̰F��O�G�~Y�0��/t!r\3�g�	&�^���CJ2 ��\i)��T��T$@;��q?���%(��h�YPRV���\.KX�Q�M0Z�0G�c�����G~n>�CnkO�f��)�������kq����܋�L��1b�UX�� �F+�����a�Q��<���Z��ρ/?����"�a箽��߃���Ǫ�k��Vw��ŀN��~}­k��Q�}�L�� 5��F� ��L����!;�&M��۠e�&�rK7�$ԃ���V�5���C�Fw�y�>m���Y~����[��<���|�����TXZ��d�����P(>	N'���6.Z�跈�E�-z�#](�����Z5��t��R�5N�u�\�h��:��&"�Z��$!��py��Z�DDEA*ʝp��"**!m&}QF�V#Ar���t)�,HMK���o�AYBI~!|�Rba�k@�sO@B�7 )��6^8Xmv�l,C`��M��T�V�;]U�#@��4
H��<��(h�F8=�y%\ȯ@P�Cyy�o\�޷����3gLF�֭Q�p�G���������s��� ���U�@��F� Ϊ�S���ӏ�I�@iq&Ο���d��c��-x�������_.���}�-Z��F���^����~�~�5DH%C�2-�*#t�~�ee���A���ѽ���i��]+�o����-2�)u�������|4�_o��7�սE�z�����;�S�@�������ؙ��Z�cK~qa��Gb������STL_$��~o�
G�L�.��X$8#Hr�U`E����j�U��z=�����e��0�4HK��AZ$��EG�#����f��B�kѰqSD�#�.w���S�XL��ѧ�-0�%�|D�&`٪���pK:4j�V��]�Ν:��$!�T�g��P$'���#��y�d�88+�����x��[�6>��'q�O�/����>���AEG�L:+,�N�{6�;�ՆPȏk�h�]k�C�8��=���6p�=H�UC�G�Ӈ����tV.�q	�EŢ�����N��v�v�M��/W 7��u�����b��=���v�׭��_.C\|��� Z�l���-ς��C�*��.����^��C^N���|�voƢ�seŭ7߄��Rl�~Q�u`��A�ӏOM���3�_���خi�?�������r�
�1���I�Y�wl-,-J�f�(��`$./G��~)PE:Lo�>��]^^�J�rz�ƀN��t-j�Ec�� Z,�vzoVVV�*��]�׉)��F�FqX��st��65����Ӱ%ă<Ү��jhe��E8{��=��mX��K�_�1�Sbp}�����>8}��lF�+�r?8)�9p �χ�h�lZ����8v�0����?[w���Ebr:"#��"��$��:������/F�b⑗�#3��z�Y�j`�Y�G.�-i���:�&��A����dFBR
J�m-��7��>"[�V+t�*-�͠�A�#�,��.@�@�ۯG����I2��7��u6Ʒ�W#!1}����V���@�A Ls�����{��ՆH�5�:�:T@ '+Ç����o�v,�f!�I)��{�ixa���@�D�MǮ�9n�W���Y�NtYM�Sxܚ��0����_��������5;�;JS(�>��w�,.�Z����Q��0J��`��::�� U����T��p��<�N5�����*�v�-77�����qA���f�ghUǄӨW�v�;�������"���\��?u!EB|j$��Z��3�Q�Hk� �o�sH��e�6�SJ��=0����i�e����Z�=�<�<6n��ي��ڈ���
!>>Ae�+�&G���	����GY�a�Y�W|,�K�^of@?�����.l��4��+)�A�Dz��_����!�~�rt"��..�����F�^A����/��9٧Q^���;�2)��_Ｃ;��>[�b����OV��TE<�E�!�~In��� b�n~ t�������@����yÆ��7���wc���hҰb##P�A�m��ne� f�%��(�MM�>�g��k��ۍu1��_|&�q�i+vn-()J]:et�S��_�F�Ή�N��h#�V�����2��}��!�R$�H� `I�nUɊ��χ��`PQ�����xﭗ�p�k��S���c��P���a�F&ë�h�:9ĩ��NA	��d��Y�n�|�hZ�7����p���>W^s%4z��z>    IDAT��V
"�
L�*�̘3}.^|e0^~k�9�,���$�A��zLl��z��o��k�z����7��&"�^ˀn$�͑��h�N7��;Q�kGyQ!�� B~^z�i��Ƣy��<ǯ����$-d���d�,6(n�r�����O?B����]�ZBX0o:r2Σ�܉��۝=P�qS,�t1�C�<�mk�W��!������_�6��2X�0F�[6	�5:=d��� �b���&�>.��gf�Q�4�k��[��z|���o�����2Q'%i�跞�}m��G^��z�a@��/��sp��}V���۶e䥮�>S�}Ia�T��ÀN�B�E�-ұ}�HN�����uy�؅9�4m��b-$��2��}�����ш��"/��������];݆��J��[���ç����z���#��E@���Ǫo���mlzҸU���i�Z i�����0��Pd�7oB���'˗NFl�ΜG��o��O����\C�G�2�'$&�"�"t5#��өN.���ΨJߺ*`4�]��PH�Hk���tZXb�a�1�C:�4F�=C_�&�j�Q���K�����q�7�Oaa!�����.��\,��\x�<���o9t:\s%�v3�/�oX������}*��٢b��K����>�(G�J�V5q�������{��3�SO�GD���!eh�G������_������#�3s"��p�7k�N��@g����)����G�!�f�9cě��7��C����/���������I��6��M{�:�i�r�6jJ�8�N=ܔ��v����	�	�	�i���6jA��,_��T���gh�� �ޓ��Se��p�"����c}�떶H��� ���ØY_C6F����Mz��
�q�t� �:/�{�h�8^g�*\�2m!J�Q��Ѿ�5�pJ�����9�0j=x��.hX?)��8w� �܀��r���T��%@���j�q�z���;��Lu��@�5�l4��r�+����i_f�0�p�l>�ee�p�8L��"I:ׁ#��W`ʔ)x���q��)�=�2.��}}o|��: �	I�`�hٷ���Y��p:�Q/Վ��hdd�`�����������/��#�=Q�r�0�_=}�j� BZ��e%-�~������˘0u2��)�M�O�8>k7�%6�΂3��(�H���=f���;�i�O�<.�%?�0�_�)��~0��z����ZXZ��Մ������:w��IO�J���Y���(Z��/t� W=2�\���:�&G2A*��Ɏ"xw�H��!.B�����K��Љggr](�*�z\ױ#�=���;E	@k
�i�4�D�x�WT�ܢ
����ƊVTC�[��;�nA�@�HO�":BmH��'�J�)z� 95���z�Qo��#XVTӂ#wz�QH��?x|nx$��b�T��m&9}8��DD\<J����x��c7��)��z��͝�	�зo_Ȓ��C��a�-9��y(�)ĺ�kp��Q��>�}cL4=����p_�gg0)�������Dlڸ��������>��c���z'�S���TG�/_�G�r���	��<����?d@���0h�����5���cD�
�h4�Ww����;�VS�27��E��a��yug�ڽ5�0?�X�K��A��,&yQm�X��5M����Ye���^��p:�7��^�8Z �����.�*���EEŰ�m�i��d��u �q���#�1�"�E�ƍa2!y|(�/ 42�V=l-t: HZ�0��<�%z�V������b���D����#'+fK۞ju&d�ѱ��F��p�	�e����w  s�N�qt>Ծ���P�(�s�������12g�P�zd���o���}��U�����~m۴��bƝwޅ��xu�߰=~�o������9܍д~�Kгǝ�.�Ņ'Тavl�茐� �{�%��b��}pVxЛ7o��2©3��������.�#uLH~d�;π��عk̟���	q�ԩ+m���ؾ����d@O���>��7����K�{W��r���Иٟ֙�z��2Wy���`���Q�WȪh���Z��T� N*����"O`���]����W����)��O0�H��rj^%��a��H
F�	f{r��e��_3E�+�4Ğ�@R|)�)�$mv��i*܀-"Ί
�m5M������\�.hu������hɺ��e�p8UG,
�����o�e��9�F����(s����	:�{�π�3@��0}�<����Bh޼>�>'Jʊ�V���
�����f��'���_z#����/b��X�h!�N��u+�E�:�К(/�×��Y\ �ۇ�k���G|r*��>�3g/��$,��Z���������#tJ�O�9�����!�4���xԭ��x:[$�O���:�zi��f����m6,��/|�~�O����K>���k�Z��X�>o�8
K��R���@�Nx���\��	;UA���>���wѯN���VU|N�xU�u-�0��ϋ6T1YT��VZ�r=�$2e	V�f���!҉�K��f����n�9f8�:ؾ4�h� J�J���^7�����	�
��Z�|���t�����R�����h6���,��#�VzhZ������
�LV@�bŒ�1m�8��D[p���m؀翸ȁ&M������9���Y�L�.	�$#!6�O���M�`��	z`1q��n�f���3g�f���Տ���
K0�ͷXX���8�^ٺv�o����c�+!����!�b�q�'�R���ѹ�5�Mп��D�2�{CZ;�Iq�q1��?��]:�*O��s�7��S�~Vkښm�2r�j}9n�}2�*�.�⸷���T�НN'G�������~�"���	�q:2^�~t�~��oA�#��A�֫��R�z���$pYS^����J����g��T����!Lo���(��� ���j��kz�No}�R��B�}�
i�]��O%�O�g�X*���-��)����xVX\����(f���
;���ь���ѣ�m8�g;Z4����
�b�`�F����_�5�v!`�#&!�N��.X�zvik���7^	��\�e"��a�J�綵%K�e-w"�}���,&���/WS��A~���Yj��� =��*�����{#p��n̙=	7tꀮ7݈]�!"�6��@�_��Ukp"��	G�|�֎�څ��j����a@����$��?kV������;k:�-|��|;p�S�D�S]ш�f�Y���?&&F�&���W�|g�2��C���"UD��9��� ݉8��đ.��(:&Os�Q%$��j���v�� �$^pP�L�˖����*'f:��T�W��IT���D=�"�
��u۵$�A�ٴE���/#2*�[e�+�Nz�t��)�Z"�;Y��v���}���%��X�QvlQX�a�=K���m��e+DYM��<�̈́��h�8�a��@�:s$V��kZmh��;=�N������Ipg�f7��q��a��m�w��	���>�,v|��:�}2^}�ut�B�`O�V�A'e2:��V33 X$�]����k^V&�y����G�q�=)1j�B�-���l�;��#dO����{�ΰ�Z�\��a�0�_W�>�S�֚�q�ֲ���+gLƒ��bߎ휾&��Py��Ȣ�ˑ'1�	�9M��dj�M�k�BDC��E$N���u��w��FѮQG=ު�*����,գ=� �����v�f�r���������s{�G%��}ު�;�Gm+��A��Y��2l�*��7��HF��+���"�����+��)·X�88��$R3iU��(���%�;g\��pA�񂣴��7E�׋R���#'���c`�G��,���:EF�F��S��(�&=�B���9�.p!���z'5n��|�Éw��,wġ��@�p��-y���|�w��3@j�� 1%H$5���B���@>�wl¢����v !2m[����(��� 0F#%!z���_�um۰����~����s�}æmY����?�V���͛$�5���B��@[ 7TYY���Cit"�	���@O�c�2�~�H^��п���@���hL�V�U��AqIby\J�GXmPB�j�j2� �)�NNh:�J�#���J��h�����%�������8Z��3������` ��),$�`��A�T�'�w���h)�O /#�nCv�g�=@Oa�_��?� �
��v��KZ�!�/�6 K�m��Bb�k��(�F%�(����܉�����4�:qK�/���ǡ(!�;���=� !>��Z��AC���f͚U:/��笆X������v�DI�Z!R�g~HQn���1���_��(n�tn����d���7��B��k�m�����xu����ey����
�?�5>¤Yҧ�Y�=�����qc�m�R���i���ZW% %Pus��E��Hn��\0�YN �`��>��x�_WJ���:פI^�T�t:O���Ft���.����Nrt����Ո�"��z<��d�қ��(/wTF�Z�D�^x*'���b�G�)&,&kUƂ�EoвY��@Y��-V	�k�JG���
/�Ng�F�$(�!_(��l�� ���z����B����+�@RT4RRR0��7q��Q�1tVl܆CY�0E��窀��M�1������ְXM(/��'󧰶=-2�l݉;�u�5"k�mD^~!�5M�5��>��
���׋:­�5����(�%Z��F��Qav6�~C�z'OŜ��ѶMt�r+Z5o����(q�0'$��3�d�v������=�mk5v9k|�0���%��`ܴ�is���^ꬨ�d�,�d.vo�3���p'P&���iv�?h��isU��j�ԓ�Q�.Τ:��:�
��_A��}�S�b2s���,��n��X� V�Q�v�V��,����S�ܪ�����왧ł��F�R]����nR�}�&����Tӧ4�ڲ��sTk��-dbc���^�qqq�i5�z�י b�ktL�#�/CD6� �M���/��GBBLײ�c�����ګ(s�c��͘8e*6�9�o6�CdB���p��Ѕd�!�A�cG�ň���̉#qk��زu9���܎��TtZ����+hڼg(�A�v��(6��{x��i�PC4$� �/
��0x������ν��G�^w )*'��F�>�¯��\�-^�Y%����;i��=�)���5>p�k���0���Rg�ܴ3����cFs�N��#�:E�������ggg��z��q�Z�	l�f;�i���*�]�DU�E�p" b��)�P���r��yj#?q���r�lF-=���|D��n��	��c�=2.��A���@�dZ|~��l�(-�٨��jf`B�J%�Փ�f�<WS��{��̆*=¡yr8ʑ������iC������4_�مe�,A�t�`�ү8�i5����ے���s����/�ơ�G����X�u?],ETb-������2�r��*�ݰ�l(*����BN�9DFD��oW���BrR��f9�~CA�&͙�_}�8�0������ ]G�N�I��%EB^F�O��C�ٷ�fMB��uqC���*�`���H���Ɇ�R`OD\����a��ݹU���;���59a@��ٿDc���r��bGy�GÇ���رi#����Q� �"eJ1Ʒ`xWW�c��S�+���.�sJ�ӾH�R�QQ^έf���#l{d,���2�L���)j�=(�`҇Դ�^g���U(=O M�p:~"ӑMkH������Jw9R�sy|0��(-u@�'g5U����hLe9��U���$4��N:n2�	jX܆#t����q"�!�e��f�2��³�p�~<��;�FBr�L���m�K���m{��hV��H��$�;��lF�(�������uq�q��~8�.�#�qW��hP�1�._����{�7��Ss/�*#�0�_��g�	�d.3}A�� �	�Fa@��0{�,:�̓pB')�pյ��4 "���!���L���a-����5=r�k�
\��'��,u�����>:E�k��k�0������`�S
� ��M�����j�]��B)mՉL�ګ��ɍ�C�+�~2.�GE��G��ud�Q���֠��+�`�"MV4o���̭qy9Y���hҨ1�L������֓fk���+"��8����y�����㢱a�w(.�c�'�6ۣ���.p�<l3JlcZЂ�T�h��dd�t=��DǢ����YV$DE�Bb�9U�f2"*!���KD4��x����3�*кy3ȒEE�� �FD�^�ǟ,�K�`�LX����^RT )�y���hݢ!4z�?~?��{��b@w�}���;�V�.�o؂�F����7m�}��3(a2�%x���!�E�.��V���{�"��2f̘����3&0)�_����z��k� �nS8{�M��|������<���7_�6�:������/xQzJ�g|������/de���h.ϙ��{� ���P�l�2U�=��W�(�T����X����Y���eg2�����ϝ�N���"(�v�JX-�R�� ))	3f���)Sٟ��N�X��aŦ�P$=-˾��Y�a�r��$co���� :\{+�p9tNG��N��U�p��Q^<hu:�'�B�N7����n�������js-]�)wJ���]PR8�N$8����<z����H�j�[H
 ��g
<(شtJ ���A�z�k�۝�s���k?�1A%�cT"\�XDŧ�2XyI!,=��m��#}0y�H|��صs=Nކ�H+�^�_���1D�%�o�#2*��V��t8*�</�:U�>���hCL���Y'���"��x�Uv⻐q�&��bD���M�@�F���k ��=u�D[��f�x�G8B���Y�����~3>�*e܊U��k�|s0
N÷_�D0B%ӛ�q�Q�]��'''37�S�NUi�S�n�[�z̅����W�[d:��'�_����lټQ�&�H�y7aͺx󭡰ڣq��1�Z�_��#�Maт�(-Ƞ2;���m�k��̀~�wB��?�o/
��P�N:6�����AO-f
4j���q��]��Jց�sW�����(�N�:?j��l��CAP��/Sﰖ�ZRH%B�=V�<�)w��2g�:�Vj
�>�?]�Vm�`ʴ�о�T�D�i���}^�fì� ڤE�h=4�Ǝ�pb�GSѮus?y
�6lēO<I��?
�������4��s��r�E&F��2��f����C�$��H�ɀSG�`�ȑ=r�ރgM�-];�VR
⒑��щ�a�O��／GΡ~���^~�{��5���5<p�i��p)����%k���<u��}�[֭�v%���ALU���X�*�~�%��R��v��I~��)B����f��U?+LLպ��D'Z���}�V���U��;�AC2���-�����ɧ�FL\n���eL&|��b~_��M���yp�@	XS�n�&�~9�����B/t�Ǐ�����W,�
�Ng@'Q���zܻ}��y���u��g����y"�Q-��uh��em��"� �(�Nj_:�Yu�SHJ������`��J��"���''!&.=z��_���зa��C���t�̉ḧ0�q���t@�-G�]����iצ)��M0�d��c��x��g�L���\S'�����a�[�TJ�Z����c�����h��W�F@��F����q�`|0�}d�^����ЪeC�����7Kףn��p�@����6t`ƈ�m8��w���7��ݟ2�    IDAT\C_�v��������q��P� �SUN ��.�_�Ujm�ni�v���`�>��*FW�RU�5B� ]�00V��W�X9����WU�#
EAQ���܃��D�r�,�b4����/y�ѲE3̛5�Y��F���7�U:B��q�]wW�՝={�A�E�F�f�"d_<�&��q�-
O������7ue�T�A��,&�՚?��+���S	�5J�	{�0���-jt|Vr[�Fbϙ|��!9V��c�֍�km7����o0�<\��z��������P2�X�!�f2��(��D�UMy.�J�]�]����8}������{�j�ĩ��PV�°!����e>~E����	a�{�}�S���2{
��t�?yo|�&M¶]�1}�$��a�Ьi+|�dK�Z��%���4�JI�9��z]߾}�>��.k�����K38��u����x�pdُ/|#��p�X� *��X>է��&@��N�8&��t��;1��@��6�S�)�#f�uz?m�V,�����ka4�E�z�����nꂴZ����mӂcْo��xe�v�9c*J�	)�i^�n]t��3����X��;���ً+۵��?F���@H��ߠ	���sX�n=:u�����j���Sp��� ��
z�͊@P���L�ɪ�<zHoƎ�����a��U�������Cs�Έ���������l}g6�:�=�
У-&��!P^�Y��:��KO=΋��<zb��39C�����2`�ν��<�M$&���3��
_;*T��.�M�̀ t�@p���+{@��'Or�}�ȑؽ~�1��V�}z��)���Ł��h��ȫ�vr�ι�Ѫ~������~����??m���W� =��,�hLt�2�nB&Ux�S$N1�����H�](��MVDDG��Q�����2� ]��Eݖ ���b�7�zʱe�z�F��\�� ��;u�������.^��n�Rt��cǌ����{�5:���G�>(*)�m�w�z���38t� ���̘6/��Ť��'��a�!X�v���:�c7�̐d����bFe�1����	i!�u;�7�����M��zP�a|�� �_&�,Ŵɣ1����./�3O=�V͛q��nÖ;1m�t2��ea��,�bS�ҋ��0-3�C��D�=�߁�� �W�_���[Ы�}hw�՘>{��_|�5^Q�>1�%Y%�_�9!:���Cp�":�
r'H�|tR�;�ofM�����������L�h�m�4G�+�F���P��q�>y�,�n3j''�>�a����b_�C
�%��� }�-�.w��?xǶobR���E�L)r}S�"!	+�]	tE*����&52'�ur��P�"3?h���2�[��א$7��
�ˍzr)}M�`O>�����ՓA��vlGaa>�v�'�%Ejk]�GE�wG���w��~��N���=�йs'����8z�0�3oTT4�.Y��[����7�J&'�2�F)Q�\P����P����lM�n��&��-/�#�^C,�t��⃮2|8a��*ʊ@�CB��:`��}x���L��(�ݹ_�������[a6���CJ|�ʤ���7�G��X��v�jt��f���^̞;����y��@o�@�F4A5�N�t����z8	�)�NϚF��5��-[0o�2�k��{7u��6����nŅ�RD$�a΢����YD�{g��r�vM���Sk����a@��+p	Ɵ6���	+���p��,xo.܃�_~����W˼�<fh�yWAjf-BA��sZ�#�p�2��z!TC�gkS6P�A>vْ��x�3{:6�[�R��Y�Y��O�����.�܂��2>��;w 77}���e�E�L�3�������G��}�$fO�8�����W���SG�<y�!���n��,]���މ����%�dU�\�{�|>���5"4�\N��WAg��3/n�r�h���Y�GD������.�c������SкeS:{����Y����Ͼ��N`���u64�9q���Ï�(=n��	�YYȾx��7@�fPTX���v���7�;�c��i0[�x���HM��z���\�N���_/���PT�^&_ ��A�qw���Y�1꽑(sa��ב^;���͛�##�	��Vt�s�, h@����7mPo�;�=�#�r��kZ�#�����%�X�S�n؞[XXg��W�s�aδa�X�lF�؇�ku�&�7��N�I ä8�ۍ���RT����:M�����X��#��/�#::�%`�R ���?q2̖t��3��X��;dd\��?�F��(e7R���m;v���㸻{OU��b���ؾO?�͛5Av�E>�~u�<HI��ѣ�ছoA|BA���U�?���/R��|/ ^)�z*����6����rs�M�~�قF-Zc�����������YR �<�ЃHIM@qq!Gc��x��*v㛍��
�F5�,���A/b,2��2�'��.E��Q�w��i���qM�Nx������G믶�i�[O b�S������K���!�f��{I!�B~���;ƀN��{��0� �N��u㫥k������`�L�d�BRL��٣_�����%���À^��i������+�ߞSPPg��7ql�&l۴f�����S�{�nDGG1��"���V�����mC5����Q�&m�wo�Ͽ�s��{+S���6��FEEa��i�k�X��2̞9Q��A?�S�&L��`H����zxѰe�f��f�чB����r: �0Y�l�Bl��{�������gegb��%0�4�_Ξa�P"��Ux��1���pw�ް�#95M��ܜ>J�	�� d?��5ݓ������hݖ������j-}�	�����
�^���)q�(*-FI�I	q�*�ko茷��Ć�9��"��������@jGkpU�FhҨ)�%��=���N���	�hղ={�|0v�ԯ���!%�64Z@�^A�\H,}&ʑ%G@\�_sW���;q&����(��M[�������Ou#���Y��W}~�O����s�Ӛ��"�U`�j��.,�d������%
�����N]��ި%�����7z|L�у�ug端k��҅�����腭~Z�r_�z{��Y��1c���j�2fJ�v:��Į]����Dfz�&9Y��lGJ_B�f�h�f��F*l�j���
E��wѲ���ɸ%�F�Zܞ
��⯾������_���!>!�Ǡ�7i܌AIo��G�ޜ.��z��u(*.���?�v�ڢ����g��[�;���O������kZ��:q���F��=��~��qzG�e�^�=���oѪU+�����$�:�\p��,����o�6(�%�?����V�Y���<&,}�y'����i���{��Yú��E<�����ð��0}(*�G\r
Vlއ-ǊP��3$��fRl��wu�խ㚫:`�Uسs=��28�޵�u�|���3=�܃��Z�j,�A��u�PPmd繟 zu��E@�v��7�����~]j@��������- ����CAJ��bXG�C )X�N�#;�b��Y3~֬_����A�d��W͛�F����H���w�L���a5i�=�g���3~�8ï�5g�>O�Y����
�kv���:b<y����T��I���_B
��ك��xv��E%��b1f��&P�٦�Ѩ�͠��3N	r4O��S��]ڟ��SI#݊3'O��u�>���a�T���H���#,YZ�~}x�>x�>���z�Ma�1E�_�գ���|�����[RR���MZ�����H�MK`�pV�J�jדf�_e��Ε�	�zph=C֯����u;s?��+$���7��]P�iɋ1����飸��~x��GѨe+�uZ\ۺ9��֮�'_x�rdH�X(d�*�`�}��`���µW��RA�]�%��Dq�9�����[z!)�V~�
�o�v
��Cse�����΀BER�̲"#��m���H�r�# ���I�ߴ���z�M��Oq�?�� tr����t�S$Dz�ļ��{�a��q7y"�o\�%�~�����-�"11��4��0G����r�6D��f�?⮰}�o�#�������w?i�W��V��[PR���С(>wϝ���H�s��2��=55E^��=���j�yRdM���h��C6�*K�l��� ���$�Ϡ+ QBmU*_K�ݕLrY
p$�ѳÉ��h�%	T����j�{����U���鋞#y�PK��	y,���臅_�d<##�h��K=<9���B�9��U;����dY��������4t�ԣ�5�0n�B�-�����-+��7^�7�?èw��k��I�ֈ����E�v���/£����"h�C���>xOa.�?��
��II�8�gt��nR���X�j5���+0mؼm+n��V�n��I����:� t������_�,g
��������[#t2��-�/e0~n.���B���@��_a��_�C�Upr�!����;zr��1s�$%�`�s/`���U�C��m��e�AdU Ƣ?2y��ulf���k�g��o����g�7:���}Vk�Wkv��ޔ%��c��eX�rG�D��h:2:
[�nE��yf��F$5YQ�ZHj���e��f����� I�9��meݙ�WE�9�;�UҲL0�eURV��$�ٷ���5E
��<��ͩ����%D]`Vի+{�	��>�I��t�t�9���F6v��KKKa�?@��YR���8) ��΋�>��_7���������3gpE�kx��6#�ݕ�#�nc��YA�� ���}�tC���0'�W]��W�C~�9���K(p80~��X�/^�^��W�Pʝ�{�a�J��=���\�N�6C�Z������C���C� *&�6mD��;��uF\b
B��
q����������F����P�Տ ��&�߂:�|��� �'�7l���=柜�OFW��������V������q:�C+� ���c�3*:v�����`�"��t("* "*'8�k���}���׹�y��\���Q{�����}�����vN�y�k{�H@��m6㩑#1�՗��j&��\.}z�BKDÊ;�]p�Ϙ�>�?��ܽCN�۷�8%m�7>m��o|�~뮏�8�lԧ��jhii���/�y�n��]��	x9A|��W�ҭ�OA$��e;��רMM����|��#��G,�`����g6;�膁H8����mP'����n�;x{�L��^h�A��N��T����(���հ#_���ɞ׬�w: �Ty�Q���y;�y������nz��*�`�: �D����`��������**����1l޴g�ٓ�MőW�_}�#I��r�.t�TE̢����2,TWQ�����B�2��j5���deX�7"��mG�Àjf�I$QT��_��1c�G4f��s��=�w�/�i���>}�!7���p�f� @�����B����k7ܯ �����{�����~��I��~�X��c��=������[�qkz!-�haEeze�$$���u�1���ĳOcc��h�jQ,��g]���@�汿�)9 :ЕݓF�?�-m���5�w�����^۟�l��S;�8��ʚ��F��n�ˣ^`��Vorr+[�z5r�m-�%�޽;�9�8�DY�E,�{��$U��cb2g�4�Ku!� �x:���3��5�*?�,���)�ԩ��fR��4S��9���4$
d8�1�S���TuR��t�4�l�I�cܺo����*��i�@�Nb���dbc/RH���0H�vKKK� h�ۋ�@,�~�-�/_�G��s�nt�݊7t޶��p�Q�����×[�P}=ƍy[�Y����� �H"��g���⮺�ZL��_��	�D:�.7�pF2
!�	Y��[��C�`Ѣi���E*���}�GYY,X� \t1��w4rra�t�l�;�L;5�P���uh�&�W�"���_��#��o�_��M��;�NķVP線l�m��ϱ̿l),d����U�1v��x��g�����⹼��(>t?b >�x	do>$⸨.��9��ؽ'�<�g���!�\��Cl�C�¿9yv���,�vX��{X4�#�X���A�,����&�U�ٱ$�w��z�:�4�����:lذ����E�0}! T�*�B,��А�=�������M M�z�
�Z& Z�&�YśL��V$U0�N���Dr#���p!k�?e�[ݴ��;�D�x�@/2y��UL{q�Nqg�����y�M�{�?���HfYp(��g͚eW�Z�'�|*�.��J�4D���{̉���W�h������F�����
�p�#�����v֣?��sغ�����@�¦&x9i�m�!B��=^�?|-f�z�9��X���X�=A,��k�{�yx�q��-�����se�	rF�&����7U���}p������������ڷ�8�׀�o��~��b�/�G��ph��~��Vr1܉�B�$�da��x�	>�ql��f6�y�$\{���' WDU\����jU���C�O��c�?~F�>��|� ������}5������Z�&;Ž=�M8ԟ]�HN@U]Sǀ�H�p�עW�^̭�g�-��5�Q% *(�C��q.�m!kZ�NlxjM��0-&�Ѭ��h��ry�L��5�6���*�t�g��ļ��:m�l\sssA@-+�"�씪�v T�j�5��Cu�l�B�I�B�"�ыg�T��:����y1CU:-4HOߥK���-�F�2��:�V��cΚ:o���G�б�]D���~���@&�'3����/C,܄�n��p��wvlۆiS�bѢE��?cgy|�	I��N>��d)IH@7R�>����sf�ǖ�^�=��G��ݰp�B\�(��>_��؀h4�5dsz��o��;�V�`�o~�)�\�ߴ(�����η�=�ϋ��>�����x�T�
��`d��~�&��}�1l/߅y_͇%�hj��ҡ���'��_ԑ=�%E�a�(p���=��O��&[��y����U��ϟ��7����.�X�|OEE�i�=D����#?/�[�,Cs��c���I1��O<�D����'@�9�i޾C)��$=̩�&}-�-�� Ϧ�n�S�m/������mrA`�-2�rL%3���f&��΋�@��e��.@V�t���s�-�����f�ی}�o"�i����j(�é�<��������,����hq�a���m"�N&�ѹr����tVC~^�m��J0�^U��3 S/��:�E��=}n�y�-��\�\�]x>v��Ì������K/�֝��c5L�I]�%��@0��efy��RҸq���f�b�^�p�[�^(�-Ŋ+��?\�3tt����GV,PC0	���/���; L��W��|�Y<���~u~;����m@�tJ�S�g-{<dd`e�ؾ�[n����U��9���0�g�;�ޒn�_���0�P��w�|��>{�w������>m��?}��l����v��ҕU���>�,ʷl��I����9������K������������/�%R�����՟��2۬��x�ގ�"6;�";i�utpj�Ӭ�@�@�gϦα�.b-��oZְ���bڱ�n��A8����u،v��әb�ڼ�U��G4��|>d�o���:�Z 45���g�-2���ق�8D�ˣP"��[�"	��vچ:��0�/����M��t
ޞ3������h�x�z
9>�r��{do����5h��q�E��1��WA�`�"dU
|IB�RM���!��^���e����z�w��9s���u�]�n�S�    IDAT�	Щ�$:�:����A��3߿�ҦE����o������߲�����ؠ�n��S�+8~�f=^y�E��vV�Ŕ��0��Jqí��s��W�"��|�8Q=���N2���m��:��@��|�;�;��d�ʖh��e��]�S&C���cSe����r�gN֪]�ve����^�r߽c'K�|� T���8���~E����453�2N�5�����^d.�Tl?x=K^��ӨZ����V��#�LrZmTj�S�:�C��oj��NkYTP��4�L�er�!әH4�3|	��(��ʻC�ܭ �!E 1�]��2�ݻv�1H���Ʉ�ew�z�?3�XQqC��1��	���?"�KY&���;���� I㖻��_F<���/ߌ4hF"��B'� R�L�e�%�q�%�i���pѓz�J�`ٲe8묳0p�q��r`����2�ߥ���:�*��_���ҹ�#fm.�='�$:�!���_�b�b���ݤ�V[֬���g@ߵf̛�? ��ǉ�^�?���ȦXupǫ�a֎q��C�ﵻ��g�������O:���puc(����KK�����1=�	ԉ`Fd7�?hϴ5�����Ќ� ��TWW���n�����U�y�L9�d�B��Xj��yA@��Ɩf�&I���2��ND"!���҂�dp��\��:Wܙ���f��/u�Śl@C��T�g�,J��H��,�#�u~nD�b`�����^uA�i�or%��$��Mr��?G��n�o޴�G=x$PX�����5�x8�G�G�@��0��]��Hǚ1��Q��`f"�;�������/AEu�ʛK��2-]�@�)�g�<�,���4l޴N�&q�Q��{ >�l��|�aH�pmC��1h>�ǳ֪�������
�������r���=����/[�6��ω��Ǌ�FM
����ͫ�`��W0|䣨j�Ƭ�3!�i��ǵ7݇�މ@QWXa�ڶ�����'�8������<�m{�Ϟ�6@�g�����͘��噟��onn��#� �P��y.��>��t
{��AN^?ZZ��m���oW��� GGlpbd��L���1"���h��f�suz�*�Td�Inó<���N��m����Fv�I��I�KD�t��c2�q(2W��X�� MmGͤD7�x�u��bG�i"�Q����Q[_y�����O�i�n���c��U�D�����A"���gr��3-r�t=n��L~�&2)G�Ϝ���d�X�Ȇ�#�v��/>���}��uM	\����B%����რ�$}�nJ�Q�$e`d�PD>o7�x֬�>��[*��uG��ݰ`�\������!�σaR���47�A�B�Z*�'@��g������_T��lU��'��?i��/���m�NL��^��y'���Z �_�L��·kV�Ï�ǽ߇��嘳p&��fF���������#'#Hr��z܈[N��I�f�����_�m���9��_���ٳۿ2��5�r�9j6-]�%�?窘f�Ty9gÆ�JzH����l��AEn=�������Cgdu��]���I�:�%u���������Y6��g]#KR���;y�9-����j�����-�H�s�v�gm���v�+�!��*|쎲���<R�;>$"!8�DRYT�����癴���K���|Ĩoe�/�tn���z�&���Rw�[���!cfl�}<���;�L��/jV��IB�����8�gO<5�$"5��Z��N�x�%�� ,g ������蜕 �)�c�,�iO*x<��mx��бC�"i��9�z��k���������R���%Hmp����~0���7~���.�(��!����?���g�7�ϕ�C���~	���v���٩i?����]����v��Z$�X�A�eJ��Nݠ��Vr���߈��*��t*�9Z��m�j2r�+��e����f��;��O9�o�l����֟l�����v��_���zMum]��c^��m���)"77A7A>�iJ��{xn�L2���:
���M@+��o˴��v��	C�`�N�@��K�w#�"Ǳ�e`�[�1j�(l۱��<D�	�T��+�D4����IgT�Μ=[�~HNH7�^?�2���Mr4+��EI��5�-���1����n��' M�xnn��H��p�5W㼳����61C���{0u�9H��p��d��]�>�tV�tPT�CǼy���X�����^���L��W �P�%Ņ�47�{����d5$�)�C�S�����4N>v �����r�b���x��H�2�:�����b�;y�ӌ�x
Ґ-��p�1\u������p�"���#���,��+x,�;�8th�	W z�g[��ׁ,d@?k��%��q���7���-)���.�}�~����̭l��+�V�{ �:��{(�k� [���B�qL���G��{~��_������/#��p?�
�Ց���v�^4�2<&`����(JģX��K̜5�]s95�is>��raOy��#��;L�ÀN�<G�V���]'���������� ��ε��G2~ƌ��3�il�����d<7�x��,�����솟6������ÝK g�drkKe��Ѐ�߬C�@F$���GR*��O�Ul~ ����x^�uע��	JQ	W�Ł\�"a$�t(��ݷ]���C$����y5u-��k���GV�ÒT��!��,��^�����|\�`a��}x�T�oj���C�� ���RУ���Å���O�Pųc�.���������!�18��*��?�yPANw18$�֮D]}���	�ˏX�D��Btz�Y:�N\�����������&�{���8�UxEg7W\|�F�Á���/��˯����5{��}6xRD-=��$iJA�,(䏟mƝם��?����<����w?�?�
��t`e���P�H%�:��2)�)����ߞ�t6"��Bq�����h_Z�j r�� �ܑ��R���]*wk�o@c��:��~�/>��;D��D?2ҍ,�浒�n���(m�d��C��`g?�ݭ�mJDX0H�g�wDI�{�#HI���Dv�^t�o����%du���O�'B����.-.9XH�g�8���?dck��1�aP�
).�p��Yg���G^NY�h�
ꖆ���!�J�&L�Īe+1g�L�p���f�.�������q���p�_FÛ[�����E6���kV��Н��l������b��~���_��ٚPK�d���X�r)�L�ɡB�-D[�aXD3��J��% ���{�[D<����F<�����}(��EC$���`��D2(zH�:2Z�L+�	�0Ϗ9Ӧ���/B](-��x.S��킠��RV�?]�p$ꫫЩ�=�8�<��(�_�5�ʁ��B��n'R-5�xp?��Ͻ��w|x�1X��lٱ��Bh�Y)�+��������b�7k�j����3�%K���[o��HF��W��םr�	����
<�����p���Pֱ��q+���~��_�D:�d��>x[��c>X �D"�����#�C�Sı����K/���}�R.��ձo��n@TW���������'�M�"A�d:�p��x莋���w�v˜5߫���Ю3|����	7��N����5Ȓ��be���� �w�Ѹ��wH���E�w�.6�!��hn!M���3�0����u�l$D#� &�����Y�@�d�K]���<�cI�w�yX�dK���p���Éw���J�@�>C2Hb�Ӌ�O���Y�II~HUj�V��&k���������uAE%�H^�a���2h���w&���<&cR\o�>}x�4�!wE�WRo�^�{��Q�"������pyx!&(����5<nv[�cb��zhV����q�-;a�u,�b9>�7��B�>�Nò�HDǣO�Ņ���WSU�+�%2(t����o=�������_;�6@?.��3>������[�%��~�5��g�cL�!�&�2z`	z�:v�H����>�'��3�e���uH���o����U7݂�."k��L�=?�t�3q�V
ss���a��Y�q�UX�a���ږ�t�
��4��0q���밎p�v�#������;��TH�bxr��P#тsO��������2�>{6�۲{���S����-�+�h��9Ca˪���[o�2�~۶m������-@��=ك��v^'r(�2`fR�,���a���1��x�I#Q_~)����`?�S�&|��<?�e�����F]���t:�|��P2iӽ��u8D�d��������ո��Q�żo�!#���H  ��=1��Cc[ڧz<x���|�$��N8d:w�N���bB��-s[���S���fhH��H'ȥ�O�ْ7�L�9�-�#7'Ǯ�@U���E\�fCt"�eY�GF@D,�ʘ:v������{_��0O���rNj	���?�ҹ�����Ug;�ٳ�H�����$����������'���������+@&C�Ĺ�cw(���`�!/j��Z��ڗ����x��me��L�ڷg�O�3vڠf?���Eu!�A�~FEB���Q����fB�=�-�`;$�c	(��v�z0��������҅��ı���ӣ&qG���y��z���o<��!��t��s��ы���wz��kC�o��Sŵ����)\�^&�Y"܄�{��I�3=�.]�`����6�X$��@eU5�KK���_#��C3E�p2���H�c��U�_��<Lz�m\z��'���J2�]>d"ax��U↫��c��� F���ߛ�P$���*͘H
^XT��R5ѫC }{t����dA3u4�B�:e&��"�WQO����0����{2�F>6j�Jb����:��C(�!�1�p�Q\\����@ia�����u��vXw<��s��b((*B4�cky-<yܪ�J~��I���t�[�$��U;���9��W �\��������F]K6~��w���ކ�HsW����V2�X&W�
�"p�6�؏;o8˾���� 􌎒�2?h0���=�L*���`�s&Mmh���6�Gt�el}M-���d��y�l�K�L�OcuQ��=`�K�r�0�H��ʗ��~���Ӷ�ȒtM	dmU��
z/�)�g��'âVo��E;�e��=�'i�A�:��P�����&)#6i{�` �h����F1�ċ �ے�"�E�a:�!	#''��-Ѥ��{��0WޡP3G��y��9'��<v��e�-Lh\D�Kc�g Ny$Pׁ��D����� �t�΅H#�MBϤ9�H4$^0��;�e�&�Y��)Crp�u�����������X
y�lØ�7�p֐��t�賾�B?.�;�gw5e����p��>��=;0�ѐ����h<͕����؞�q��	th_�)3��3QxV^����~��B̤�X�B�YQ�!��JD�]^X����|:g2�?�\T��!������Izv)�����ASCrA����ٛ+�]���g_Bu(��H_ ���sNF�#�1�xou9:u�#��B�)�'G<�m�*��I�%C�����ki�e�յ�ؽ{7���c��/X�[~��m;�[�n���U��ODca���`����ѫ'W���|4���jIA� )"�k�1�z�:���|(� �ZLx�E<����TW`���q�����sG�47�#���mxf�S�no5���xd��!+Y.Ju1t�����
���oD�i7� ~����ر������z]\%�C� s�v 7IJn���y��n#k�,��$�)�t���Ģ��d��ٻ �\�T'i^_���T�����|U��Y��O��}dD�wrhFm��lt �r�[e��T�3��"�,�Pe�E,�d�`�T�d8�������ar+� ���*d�G�4���<g'K�H4�����@�D$$�>�8�H��U>��5j�x�IN�ڊS�LZ`PG��x��,h��I�@�8Ŷ8VtZ6�����CU(C�t���ǽ���Mp{�M:���q'\�[�x
�� �p�<6�+٦��m�YC�n�C��V���Hqo}�|mm}Kɔѣ�o�6�x�i��d��h�$\���"�JF�:����[e�UN-M!��77���!a	�C���řA)�x"A�PTP���<̝=w\wV��%=z�1E��f�/���^x���a�7�WP��6�����'���������P,���>S�y	�mX�����c��u8��SqΙ��%�X�ŗ��OJ⚆��aʴ��u=��I,��0�D��|�O �L��t��MCN9��&ܾ���e˖@u;�qV�Ct!(A}Șn�����_��ɓ1w�F@r!��b�p��D��
s�p�J:���%�]U50O<6�*0m�;���J�ީ�m�cf�L&�����1��[�ł)���0�^��C`B&}�:u_TdM���x,���D*��=m��-
�Q��s�п�1�>c6b)��¢|���7k�Fu�n��PPPA�������8�sر���n[�lF�.��#�y�����о}w@H��x<X��2a�<�7U��w�BUU{�Su��'y�?�����XU���ZTV���F~~�Ĳ�~܎��v��.C}c��#�CU7u^h�@ �i����E���!���N�:����裏�a��if����H�N`^��k/���9�?�+FSS#�W���j?�֕�%��T�ՠ�S��p*���I
r�H"e۾f5x�>��Ux��M�1@Q~lZ�=4�_�g�w8�S�J���$�fӸ�n>��9Du��a�U��-���e�X�������'F�)X��;��s!8�H�uh�0�� #a@�-G����n�r��"��h�w�BKBCJ	 m)Pe'(��2��=�PTT��g���=�p$gq)�Z�p�.т���G�"���{L�6��|�]�~7�\ݵ�(
B�(���U�m�!�H�����1Gv�$ƍ���%X�q-.�������K`%3���k�uG=D���G��ŗ��?��/�0
�h
-�M�N�9dzC�+׮������0d�)l��t���Ω���
�SFCS#W������@CDd�h�|�ɻ�hʇ�d�&d�D2����]�ߟ{2�j�E�c!dST�y�e�Gr��_�5{È���sV�id*C�@[�e�"q����(<^���mEy�n$S1f2]S���n�۝\�%LU�J��D��~�����T��aL�6� ��sσ�t¡X��+�U���^���w�þ��ش�[�q�8�w�5R;���ѵkg�~��X�~-w7V�^���ϻ ��0$�_.[�x4���?������M�x�u�g2`�g�E��%2d�I��vcɗ����^:�
Ϊ'@޲edE�_��zC}3�D�c��>o���.Z�}�8��;������w�bݺuL,$�"-h��wB�������A� ��p�W`��7�uӷ8�S�����WUagE|E�H����v(���DD�(�ă���(!���~��&��})�m������?��+��d�*�XE4�y�Ɓ��4��x��⯜�6@?n��~Z6���É���r$C�#�=Kv��C(៕�ѭ�~��q�}�R6�0G���t��d��={��E��h�YvB��=�d<�3����vm�y�7m"����UԲ(�X4w"J��>� :tꊊ�J�u����{0����q���ݕ�����3qX�B�����/Aq;є
���(7�����أ�b��H�Y̙?�� �Ǭ� ]�������s����DnE�ܕ�G�b<��3mKU�J��Р@�G[ԋl�v�7���y�a��������h�TL]��B�^��x�    IDATXi�I��CH�C���G?�Kν�\|~�5,q�����d��'b�JZ+��e�bK]2�!;]"�)0�E��S�����<�]"��Q�j"��ڿ��FG��N�hh�
�p��T.�D�����S<�?�=,]�OB~A�k���u�Ep��nE��=�v㷘9g.{�s��8���P'NĞ=�pd�޸��K�j��ٵk������g�E"�Ƨ�-ƒe_�y6l�8+W��pb��}���ܹ3����4�?��ù�&���/�D�v����w1�~��)زe+�����:�0 S�L��)�Owޅ��������ɂO��p���a�3�~��bT�W�C��r�)%��Mع{7W�=�$�zޞ��۲�xw�{7J���g׬Z	=��I���i'Ayy%>�� -��`	A@���`!����^(�x��qA�r�M4l5�ۃU���ʨ��G��3�db�9S� ��/5�1��cNkc�O�_?�6@?.=�����b]C(^4}�8lۼO>�<����&ƴ�N��r`�1j�c=�C��FT��̂�WI�2��\�56ǡ�}l|bZY8��&h	�gڂہ��Z(Z�u��[�#��3G~���g�푹���o�	ULO<�(F�x����8�~��ڛ��]��5n{�����:i
?�u��nGtGײN��I�0` F<�4�/^�X:�EK�"��@������|��7�N�;���沤�_��F�%���;�\�䦨ȦӬ��6I���#��U^���L���vu}%&}�6|�-����;zp)N��%w�;n���r,� �}�x�<��q���@i�	8!��O��d�"�<�XW�������@"��:{���� C�y,��Y
ʣ�v�[��03M�����~�ݼ�+V����ǟz���7�⋐�s�ә�ODQ֭�=�x�>���ӭkwn�WT������i�a |��W1o�|*Ǝ��U��[Q�n���h!E�v����'_k�޽z�c�a��믿�������íwލ�+V���c#�#�҂��ӧOG�.]��o /� S�NŘ1o��}��U,�#	��'� �ۍY�f��0���f��7߄��]��aW��];y��ʫ�s��GG`��y��7w�\clܸw�uK2�|�t(i��!�;��bD,��B�ia	r�ֱk����� ��6D�a��M"���A�E���%{�S�����s�$
����ǝ��cw���Cl���{`��/�<?iΚ���ƍE*äI2�*���(�!���c�z!���@%�/�e2:��e�C�z����I9�Pe �Gn���3��A�r�hڷ�Ё����ܳ5��1�C(�-a��؅�{ʑ�_�m�u+��������n��o߇� ��Q��;t�����lS�jA�~=9֕��C)|�q|�d3"�$�/�	M�iy� �,_���*9}^�:�J;u����X�z5:u�Ν���f�d�=���D�P%���M��_�A�,Byuk�_z�I���X|�b#��<���a�i¡���΋��oׯ�;��d�r�u��m�@*�f�D�S�}),�|[�9 �=xnN,p-E�4�W%�&'>Rp�&2��i �6�BM�0�IH��Hἳ3��Hc�ƍ�펻0������PQU�L2�+.�=��s�u�z�[�G��������Wp��]�vx���t�R��޻l�K�/��#F<�;＋A����HW^5���Tկ_�����t�=3��=W�d�s�Wb�M�:'�{aI	x�q|��<��?3�1�Jb��s�i���cQSS�Hj���`��x�B@ݳ_�r��5k��Ӊ��<���g�y��AZ��#���E��/���=˜��3�cܘ�||�W�����PZZ�3�<�� >��	\7<� �:�b�a�s�;Ud�EOr�a�|�4���`Et�!�Qr Kא=",��A�?
��)�`�$��%COd�2�W����~w܏�擮��*�C��0m�a��.\�
y��r=���T2���<&�8�H���`�'�sdo�ݽ�I;Z"���D2���"xyp8\�֥��)��'PI"kDn��t���	E];r`K��}()(Dư��^�v��+�^���mdӏ��T�4��o�A]m5N8v ֮�3g��eW]��5�&�X���Zj�R(�!���u�f��atl��}�G�w'c��M&�z헨��7�TV��-?�����9g6w�;�D44��8��去
ǡ���z���&�%��Rk:��2˞4��L����$B)���!�X�ݍ�CFIng��u=� P@������&�S��8���m=}�B|4k>�5��r'�"]��;��T�qI�@B�lI��	���S�q�����IHj4������T�u��Rat(��������
w�y��x*�S���N��b��oYP�o/F?�4N?�t�]������s�q�J߱c��P�>~�[L�������k���ODQQ�|�	�\���<� W�D&�>u��]�{��7o����Y6F��#F �`��O���^�o�{yA�z�M�����ޚ��}���^��{2���'!?/+W��Kc�"Ob�С���+��i�@��ԟ�yޏ.����%��kY�G�O��d:�)ӧ�g�^x���x�n��8��3��Ïb�GS����"����C�t@��G�N4ɮ�H-
��A�^�Y ;��8`)'�I�y�y��?:�A���Z�!�U��=�挹��;o���T6i�a��m+Y]RYB6�?j�H�9d<��N��.�[b1-K�X����ťAm�t�&c�c:��y��v�^Bq��,D"%�ܹKÌ�#�����3g�BAI)���r��G�S�nx�ٗ�v���_8�S�8LlٰnՃH2��X#6}����~��[�+�l�ĩ���3�(ؿ{'�,Z���^8}^477"��zx䗴�Kc���/`9�������� �֐��v���A$�8��%xr\h	7C7$�"�Bp��uz�V7Ӳ�<�$�5ըؽ�h3�:�CSs�hوg,&�=|��X�t5ޞ��+"ɯȥ,IndN�2�466"�Aai��D6�S���y��*�G"p��#Y����Nsd�+{`�d���ePm�T��&��ʪr(2��8�]�{��[M�\��c,�j��k�x�~������ѣv���2��z�=V�l[�u�Vmբ���f�4������ۦ�|*�����Ȥ}I1v���#	�62�����uNN.��r���#�|�����.��Pp��*���ү���e[�4�e{Ա K��ȣ�ѩS�x���]�x�wtln��6�<}D�qvE�!�֡�p�����N�B����\ȝ^-�hI0��,��:� 0�h����ZiE.�^����۬_��</��C?t���is�x��O�Ꞡ��2�MR+ς7@s}R��J��C�,/�5���DŊ�A� ���s�h$�9��c�$�Z��F���v;!�"+�2��pI
tjZ��1��7+���u��k�6l޼�SȠеc'|��f�z��xu���n�TTVc͊��ض	{w��J]S#��a
&:�k�bqi	�	Sf}���yO�S�k��:i��ѹC)�L�������Ź�Ͽ����,�>h���%�=*Y�f�4���	�dooÊ��s�3�O�GqA�T���3�BS�̙8��v+Zj����m|J&�� ��}�AX����%����)]32T9~B�..��L�r��=���yk4��&�}�m(+�Q/����>��%�W��W�BT�$'t�;UD���<o/.�G,b6��)2P���L��7�S|>��$�iQI�Y�>�Q{�[�q)��A�����k#�t�;����[����i�iy��_�Mea��|}�)d���!7�յu�� �;��r�455q��Lg�q9��֊�E$�,J�ߧ}�{��MS��R��c6�!G:Y��M4�;*n7���jF���u cXv:ai4�Dx;�S�I�t�� �6�"��$��GRU^�q������Ŋ
�ERfZG��
���u��ԯ�)��y��Ց��!p�}����>^Tw�Lq��M��V]
��)�#��LRId�:��ө�t$v�"͌���tB�lKά`!ih�ȳ���aĚ��^خt�M��pkh��ux�l�%B�*�,��;�Ǟ�۰b���UV։�рϏ��:\~�0<��s�[U��P˿\�D�>��tKƎ];QS_K7�TT��RJ\�T0q�|�75cٗ��u_������]:wFm�>쯨Ď�{a�*.�G���4Ų��x�JXGNc�H��u �N�o��V���FڄBd62Gq8�NG�p%Κ�o�;��+~�^=��G�>�1o�W<���͊��v;"��A�Tu��sΦ&4K��J��D=�d�
c_}Lx#�[o���<
{�U��ݻ�Ų�vݭ� B	�.7���D�#8[���3i�����m�t�9�븺T$��q~d2���FQ�B�m�ʤJ����CUm�-c"��rWH�����
�'vk�*+, �&���������]���l*ɠl�B�Hd�̱����������,� ��Bc}��O�`;yhaT_[c�gт�ey���/)0%�y�a��\��t������A��9yy<n!6��pC�X_�6��Һ�K��M��/
@���
���r,C�ȼ�Z�;�	n�Ӗ"J�z�̢@͆_�ˍ�����c�W���+�����<7i����p���$CA*�CX�-$u$�q���d��+H�_�?Բ���8��I;aJ�U�)��Hߤi4���t�vꄌ��kz}� {g��j^�=ь9S?����Вh��ACsg��1�M��~���p�c�aOU-�ugN��_/@qa.|���
��l��p����ӏ?���3?^����0��o�S�B�5l�~���p4=��������%q�g��)�5�GƐ��E&/�oI�LP�����U9�$�p��L6�tڀ���9�u�
Y�6���9�0��G�\[��:A�cx�ч0}�,쫨�֭[q�M7"���x)"��lk"&��v�LxN�"��#O���A�t�*�ɬ�x����D<p�p��ivh��_-��g������ $7����ʐG;������YzE�D�#;_�����E��c��x\n$	���Nj��FU-$����)�kGill�5�B�GLA42��s�V�	��J'�$ ��?k���v)P�������ΕI]�I�����!+N��f������"o)�����M|hVo���G)��%_�T*�ҲN�3\(̿fVc%����Waw���h0��)xŋā�Gn ��iډI��:W�:D#M�dMǋ4��E�d9 X�ݡ�0�ţʐ�.)��}�G_��w<��� ���oN���YKVEe�7�'y��	-��"HE��
$q:�֥**���-8	
��I?D"�Q����l�SU�J�8@"�hC=,C@a���<
��Dj3�L��d�XD+��{ N!�`��%+Pz�Z�p�$X*�v��y��3�$.<�Tto��� �`a������Bx��x`��0� �@Yi��s;�̜�2PҩG�����:��r�^�G�T�3o1����HY�����yO�r���"�e�[��T>��Gɴ'��)�T\0�4�L�{�?�
�N�+��0߇�G�`��܅_�����YٍQ�Ά��犗S>��N���| BT�$�ǻN�W���T���ň���7Ǝ��x1s��8�ԓQؾ���p��C!���S˟4x��D6M I�.biQ{�"A�0M�����"R�tRLH���8t�h.O��T"�"I9�Ԅe�p{\�h���\���f�H�d��1@�̜�kj����R���$�`�^��������XR�(K(��e.��eX�ɏ�.2��X2�:���
���q�y[��F&-�9Je#9)h���fy�����������syJ�#���&�Ñً//���qu��h�D��h�����bX�3�J�Z�t��i���nȬ�$)�M�x�nI"��N֯�Wｩ��g��:�6@?.��Y�z=7u᪈��|�|�]���ܪ��H46@��F*D$d���" m}����F� 7��(>7���������� �<��p4���m	��+#�EQtb���m�jlٴG�p,��c�o�GFb�+�Т;��A��tI8��T(	LBii1�++���K$q�eC1≧
'�Ԝ�`=�ĵW_���}�ޭ#��0p�Qhi��9u�'ࣙ���-���+Eʒ�6d!3��,��A�HƎ��p��o;g��K��0�gj�+l�C���4bδ�x���I���}�%l\�y9�hIix𱑸��PMc��k ys`P������%��]��|�:�C�?���Z��Z׹�\�54q��q#��"@��v#�Q5K�]�I�G�Į/H"GU+���1�g�t����4i�	�,@"na[������4��I�bp����)��3�h�Z�d!,#� ^�	w�˄I��ߩ@6�O���%MTֶ�]Yd���(r�d��r�
`*N�9�[.��T��0�VU�`� ��h�@5^Wϭp���}Zڡ���yr��΅fZ(n��,�����a`v�p�Z����*��W��TڄC��{�g��(<�t!�^�_�@�Y�SE4�`�_���KH����E�s���;��� :e"�E_���/lg9��m�!{�'������Z�R}AJ#pH��\�s�RO�M3S��)jV�#[,��$*� ��\6��CVv:�L��zV�𓔨��+��v�^v*+;�3"J�xΆ(,��$B�voszUXze�A���+�Y�o�C4�k��Fi�vpy���JT�'Y*�L�������i�OČi�p���X�|�Yga�g�PY݀P8	����ѲiN+�z��8n`��a|�n5���8��m�&�9���#�W�� "3dG�H�]��C�T-���yܲI�s��fƲ.:�M�E�n@�t亹3�@W�*��"��x4������f@�@��>�~�~��	�) ���f��i�A A�+z1�+,X��\�Udf��� ������2m����rX&�9��<;&�{��ˆ�-mÒ��ʐ�x�w�,�ꔸǻI�b�Ds'-<��E�;�ch�_{�%E���U��=y��	U@0����zԃrT1a@E8b΂%(AE�zP1G2{:w�w�.<［�]}������XLUwծ��������g����q��cዔ�rEfJPB�|A�ٻ��F"����!�i|����3�?�W�t��8$�`�5�I`'��!�"ܪ�{p߃s��b�e�l
�$B��T�Tk+|4f���e���-t��J�Lw�gRI%�a�nh����/+c׳DC��A)/C^P�[�2'�W�&BȲ�&;F�d�wZ�Q�^"# �����IV6y!nz>�3f�
�5��Z6����9I��M$���'�U���O�B���������ޅ�}Ԥ�N�y�y���!�hA@$)Q��:�03�6#*�lO������L:Ӧ9A$Z�f�� �F�3���ߵ�[���1ä��
gg#"2����RK2@��H��YC~��CЧ{O�<�;���K��|�u7>��#+�l"��0%7�j�K���٭+ҙ{L����h��&�Ӡ0U�� ��d3IX�$j۔b`�^�jS��T
o���mߍhQ�hl�ꮂ�c�*9�y݋�f�5���� 1��N�`Ôu��%ƻ�B�$�)�i�nf.�N���@M�
�qF�o��k���E^�U���2dͣ���2�υ�Z�%�k:���E�yڇT娢����*�JLB��z�P��(Q;'a[�y	���ͣ���'��Ht9�SK��sԹ��N-~�ݩz�L�k+�������    IDAT�ű�:ֿ���%%_ D}��$ٚ�?�%���3���}H4lg��#G��t�F�p=�6s�ɥ,��:~jG2_ͺg�=�������B�e6�OhlB�9Q��dO�o|���6|�=��'�*�Y5���N�r�B�%Ο]Z��%\Q'��BHvı�JdH|�z_�
�T�w󀑄�g�����ȥ=Z"-�5���ϥ��)ȶ�Y����Sb�
\��6Ĥ�@�V+�
��}h�%�G�o�~�X+\��%���|,�z�׭O,�0�Bz*� I��-�I�A�f�s=�b��F�>h��gҳ����N4.�hӃ��cG�ݴ:9�]"���_�  �G�+����BC+����UuP(�dVG8�!��ٶQ|��Yt�} ���f�A�tXrd[�E���p�%:oF6Ê\�M�4����g�Q���]��Xy����[&���02��H$�$Й� )�d�K�=��%(Jp�j���>���%t��=�W���PL�pl��$vV.�������!wC2�����b��W���aJ1�R����n��R�D�+3�E�Z��?O�E��*�9+��]���.��iq�:%t��v���Q���6S�f�CSb�G.4/wJJ&wsh�@	��T ��T�8pB�b%]�ЉS�+͌@_�D;J��ĚU�p���%�]Y�k&Q�[�.<�����߃_��~�6����8󜋐ə(��ѫW����X�zsc=:�V��Tk
���V��ڍ?BԂ��g[�.'��G�SC$�"��2��n�.� _����h�+x�[�5% �6���~+��� Q�V6�#��S��pT$�EZ`�]f�;��`@U���f�ڰz�@A6��"QW�@@��wē98�ZI)�45�~��>+k<4�#N�����V��BB�??�,[�g��U���/;��Y�YE!?2��9�W�B�X[É��妠��%��u��W7a?XAwE�@Q}��2h۱�bVM��z�m��W#	�N�T�`[��
QS��D��{���儕MPU�BS]�Aհ�0��J��s����S���1�J:���f�2T�œ(.+��"�Ȧ[��M�jja�,a�0"a8>�+@j�Ӣ�t�)��fr%Nml�R��-υIy����Ʀ�ц%�</v\�Q��w-�4�ϠK�6����(�ػ=zu�f]w-ďۛ1���H�� v6�aI!�	��ʁH�@-s�O�V�A�q)�{�4��]��w�؎m�ƻ�Q�g�*[n��k�ӵ�kB�
�ꂪ¥���\�3?�1�6��]9�G�z�Խ��;�/�@���km���wu���%<�����;#Pq�Q#X+���������_�I7⋯?Cm�C!�
l[��_A}CNu/0~��;|����IX�t���<���|��ؔ���3�WE�$�; �w��/M���Ǒj�s���QTY)����M��{7�#�^�j�W���a��L�,��D^"��!*�Z��#�&�$�:-@\R۵�n��I�B2��T �Qe�i+��P e8x��uH.|%5h��Њ�̜3���=��ao�O��U*���30���o}t����h���������	矱�mYtU&�-
�ZJb��/����;�Ti�HGG�;l�b�[Z!Q��*H.����!�t�Bqm5���͐�y��$���JCH�P�:�\�A<�E&Q�浄\�uT��9!�Si�B~��;'�(j�	G��Ց۳��BqQ����`�t0T
�_�_�ֱ^�*m3�HXE4���a��h�0��S0-J�5m #L��j��۔��AK|g��󃜄KdJ�.	�P_��Dj���-C��.�p�'tB��_��@m��;0�;p�m7"���ѡ���@O41�o[}o��9N;����oA	�~>����	1NI�Z�4���FP،ސ���9%_��h#�6)��.��q�i��k���Ŀ斻@�a�{3t���/����KD{�7��I��S@#�����K��0��焾��%��F
'��<��	ӒX2��qcQ�/����d��Z�6U�x��y�Ǜ��g_`�1g0��kU*p��X5���P��?���۰	[w�ă3g�ť�`kJ@^Ta�yh��cc��m�3��#F���d
��Cah�0ϬEBKS3�%4�	1��$�꾼���&t�)�j�����+�K��3ivʙ"���e
���� �
�Ц�l�ke>�ӣ˺�=���xS�τP�����?�j]��>������D�e�N����G^�<�
�X�������/�pϳ/��?r�J"GH��]�f⻶�>�k�J��}���>//{���v���e[`�+��UT�u)�d2�'�.)=��w�D �c�+�P�l@Iq�����K� }����������㞻�DǪr�(mn�gpS�OE,��%+pϜ�Q�� �u#ф~];a�7aώ�h׶���gvq���),���Ԅ���o��9ФYO���J�޽����O�Hm����9��ոMO`#�,)�̦�dF�fa/،�*R��p2%ГJ�e0ʜ��-wZ𨂍����҂�q˵W�$(����߭R>��;wC����8d��Ǟ_�PQ��"+ҞEF�j��/�E?S����%d���x����m^�� n��_RK�{-J�&ϟ�,A�@q6�������i8���|�C0I��oB�{(�_��r�ZWʹР�H�ނղ���[6�y$29m�+0j�ܧ;2���M����;����i3om�G�l��Ƴ�m"���@�>������b>P��O?���|�<�k&N�{�l�[Z`)D������OÞ];1��aÇ0{�l��14v�%U�� �t��&u!�^_I�%w[w����JX�>S�=E�>E��Ȳ#
=Y�T����f��+23)pM �D���vEihmM��3�޹�?zb-\�����_9v��QwL�U#��]3��8v��!��']��~�x��Uf�{�=S��R>�Ğ�x��9i����������85�7�olM�ƺ�h��/��Iv�
�D�P\U�T"��ĭIlxg6�h�u��Z�x奊�
�RM����ٔײe�SB��{�X��7W�t'B�!����1�o/t�,�3f0G�+GA�B��$QJ���gJ��"��N�JH�<��s�>����_y-R��D0R9b]wj3��<����`tM��]���D��i�*C`�/j){�h��k�Bv��K���3�Č�o��'qh�0j�H�CMU�z��|�m�:�|�nI��ϿF���H�:!{�U=F��`.�{ �IB0l�AT&�+g:�6P[ݶ�>�R�l��)V��F�7���8�Nx���a����򬜖.I�R��VDo�	�'�BR�T�(���˝�:ԥf'8�� �V<�F=�y�t���!�ѳKG�Q,-bXh6���mQS���x#����܇aC�C�!��p'�g�.����>��i{��~+-]�O��닰���(��XO>��صeb�"���./�R&�B�1����ʊx�a:���ܖ��PD^�{��'�WYA��iZ�h^W�%j\S���OzG�=Y�<zwl�/�+�����_�����ߟ~����_2�ɷ�R��6f�z�G<W �fa��"PH���-n�k�f��d����-�����^);������ׯ][��w�
���g-��D`z�8y8>��UE��v}=�{}5N:���P6��VN��`���d
:y����N�7�Xdi�đ#G���3�?�8"�x���9,,S
`��w�����XT���^�!���_~?��En��bd��K�/��\ ��-2q�-����R(ARD#yU���	AN�r�"�8���Q��r��R
�E��Խr���[�i;�z�5����׻�C~�d�L��i�nڄcO:Z$���^w�ÿ�6��������̜��.�6濲�l؀@0��<	�M�����#�Z�I���&;ڞ��#�\���y" f�g��P4��=� 	ٸ2y�p�T�`��id^��O0�<��m��]XQб��A�(�0�&��#���}lt2���3�4�7!�\lٶ�|��~k-�-��᧟��pn�w�)A"ш�f�d4<�.I��C�U,mv�Ǭ����O`K�BʦI�Ur!�S�X��"�?/�`�ct�H��	�pI��8$c\G&��E2�~���~U�� O?"����.���x��4��;��"�]q=ږ.:}��KO<���~/i�SƜ=���:n��jw�t�C=z��TH�%��s�-$��9��?�����;���56jS����k=���O�[/���o��+kVo�ak��_|��kE?�� -d.��NChj��+�����;oB$�b���`�U��أO`���L�fyY	�v����u��Q'a�������=��z�ZƢ~�ƘSO�a}����㢿���>Z��=��MM�}�i_�kS�[�q2<��S�Je�t�R<0g6�r�����E�z�_Pվ�:oI ��CP4���%�T=�����?Z�{���HF�d�A��Dc��R�&T<���&��٧p��W!���Cz��K.�ꕯa��ñ��Uxe�J\>�*�?֮]�V�WL��C��C�]�iwMg��|VGiu[�?�2�v�t�.i0,2	r��M)�9O#��ѻ{G<��,��q�om�s��i8��1(�l������Sg��t�G��}���:w\5̟�F#��9�d.��%�|�5�ڭ\͏e�_���s�����0�Bl&by_�b���>\��@P#��,��O��hۦ-��4l�e%�W���ɮ-?ᓏ����M@�z�mSEv��?✳�b���[��ڷp��ix������͘>�v,[���r,هP��
�<&pm����r2WCa��;[��S��|>Ċ���YF��-	n�[>Z,�xb}P%�2��|���I��/h9ȷ���֧yx�5v.���}P�㮼�~��򫯾j{�=w�uک�t��.{��Æ�X����o($����/^�j�ԧ�sDIxt���-g1��˿���9k�����%����C�� ,�¤��XeT2�7�%�1����vұGaҕ��Ԃk���K&L�w_�}z#���[o��9s��Ư�WT��|	��ꃃ�˯���Z��t�N9���ƲE�a�a}Q�gν�Bl�ǧ��h�L�+����O9N6�����T�����5o�G�~��A\s�](n�����
%}��ڽd1���{�ĹV�R���ل�&�9J�4c�(��p�m̕���e��Ԇ��{k^�M����_~�e&��ڀP��T��R^H�?�"�t����7�������Ȓ�o���w�A8B�1���m�t�B8��x�@��E�`�Y[f�j��~;�x�U��qXFÏ���Mw܉X(��Ӧ!RR���7^w-F�s�}��b4�����Ÿ/��7^�����@�=p�%1宩�}�@y܉P#%�f	]��O�*�iٞ;Ѵ� ��]x1d��F+O�F��mצ=W�9Gg�[+g2=�\��>�#F��TIiG;�w�b���9�ջV��.��q����/������V�<b��){��$��A,�rǉ\��l�,���ˣeO���)-f~:�Z��a�f!i��E@(��O�M���5�Թ3BT7�Xf+�W�*��%���{��t�7]���;�ޡC���6X:��Ba��"PH�����x�������J���5=�pAȒ�7oo����������w�Z2rY@����ycQM9|"km�+/>���z��,��Ɯ�}zq����W2��ǥ\�t2�����'^�L�B��	��z=z������-3fC(n���X�{p���8���x����s�e���Ba|��wxe�j����5��'ӈ�S�ҥڵ��O[���L���'݀�N��u}H%�H�[�E��C��
�̐,*!ۙ&�I���Kr���HF����N0���E0��y�v,_�+�o܃l>�p4�`3B��x�/F(�܇Ɗ+���f��m�*+��c��c�A���q�M���o�f>�V�Y�+����Ȋ�����" ���2xx�t�{kҩf�}:.�p"���z��"�o�����C�ݰ���dR������&���8��ӱh�t��	�;�]z)�=��x3�9i42$L�|v\K�,��6dգ��0KH���^}GC�s%��yvqs�^(+�51��'Op����?��:�?o4��V>��Y�� ͫ�OpY>�$e�;����1k�#����d�qD��H�5���A�n��R�,�d�;-$sL�ѭN�c�WJԁH����њ�#�$Q�� SI����mZ*	3���J�1E���N�h�pP�n'?p��~�r�_lXw�'�ظ����֫��X��7������cE����X���l^^�b��O�0{�����է�f�r㉿��B3���o}tt���%�$K`�V������hƲyO����0h@\1�BTU� ��n�)g�����c�s/b�ĉ�r�\p�x�K*V�xj�}��2`f=��h)���p�)'�o�n���k����oi@��v�񗟱e�Vl޼�}>��c=|(+�QB'���}���O�#�=�K��NEW�� �y������l�ҧ�{�	�xI�8�W�,�J7#/�f�ϓ%�P'�4��b"$�*6J�1D�L'�1Ou��B29n�S���5��f�P ��&G�����,�H]�2�� [[�L�&�xf[���c�P��{�,�·�م�>�{�~I�%����^�s��W;l&����(<c?㴓9y���A��d+^���o��~C�A�^�+'!�ᬱ硺s��m�M?mf�>��u|!^p��mPI<�`�<+Մ%���SND��-�#au�v�. �ӓ%� ���*�&���e7�Jo� ����2���n��I_��a|~X���=�߀�V���4K�ʲ�����H������'ݚ`!�|� ¥Eܭ!�����I'�G��
Y��m$�^�K��P���!�� AW4R�ki��Iz��t�$��P�F��X�����8n�������-�}�~ç�v��!ѹ[ב�HM��}��q������󙿴l��iO̟~�i���ךּl��ߝ��M��ztыK�S�2�#.����i.o!ڮ
�`×Mb���0d�A,�zH�Y�=��󯿃����4jʪ���ʍ�G���~�ݛ���k��G�De�q����:ɓ6����CѶ4�Gg�D�>ݘ�^\Z�H��?��+&��d0�����۲�TVU�_6�i�q�WC�9&=�IW�=�R�7	�ҧ���5���#uO��@$�&QB �⇾�Ȱ	3�z�aM���!*G(����C�d��N�CR5��%?zj�S���$dR)C~�?��ap2!:-
�}��Ln^$��W=3�G@�1PLvl�Wz�@�9��L=����op��#q���`���J��@R�M8��c����CR�\��w�������qPo����*8X��eth�]��@I۶���l|�e+�Ί��]@f��4�܅|�l�D3^|�1�9��e**+��(���T--T6�ڊ��r^�I��֦:;�H|��hnjEuU%;���Y�R�[q��֦������:�me���;��y��eI���cH0�D����'	�4s�IŐ� .y���@��8x��RYD���Y���(��?
ˑ`�
w���'S��=��ɭ���H�&N+ڗE���+�u��-����w;Ʒl�-Y���^}�9���BB����sWH����Og���o����N=c�un�b�С�����`�9�����V�eks+�d��:L�AQ�j8���U/=�^�:�$ !���%�,��R褚�h��L=�6�U����0���Ɖǝ���շ߃��}x�H��J����NAPs���O���K ��4'�̥`�IF3~g%�  UIDAT�ri��#������]�x��U��p&����Ma�s�ٜ��,��E�w��r�N�kh��TE����6� ����(hI�>�@5e�ihA��i�����M�Fz�^�O	�	�}�e��g$���ӆ�!4�����c�-j�࿩�6�<$�+z����x6����|lUJ����$Z���;2�C~�T�eQ�B%=w3'C�������k�k�Ke�ڵU��	ybP?Õ�ͥY������%Q��*a��@|4@w�p�̬�`$���BIiR�,R-�(�kAB2K`D���F �����P[�D����,K-�E�ؾ�	Z�,�J����!�[,��*@sE��H D>�
��V�W�t����J���0����u��u�4(� b�$$�B$�u�D�^Mup�i�,��V���$:W�6_s���ǜ|���{�e˖�;�֮�x`�l�^�GW�*��k���F������n��|������3��n2�#�O:��s�������U7�������lț�HL�E��ðl�նc+K1�ǫ��DkC#��E~��"�06}�5&�1��3Ix��oB��ʉ�����p��greuǔ{�x�
���P8��=?�4������CrLO�(�%Ռ~޶cWMG�'O�� �L�g��M�uɼ�Q���3k�_S�&�RAT��E�.D�"�ɩ��|�)a�+�J֕pP� ��"eIU����O1�;
c{S��Y$JcA����r���3����њ�@��^�`DO��2�,8�(+�V4�4~��? k��EYFK:	Q�`�*���hH�&�Ee,P#)��REKjw
� d�\��W��'��A(������"�l
>Mb _��� �vo�� 4�A7�Ƒ�&!�ʛ ����^sNu<�y�q<���3z"��W��W	��C�i�c���|��ⲿ���q��w��]5ο�4�7��/���Ϳ����0��z��i3���_��_�9܇��jp��q��I8�����q�M7A��<C�$��c�Z�<�w<�����"D~��,��jE��sN� O@O�
*�	Q�MRXS�S�gCK���&!�XW�AR��\���+�n5��^v�����ݦ*7n�iӦŽ�u�޾s�S˂e��w�pܟ7����w�|�K_[u������ǡcU�{Ǟ|���n�����X���u�Ei�@��S�H%���ԅ�>0I�łF/�4JB�V�+�P@c	OYSoMB�m��Q��U��m����ߜ��O�i���D��-��e���75�q��1�⊶�2j�i�	$SiFKS�rlv�"K̼nrH���Y,�!s��\&�~�?���6� 6v@���9��$t��²������;�#"��Z<;�>N�?�o��)�8j8&]yn��*L�r+��q���/�g�s�8�B�;�R4gnU���M�9�N����9��6��t3���>I���`Μq�y��+'�s�>����<� R�yWA��|����G4-a��8!��.hqC] �G����N�/��N�j�ﹷ�IE$
=�E�߸�ݺtF��}��g����W"���k�v��=�T�rұ�����s�̝������O7~������;/-^���#G��Ï<�c��cǲ����-[�A�T�m����A�~��x�gx<p���;�A�����CM��hߩ#N;��K�@�JS6�!�;B�SW�: �y1�?sF.�d]e	�p�1�~������5|�(�(�0��ȄG/2�o�Fށ�M#�N�����0��8��*��^������K��v\���)u{v�ֽ{��C��7,#�¶�E����������|j��v���k���+/ׯ�_��{.���/_�ї�=��?�bE3_0��j4/&���v��If I2����q��a�r����z���s�Ű��t�0�������[UQѦ=���syz�76֣��E!Q���©'����
��[n����~{�Y�0�����9�N*f�'tV��hNmp�Enj�
G��R�k+J�l��)��5Ѣ"L�\K�b~4��	�\=����\�7�E]PU[�ję'һ�ɆOp�q�e7����S�GD�@���g���'����=�l��,�:���q��`S�����k�'Zx���c�-���f��'��ϡ�]{<���X0o>����}�F��a��v]{�Ǟ�.�)u�i�{f*�G�m�ǻ'KJ�a��|ީ���r���%�������~��hmA,������m��w߰�}8�`�3p����Wa����C6��$I�3>�K�,��g��iӦᤓN�q��m۶a��i8p ����q<���[���	=��KJp�\�;P�.U����b'(�T�=b1jS[J�X�)5��ڤ(��{�VI���jQ3�����������9������}��\7����f��>��(���b0�V�ϜGl��u��������+w�u�(s��m8t��s��A�ٟ}U�β;����ci�U��*4gì T��kp S�-�5�ϋ@��ɧ����(˓G�A���-63���y�p�B��X��Ug�����`{�~�$���+��_c�=o�I�Y�HZ�����]����C��K�^�������j˽���m-ErU����6��E2��O�͚T!�!�7_R��$�(�흗z��bkZ����*v�ԲRW�P.��H��E�c�VJ7��
�k&�U�D՝�\B�g`K�o����F�;����B9�m�wYFrǰ�ӏ~Jw�ӐV�%�û��;G=��)�*m�����eZ��L�Q����A�T��eN��d��p,��LUK��2����#p$&�]BH����73݅��#�{���h�a[�`�
u��d��	/jpه��%A�:�S5���q?0C[(<~�򥠋���=��;fcl�*a	ȟ�$e�B�ۨ.���c��ã�p �}���+ &��.��z:���������i����ŋ.��/C�8v��q�N�EX���ˤ�gƌF�o9�g��8�?3����Wo {��������SM��u�|���Q�Wq�71�b�@���h�aDb�S�h�h���V�~01�l�p����f�����s�ݞ��S伶����}���{��2���%J�!�����xQ�ӯ��&�Ei�256Ł6���Y�Zӛ����;��m�)d�����7,�y�n����F�+؀>�1��<�F=��*m>�kU�hr8i�Jd��T>!Ӧ?�a�������e|Jx�8w�_a�{I9��ف�l��dQG���Yz5���:��9#�x�Q�Tɺ�H�frp�͛m���|��ވ
^�&�?:�ӄ�}
^ff���
�Ig��V��T@dlh8�����e�z�=��^F�m�{/ǚ��^77k�nGm����\^�픸��a�[�D�:��+�$b���dx���J����*��HŖ+���s������¯�������Зw�ȁM�I�\�,4�)�S ��f�3�g^�p�� ��f�r�V����_�|��5blb�ЭB#X���k��qH�ݹ���I�ZC��D��,oR�M�����?�S��f�\]�v,@�+n�^z�[H}�=J���^/�S6�?�I��猽jTw�X�r�:�@v�������E�&��t�ʵt�ra"L�V�"�T&�݌`6��	�@���F��Au��y���g����3�u�\F�ܫHP�0A*ZEi�Nӏ1�4j}��A�F����|(�J,`��Z"d���R/����e�����̧2�Xq�a���1��zk��ͧ~[�n}�����K�����u\��� ��O�V�>���2;=��j�7�`y��|N�Q:IB.��E�12f��ӷ�ID[[P�ihd[!��5��d�Jz�p�y��q�5R�(<"݁S�&���8�]{k�qu��ھ�ra��z�~��I��umT�7L�Z��"�j����Dl{ӕ���>BY�
����O p��_M7�a���!ёiqf̴�����&�y�^��bLywDB��� �����5�.��ktx=;�z�@���h����.(�Tu<���Z�9)�Ԇ��	X¶J^��잲xt L,�?����H��nA%5�&�ʘ�œ)��N���A-����ڲ^�i��ե����gOr��k<Җ�	�G�IW���%Y�_f�C>� �xBU��g�a��i����٩lܗ�	��������X�����d��[��+�T�25]���I�B���	��k'�����}�2��b��C/O�}���؄\��J��~
y4U�n͞&�z1P+4����a��Fޢ�4s�[��s� �B#r�M�r-u���S��/G�<��R���V���A����*��p��ް����KW�|����h� 99u����49��_�Dkc�_I���;P�R��~zG�����eO�.�Sx�n>��Y�N*�+}�+Aޝ��=��A�˧l�2����|�Grjh��w&�����w�g	�����zd����Bɺ��!bf��fP���v!�O$�@�Fƚ'���o��I�R���d]�Ck���g`�t�D[�I�6���@=�sT�c�jk���&=�:mlh�������o�j�I�8f?�������HُV��]���KP��i�h&��� �@��T�F�����Զ4h���Ң�����.��b�����hg���n`7�h���/�/�v�)�*������F]�g��c�K|��G��|���>^B�A�mf�C�ϋ�,��0^r1����;3Ԯ'�K��O�0]�#��7!]S�~�p �>U,�uu�4����1�Wv�";H�K'�!��{FK��C�vG�E�G�;U��\�]���`�~����ù'�"�w�1J��U�	l��h!��D�ĄB�"��p���'{ �f�ũ�EokqD���
Xs.`�"���P�hl��.��F�g��"��[��t/8��ߟr;�%p�θ~>�<�5߮y�oug|q&����Rk8>;��چ�ϛ^�$�V=���w��- Ǫ"����.�ؖʌ�p�>����]0v��D���ĥ��D/����{�S�w����!���1�@N���ף��9f�b�>5q�
ǂ}%r��a��U�:�h`�8Bf{�k���f �z�+ygI�J!v[͗��t�lL�Tc�>�U�o��7�W$�;��?��>\��5�&t�^��z��k�qW@��ѡ���"���O�)܀E:ѓ��1�V���8,N��`�6{�X�[�O��7;�p��Z���^�U�@��j�6s���e�Ȇ�!�_8==�������Z�oW��|���m����rI����� f�fE ~��>ڍ�&�w���4�,��������4I�o;������J�W�ds������%$�����8BTΏ�ha? ��*��Z��S�,�[�լ^.��Q�&A|�����@�0+��FbY��m���<^鬇E��S���` �=���r�I�
TLt��7�tX�6#)@�J��H���^#_��rl=P�*_���E�{��r�x����>a*Ty ����y=��O�O\������*�T��J�L<p:�^&���4���(y:��LmM3�J(�{j�bm�2�T���A�-\K%,8"y1���ITGM�	��v�[��v�ːK���W :�|Sr5��'����e��[�h(b@�5@�q�iLPm]����D$�U�'���*�Lw��^�d�RK�'�Jv��dD����j�*>���G��h@0�[73�-��0~�T�)Y�h��$��up�۩S)��R:���%Iu�wq�G_-�@�K��d��pH+% $�
����h׹?��?�eJA�����0���bYs�\�l��M�{k*����ߍb6L �{��wd�=l�*7C����漱��/O3�E,����(ɯ-��ŕ&�-V��6��!h4���7V�����<�
?���JF��*T(M���1 '}�>Б�����0�0ᔑH�PZ��I�	��106�Q�`>L��83�B�˛�,1���N%�3�[��H���@��M�Ԥ��Z_�qPD�ۅ?�X�@*�]�\9��y(JO�t"��L��k�d�L�<���/��4�\덿�	~3.ٺ�g���AdM�3I�&�.J�p:VG�F����(0N�0>@��lU�H�ƽ�b�}��vJ�&O��~]]��G|\�`���;4� ��|ƤjZ���"�JB�Ty�VA���ޜ�)�Jg��%Vn���o+\����u\-4�`�pgȋ�퓏�,1�
�Ĭ���!_��4�%g�����V�N�y~bP�ç�����+�GF}{��&)��b�����ns��p pΛ�7������#�]�T�x��;/�e����|�KH��U��9����R�a�)t���s��O�7��B�y���(>g ']W������ɫ��w��a��5B{���cQ�E�nx(d �9��9W�5k�h���57���y� �SR�m�3��X�E���t�sV�j��r�(:�*`z�_Vw��a$mb5�]������W )���?Ԕg�wj0�ܯy���Zi���O��6���S�/ίp�W&�w��<h��֯<��Y;+����ۍ�+���]�S`�䱵�����e�b.E����,:i�Ub�J�_|m�Z1,ۓ��p�qm�tn*Apb�o8����0�7�Zb.[#T��<A�����aû1t]�E���l'�"X{AA�
=�lx�G�j��c�	�{vA<ζ�Yoj`��Po����+rsR.����%�bSjs�M��.u��q���۴�����+#���a&.�W�(��ץ]!Wb�c�T��b�V�;���dND+��h��V@�=M�2	��M���n�R��/������/����P���pOW������y�{q7؇���q��]��;Gb//�����%s�\Ht+��ō�	�U�R~�PK   "��W��L�h� �� /   images/505d58e4-7e58-4ce3-be43-3c0c0a024e39.pngl�w<���>w�޵ku*jTՊ�U��ޣUTc'���(�*�V���3�*A��J�#�nl�+���<���>�?��W�\��:��}����>��bf�� ���h�@T�����G��T0C-5P9�o	��ָg�o��E��x��l:�`�������ݧi��44pcy���%�S�C��_K	��U����z���_:Lq� F1~���_AgC�̀���}z����Y�x��e��)x}B�}��e���y���j�N����y�-�F�\�� �[�2D����T���H�<��K��*�o�<��������������۳�_����AE�L��_"�>��۞�N��o�;/�?WAM�{uLy��l 	�ȡ��W��W'���Y�>�J#B���ʸV ����@�[�{$����
��L
����M�f�3��ʮ�A=F����:��G���@���-؟[V?k6��: O�U�9|��R-��+%O��y��h�4ТӌZ��K��KC��Յg�Kf���ՌP3�)6q�alW�~�d��y|���{�~vKV��f��u�|$r��Kޏ8�d�OH�G{��ޤ��$�����fD�1$|�݋~K`*�1+-��`��$�_x��˥?4�Ze��i���5����Y���w���F����M>A��'��A���_��  �r-��;�R�B��V��
[6��5�&��^Hȵwnl*:_����_�nL�y?�9V,&X���E�������&���T���	L�q�FG�wˡE�4�
;����5-��M��l;
����:��Z��1{M��)x͇�]u��*hQ��/�'���X�w5��V0J�J4�~a�]�� �DҐy��X��eR��Y'� ���9�7}��3����k��Η�/2_g�j�c?��ժ�&�D\�X�<<�e���S���8h��m�H���ҕ�i�����L.vL�$KjO���e�px_̓xݪ>��=R��mUR�w�0�����EJ$ݻ�ZI��K�w;�un��J�Ͼq_�,�Ps`��+��bt-�j���{�$&�B�?n������{��A�(XO�`=+�CwH5h��C��9p���_�E�<�g����mR�&�[pZ�]1s�.��N�~�A_��ז\���^��w�ϧ[r~�;Λ�_�^JOu��8�7�p���Vƕ���%�9s�W��T�f5��ĭt���ؙ���V��q��ս��v��p�e��t�xX�0�^�X.�J���W�:�p-Qiv��԰��C�.�߲ Qg�M�����~�kӫ϶�:�j�|��,@mn�^�����S�m���~�^M_>��φ�k,���u���"�Lh[{�RӌrTB�����~��
|R�(��X�W�9�F�S��3;�ퟪ���{�&S�)�VV"I�ӂד$5R�n$��o$���|�t�9������\���x�u�B���Q���������W��F��@�f=����Æ�Z��R<��W�I��\Bh��MiVw��#%+��D�r	_IBi	TD�#�n~N�����8�r)���,VX�%#�]�*X��fld���VM,�JhY~���TxM���ӌ���z���'3�X�j�T��r�pu5g9G�0@��n ������yv�Y�㓣��`�9�x>C���7�_�72��~$�܋���4��Ҳ"j���49ZYV�����[�;9Eb����q*G:��y^�<���i���L߷�����P\]]��p�΁;�~!W��D��74�B���>��!������(�?�JGk����sz���@�O�;�i��4��\[_���["�7rh�E�[�y������W��|q}.6l>�l9R��D_5�0���u�mf�m�F'�Ќh1��gu��u�j��]��f�f���9_n�޺�r�N�!��	]3��W�_�۠�G��Qn���K�{���:iΖѿLU�L;��͑'�)�T+kX�W�;::�>R����|T.ϞR�eMA��?�7�Y�9�ߑl��vD+��X]L�e��z�@׵�\!�q�S�u&q��A?'8�Iz��d��O9��Kz18=є�k�l��	��b����ϭ���Ҙ֙��yjG��C����ޥ���y'�i�L�T(yM3�����ύ���JLdD�2=:K��C�>�Q��Id�Rë=�� �rs��ĸ���׼�--�[���~�������{���怜 �=�Ԧ���w�p6��k�2>}M�n<Yy�ۑI\`�Ig�Oӌ�i]�C�J���z	���,����I�ˏ]��ɤp��j(��9��p&�%G�9��$����.,D+Ѿ��^5c�
�V��16B4��咟 hf�x�D>^��s��Y��[~���P��f|�|�r��r���oEE��VW�!k������m��4@(S������;C��#
vC
|� ����*�G'�.�>��Co��3�V�
1U.S�Ə�	Ot�Y�&������������D�@���i-^�ٟ���|k�7m�vDF��n:��$�	N�$i}X`3����G�\�O��Wy����#��gw��� ����HI����ߤ��	��p�RW2�{��CϾ�ڒp��q� ��a [y�,MJNϢ�Y��
5x�i���L�� ]��%��,���x���i�:7�S��w�PHe��WE_�����i8v�4�����ɦ\}�a���E���@a��$��A��X���y'xv��mF��㬃��Yh�T��o�QMz]��X���F��q-��8#˽��:�D(Ɛ�<���'�i���a�/�A!��c�׹�M�>zM��h Z��&,^~���u��ײŁ�a�c`b��2�K/x�ccW(&�0��K�q&�9��Z.P��CN�yU���C���En����������uqܤ�N�u��zT�Q��4U���<	�zi�H.;��4t���]
ƍ(֓�2�'m���F{pȷ�	�6��K^����!� ��������
�h�3ળ{�*�	T�R���'�[�޼/���
���o�t=Rڸ�2�K�����V ��69���t˴�qjp��'��*��7��t���0�\��N�@�t-�U��U��n?x%zm��[�����Ϋ����_�a��x���v4�WXRb�Eh�z�|��y��s���y��F���|���I�tլ�/G_y�S�!7r�Ȧ�|(������XLh)0����`�`x��*���6�"��t^rQ�`h.Ȭ��b����TE�uع�k-�~HE�l&އt�I[l2�k��� ���ӂ��\���}��>7-M�%I����7��$��	�wR�/� ����ߜa?Ed�,?��1�/*he Sb�;�M��ݚ��� �u���u�����Z{�Zq�=9:����O���P~@La:<��-�����v7{;�32r?|�	s6S�K��W�/;jsԏ��Jݗ��Ky�a*p�,���gy��T Lހ�E;�]l���Ux����@���}�N�Μ\㻉�.��a�i�A��X�"�t]���g��nX��r����(�5(���O��}��78v]=[R����X��@���o��!GkS%f���h����o�
t�J�{��e��s`O3���H��G��X#'yHE��������#��fC�	�0`(y������w���@>�<�����AV{����9rS�^�E�Ek?�tp��]O��HXuIXl9I_������#X� .E��S���]Ca��e�{_�TǞ��7�clKń����?*�η���:[v�#�0}� ����bP|0T�*rč:��7Ii���b�Ȧm&���U��J��GF��D/���nN�L��l��Wd�R� 
�`O�_��e�㤼y�����2�K�j��)�����$K8�:�\������A00���g���<�q��3�"GQ��H��b��	'���&w��T��\����z�L9[rO�}�	'��)��nx�uE�ˋEž��b=�-C��i�F.�(�!唫7��{��������#��F.	�<�M�Ԗ�q�cz��yMM�W���W��G����&<П>}=��&��7N���-�+�~���ߑMRq�kz!Y���I�U0�t��Ǉí���FR�g�r$�K�E?Z����_��ӌ�م���E<�Y��\Ǘּ<��Z������x���{����M�AX~\�`��;�X͂��a
�(-E�O6�+�����������e�:�m
��Qd����j��&�9����J^��d�Gd$8�+s��cߠ�Kw]�+�%�͟�;�Z�֢<7�>�z7M𖎚
��J�n2)�6�T�����@x�p�&��K��I*�$�d!����ߢ^��%&Hcy���H�Ax]�	�^��X��=y���	.�&����h�Ȃd�K,�<>SY���l��X�8�G������������۰���
I��0�;Rѣcjf�&�T����%͓E�vWr�M1�(?Cj�|Y#qV���Wts�a�S��"����K��P�4g����NklZ��\�h��M��E[�Swv |}��Jζm�է��:>��%��U�͸�iޮ�%�U��J��/n�vz��~�����a+����u�6��ܓ�ym ?SP�\d��/����0ܴ�s�e	������,����"F ��C}�H�?�,��Q����)&O�%�I<�J9���=�A�N��7 ��*V{�p^~kn��꒖�l�۔(ח�/�?dxï����p�4"�5��⣶�2�#TI %�iģ��(k���+,~߱�����?��5����#�m<w�!`2R�Ҍ�$l��v�K��~�==��WWIa�ؿ�3(7}�0 "����=(?~�c��GXȶ�Eg��p���'MQ�|�ʟ����24�>��&����Uk^�K�[%�6�7Zp��y�R�Y)6�S�W���;�p�Gfv!>��g�`R�J];or���l�3�=Fs�)�@�j~%�n��-�w���%�����Mt�b�7>��W�����ebff���x�OL�4h	�5�\$pW ��B�����h����D������ru��[Y���,�0��pL�bu���'&,�ˀ��L�q	��	s��k�kv��R��,,4�V�7r��C����>�x��KC�c�<�͐���=�+�vvz)N�[�@p������$t]j�K����u�V������B��K&|T��u`�:�*.*7����%,���&��?#�����s =��l*h#���޷�ؤ��!��0v�W��;�/ۂ�y��,M�d��se�҃�.1���e��7�F���fM;'by�k�M��T�?���a�~�1��=��~���[�ױ����7Bn���B�Z���r��o�c$`��[pe)=Vg)6"�!�WϨBZ��3�ѣ�ʑ/z��P���(M����:/h�D�*�ʸ�<���>J����%^��b �0�W�9�-��o_{�;���A��&�1 E�Y�{,��H��=�AXtMe�����Gy�Dǝ_<�����X�ǐC=�f��]$Ou�b�:6>�A�R@�2�i��4#�����=�����7!{�na�'I?�)P�T!�re� �~7W4{���V[WƊ��z!أ��������#HEy���������e�Hz֣�iп����b4� 7E:�U񰬬l�c��lԏ�r����!u�X�����$nP��#q��xz, ���$��y�v�CR��¹���'����@��U�7@<`�?�Ok$&����j��Ŕ�ʹ�.��I)0��_�<�s���p����5�I7<8��^���ku\>|&T�E��;mW�7O^�!)פ۔�k����RW#�)��\�%��C�ݳ}'�[�����g��9��.?��}��>�=�wĩ��{3h;�}y}�
�=�cQh5 pR�m��[����@���d�����ۥ�ન��~��moE���$������s=O�`�m����%��O�_��{[e&�?=��B���é���N�
�������d&7F`���(�Suu��g}�YWrcn_|W脿$�m�Q�c�䈤pw�\�}���"�0���B�ݨo*q��-yo݇ۧB7<wg�g�u��Ph
d���޸�v�r���zS̶�\����ա���g�����Y 8=����u����˺15td�!��m �&�m�pN٘S��1Y���I���7���l���˖7v���eUvn9w�`��u�8npG�uDꗎ��Q�8�3	+����j�6��hWNs�V����u�#R�D��������/�E�[��R�t�C�������>�"	� t���#�47�.��e�	ʊ)���Cxt
�Y�����
�T�����KIg~��g����(z�z��d2��.� ��k�����"4��� U��Ԭ@�؆D�T����k��"T���1`���c����뵠g#�c4��,N=�;� �� x)Et�W#�ۈ2�=Gh���/>�b9e}�@���+O��}�(x�O�T��kN�}�>�!�ť��n����i�2�7�i���<��QMI���M��uN�	Do�]4�!q8�g{��
�	�1�����Z�}�4��	��f1�����E��/p��|�5�zד~ΦK5�b�28����tME���%F�B��0 ��4z}c�ݸR\^�h�sI)����'��>@��)ߣ��&�%@־xG���3{��g�)U��5Q_�	[1[��tp�"�m���mkten���nhד�Y3U_�Ȥ��:bl2����?܋�@���S��9Rwu2@�!�����{a�������՗ ��GQQ��do�~uM�\��{��Z]У��g�C�[`sx��~�?��~Ѭ��?�f�Ҙ������p�{+dRn�v0Z�C��@6K�!�EZY�P�zCR�Z����t��mK�u��R���oa�Uʤ�{��j �#�⃁�ƌ}[W��*��7X,֗j�Mcp��Z������V̓ߥ�����5�:�%k q�����-]*�%�w�m��2��4Y�5��@���܊h0��,���d9(����wy�ɿ*��[��|C�GN����R�� �K	���Hи`E�����"C�Y�:zD/C��i��}}��0G�u�G��=A�Ię��17#k�QP��0�Y�%�<���Lngy��vƛb�ӍMUk�u��l�$`5�ܯ����B;2M�r4��,��Li��_�V{�O����hG�'��,��p7QW�
�xdT�2�mr�Z��%J�z�|H�źX�)�ll��G�D
���G`C�dj6�E$��Y��#�{�c�����Q��c��~�J��ɀm�������|#ak�w�Փ'5݃��}A�^��cT�m=�A��q����n��t�m�Z����>>>Eٲ��'�3s����tTV�SB��0=ȁ�E\g5��m[
m����*�V�� �Yd>�P���Wp�kӀd����D~��� N#���9ZPS�
41������[1x��������#��6�ڣ�`�T�ms6�Y)�AS�:7c��(��$��Lp�_��_��R��V�`�w��JW�(�k^nm�P�^I��ٖ��?"TUG����6��蟜mh@F�m�|���׹%ܲK��&�����1Q���CV�~)8�ѨĎ F�Grͅ��V8l���0@���{�?�,��E�N86I���lCTh��)g����)�Ր��l��#Њ7 '� �\?��o��t�p��)	.��a�MZ��9����C�j����ak+E�;��Y�K&��У�
�09������tLIGI���G�;�� B.����A?Cf@b�޸@��A`�;ԝˣ�
�W�M0w��*x����-=���q�Pr�^��
�b�\O�����ޔ�{3L�E"�^�BT�)$����~ʉ<�6;�p��toȏj������Ŕ�q�NVz�������
���-�Ղy�H�m#�;��2�8z��f|Ǭ��$y5O�1�r|BO9�V2���%8�I>�9��EW�;�������gxN���Ct�-~�O��	�1�	������	@b4Y҂��`kd�9b�?�D~c�7�s#�j~f��f2p�Ξ-�A  ��🉠���)JN��y!#'w���w��k�^^=�2�]F��HH�R,C Y\��X�D�z���9x�6)s.��l�~�uvS�u�;�Q9����aG	�_��ʲ��H�%�V$|�p�qf��d�g���@���~-<�H�uq�D%�7���6g�����s �(�?t�I3�V3��\��Ky��[s��%�F�ʠ�x���]ջG�,( _�h�ȯbR�Sg$��Da�f=E���K������uϮ`8�pyF�/��P$߲�#��}�~Y,z��xB���Ms���'4V�N���9Z���&�>���5����x: ��*ge?x�"��7��|Up%y�
�[�9HtrE��]n�LUq~Q|��'��6��D��{���~��ԪTT��R�Y�i5��"�O�<
2v����]�_wWQs�i�{rv�RE'%�(���E`j�?�9Y�O͓���)�9U�`�������N�|�]��*ZO��z,e&␥� �: �C���t\3�ʴ��<�{
�!Ȣʺ���PMU]�x}�r��Y�y_%����t�Y�[v	�UX/u�r��I�.��ժ����Ѫ9G#f�uMA /A�П"���T����$g�.��hř*�x�j���Ò4n�m$ }[�t��+�6�%*��շb���o
)�2�W��6���gp9��q�	z?dgЯ�����\��0]n#��,ڮ/�����+�N�p�7�Z�L�m^yrun˶Yg�+Ic�\-�)7���wь���p�̖)Z��E��yK�A!�7�i(�Z���i9NUܼr��������9�p���a'_]���a��ܧjw +M�Ϝ���q#{��q���7�-j�}�F�UG3�u�5y�+@ǐ��L�q�n?�0ȗ8Z�ӌ��kV�݃\���ҷ�YÕ�����"i���X;!�BMjI\�ω�\9����� 
!�^��*
{�W��	����<�W�0����x�3o���t��㚮�W��	SQp�]Ĩ�]!`࢏���>A�G��?J�����n�V�h\���c�}����Oֵ��f�v�j���^
s�s�9�3q�$ZO�6�l_����ū��,��C��J�λ��-l�@3	=+�kf�1����b,���J���y�I7�I.�g�_�AZ�q������E���|�Z����C�Ξ�ʽ�Nm��Ub.G�'��?�����}qR�����p�����u;�&Е��+h�ͦ�Bw/ōj�GF-�к�[�6Z+!G5��������̝��L�N��Թs3�HLp>V�J���\7��Q���Z��-7�,��V���\�?W�)���Z	`�9�!%w��E��N���$�0��5PG
�V�H�Rl�Z��e���i&����}�FX��z��ޚ���������)ɦ�7hqtb�OH����n��j�X��#е�T���E�ڢ�W#��eW�8����>�RV�Jl݊�4�'����Iѵ�Ľ���i]�y�_eP.ъ���s���ua�J�����]{���w��֍���x�[�K\��m�'jʙ���΅��K���V|�+DZ� 曻�� #���q" *	�b3cӐ�)���w��� ;��N9���=�]!iY;w��	������ۛ=�ɠ���k�x=w�:����~�S����`��	����$'��g Ɍ�[�����
�e={�F\/ʌ�L����{ P�S�W�� di��ߪ~j�.��p@��</��y#%3�f��sٷH�tIkRȼ���<�p���Qf%8
��
����2'9��X,,���IB�w�lâ����1F3B�p⅊7�)�&�Bz�m�?�U��FGMe25�Kų���@�m�F|�$��^$�y�k�'���2f2d41F;4Ri��=�_=�z-�ݠc�K��)�����zN�^	ʄ/�ο+���L�e�\7��=�Z�i`Syk�������뎏�^\�u(���f\ǫ�8���f����l)�v���f{?�,]�`}�h�G��79=�t�Hw��iH7(�?�t����ڄ�؋)��TP��򣢟�̺�F0����(�Ny=�C�b)mpo,�?�5��1|9�4�0q�h9x�^�{+�	.�/!p��[R\��C�F�ߧ[�a�?VfT�ϬL��>;!����_���~}��(���[r7	W;=�H���٧)Vɱ�n��
�:�Έ��H�o������ ��U��h��<H.��$e%�pR����I�\.�`��)y�>/I��|3�W�a����*���9�C��f����-z���?��/O�%�V��ˣ�J
I�R����} x�����0��G�%�G�'���o/���*����;E,^��띉2
n��4]�/���E{ՄL"��O{S'�ԷޗAB*��C���U_svac
˚`�S����#�/r�[;�S|�|���ʩf4���N^�U��M�)���X�z��t��	�@q*7��%p�H7�TS>�26���<�-9�(=	ܻ�+U�'E�W� 1o��+�:�����R�w�jv�������r�Nn<д��1�2��py��g��1��i�E��{���̶i�M&w�.9@���~߱T���OI���v9a[<��'1�fh�x�B �_���X��J�
�}2>َ�Գ��� bx��W��ǧ/�.��ߙī���4L�1����dq�Ç�ϻ뇫O����@�665����9����ihT:
�[*��7�m{ȼ�y��{8�c�Η��$B�t}G��Ln��-���B��A��|4���`��35hH��&P�>������Юx8#��V����m�a FĲ��"��A��#Ii�p�Vd�o������p�5�C�M�ȭ���r�Q�pk����P�j�n`���v����I��T�K��vT�a`�uɋ �f���U~��@�ecjf>s<�Yl�F�L^���߮��j	�=/��oo:p�=���L����!�M����g��0�Ѕsx7��k�-�S \��Ŋ�qb���A��=7J�/�����ȣ�?"\`���r�p)ܬ��N��{V	�*��Q�ȷ�ܕ�Ȼby�?|�@�'~��:�@>�_���kD����N_<e�����o���1�\�Q`8]�z��'����l  �:w��;F5�!=0(U�ZME������*���w���5���?�+��/�oU�*Z~��x�J��΋Rƫ-�@�M�F�CZ�FyrJ�Kx�v�S�Řʆ.���G���s6��Fk��'��k�s⎹�Ϛ�+�gE��c���y�����	�DE���(e��oZ!������+����['�D`�+M�Ƴf/�˲��0~�v\�	��4sL�r��� ��W&�9��{��w��DEcY+va�D4B�1�y��՚!wi��E��b$�4EP�b���S�vo>�T/����CD#|���_��
g��OEn��ݶT�C	IuJ��˰��/-O�O5LL�r�����N�壞��`cpY�����H/[)�2�{#Sf��n�uqpz����Ť�Y��O���="�ܝq�hq�_�#�42�~Cފ�B97�KK�nj=�]bCke�gR�L���s�=����{�~Ǳ�;>_)S��e��G��+Qq���%����7�_@9z���>���323� ᶦ�:�M�����K�+�Ͳ����@3�܅��g�����6��/P��:M2	D�,�Q�[�������ܪM)��$(��)�N�j9�=�.۩�E_�1+�}Ǉ+k
��zgh�q��$����'�� ,��L��?�B���D�N����ꬭ,�	��MS��	�Rs砻��I��_���j>#VR����3�R�}n�:����~ֵ᧴?�߶���2v�B��x�o�ױP��Ū��|{�oc����菌V�>���brh�V�L_��,�h��%����*Ȩy��_tR��=��,��ťb^?�ֽwχ��&u���(֨1観�\5��������ZOO(<�GH܊�d#-�h�f���r���Q7Xڴ�g�M$�>�4Z�ᧅ�0����22��i�bQ[��r �-�������M@�W��9�q�� �qWN��v�ٝ�D����BW�2�d�5�2w�tLfm�Fw����M�O�����@ܞ"�j���b毞�u����� ��9%I��悁$a<�I/H�X�U�!{�����!�E��D��2k��J�d�Wo3/x�X�Gj�7��:��O�a�!nB;'�D҂���ۅ�X�q�ny��.�pM�{��|��U��2���G������t���J*#�Jk�Yl��rx��j{��P��Yi^Tne�<���3�J?E�Fm�S����X�j��3�_��2����Wk2mZm�A�u�{Phyeŭ6���$[��-��ltɅ�+6w�H`����j���ȝP��h.�%;b�FYT�E�|zr��Mwx$��*�Nٸmm�<AP �I���r�yc�8rjl���v�z���4,��%�&jP�K�KM�m�S
�aSp���'�mL�u��4-fo���
M2ӳ��j�h9�y��`�K&�<� �X-����ǜ����ѲCz�r0��8���ӯ}�p6N�*ȴ�+}���@�Ld6��ޭp���vΓ�����5�+��G�!̈́�ߗM���*���F���� �Er-�6U������ox���ҥ�Uڽ�uF��yўL�n�y]:1�f������2Aat�T�j�E��D:��fa�%�uیgWߐ���qhN�l�9��x�B�
�h?�O�H;nB9�e����$��Z�d�T=���P���`n�!��/ɸ��D@��C?��� s�,����qXY`~������)�����֦���?G��1����K�Oсاh�X�����k�Ui�B��@p��5��Z�C�o�k'_)Z�hT��QTI��S���n�ܸ��Ș�;tϸf^���t��u���Q��e���Ha�W��j%����ۦ� �<٤\��dL�޴�uxa }篧��ۈD��y�˰v��i�[�oL��yd;N*`�ψ�������#�����t�rO��ô����>����m���_�HT��9w���sL=d{@9�A�I �Ґ���-s�z����]� Y�n��D��K^{��?]S �=������z��`�ĶḶ!�x-������#��Qd���a�Lr�j����pi��t�df!�C�N@��Q�wYp�D�$-g�K���cp�=FY����O�J��IbķI���`�/���k[ә��_�T3
��.��k�7Lc�-�v�N<R~넣 ���|S�us3���y?�����\��|�S)�*�fOn8ef���`�J�����c�XDf���.��~ǩ���&p��6 ~3N���I�I��뀝�ɤ�;��@ƚǤ���&kG�~Z���Yw�SW����:	�7��a/3�!޴GH��� ��%�/v��iva;�i�+�}>��F0C�����ȋ9�3ᱱ`A�	$N�����z�A�R�a�YhG(��3v�z����T�nVLm�*�	��%·k�s�4�@y�F�e��!�d����FD �w�������l��h���	&�vĕ�;��VKHj�k|�8T��coq.!�kRȤ�^�\Rڧ]�p�ʹ�;=ΔW��YMLn��w���p[��cB�����0�m��Zvw=�Z���u%��Xܼ��-~�"�������e����TV���#f�(������*hbff�Vn3�D�>b�!�k5"|)�����he-#T���������rY�!�˶Y0�&�0��ۜ�-B�+Q��l��>��s3�V�YUbz��vx�i5�[Zh�#	;k��Y3~l������k����^�6�M����sX��og,U�<���ӟ��n9��T� W���E�D����msl��|���,P(�� W�����A����4h�,��R�V^��+?�P��X�|�$�-��X�dH�8�y����Fm��N����SS�&�ߟ,퐏3W��M����x��Ǻ�}�`���b}��cG_e��4��X���"�M6�L���1wPQs�^��{H�V>$�f@��" �v"_����f�$Ԣ��g�i��!�Ixv߱�9�������6Bl����,[��/.2Q�)v�N��0���sJ �MAd�3u+�rA�0_E���<���\t6�Y�y|���/��s��T��H~�Yq-Z ��/~��ߊ��>�s_{qʨQ��%��|H;��A6�`���2��eљ+(��D����D�t@yk9,q�Pt�-�s��D����}�Ԡ�����.�L�ϥi�Zy��զxY������[=�aԁ� M+���D�D��[��=5ox�^�4ͤ�����l��eb��o��^0��]G!��V%EE_!��<6Usdg_�[<�ݺ� �j�cT~�}�:����8��HV��8��k�M�8#���_=U1�	A�Y�Q(JT�b
�s��������;轒�!�v�˧e�m��u�H���i�-��R�8hC_�s��AAo�v�(��99�lO��-���[q�<4q������Ϛ�3�X��PQ�#S��tu�)OE>��=4�@Zl�>3l�Y���@����cmE׆�{i�>�ո<H.�L�C��v�m�)wp �0��bF8����� P�����7��K�1EU5��7([�8I���E�gG+<��{}�Ӣ_�ږ-�[�m�������p���F���;�4���̶蚖�N0pd��`� �ǋ��P"NZ��ޑf�qM��ď�se��ަ���y��&=��x��.3�����r�>���{�AtЛ� !!��
�Y�S��x���''�,��>g�Fu�a5�!�2C���&x/e���輏��8_<D�uG�=�x��}�[��,]�{�ǀ�_a���Lf��#�&�xu�)`x�qP�0�˗�y��C�KTIz����j�͸�0������9��9y᠓�B!�k�K|�4���"���^���<V$P���W`λ6�|A΅\�f�� .�jV&K���_����9�9����#N�)_��6��|����u��{�h{� �j`J/?˛/d�q�S躊�����1�����۶$:�Vݝ9�f�(�$�bnx�P7�<�T��t~G�r��M�/�Tk�kђ���m;��n���~Kf x��O�2QTpX��\�oû�$��O�0zjQ+~}K�)���I��:Ã�ae�mg\�Efœ�i�3�j<�(PS�6�U�����rT�m(�w�-����-;���<�>fN�޼6��9�M���󅋋�۹X(+�n��βû@Μ����P���:��8�`L�[�� ��T�g��m*����*�E�i�覍���C i�g�o�$������k�x�\`m��S�h�#�P��т!���`?�=221k��\�1�oZ��n��C��Q�'G$�W�$�I��oPD�׹De�/�v��'���%��B��ү7�P1k��xhRF��J���}` x�ܴB��%ede�����7띄�$�Rѷ��ф{�B[~5�Y����(�gUm�=/ٖǲr������{�
�%�ſx>�R�b�"��y� �A���=ʬa�&���!�hM�io	
tpȧ.:���q˺�L�-?h.[�6�$\ś����GG3��#1��Ɠc�Nl���uDE�����=UM�kә��"A�
so�T� 愢J�l�� U���"��❥�ܞ?7�,>壱#��|H��r聱&'{ج��[��%�7��f`ΥD�u֡�`�����w��e�{G��t��g"WB~x���H��D�����Xj�t� A���<�u���)��;��4[=���}�-���>���3��1�T@h���!k<�!Y�G����ͽ��8�&o$P��=��% KzŦ�U󃺏:r�l�ܻyq���f�\~tF���{�n�c��뺔u�Q���0���%_$Q�f5�a�ڔ7�#]3I�}�#w���]�oj��cB�}� �������~���ݥ5 ��$y�%�V%ys�u���7�~Tة��r�/�(X�5�����HC2z-?	���νү�����,���U����M�����i�g�Ґ��ۊ��6fj--���U�?Z�0���+֯�����yi��<;�V,Y�;�\�N��孑�Ht��?K�����5�~��W(�����ż�r�S~" q�_sw��(�=��5�>]����jd�2nޫ�e}��*��/��y�6��3J�1�~=77Fˬ�.�A�}�f}���.�1x���դ����'��6�ܝK��3,h0���d�G�K�Y��
��F�3�v�K)Is�c����S�����Fe���&Md��b��-��j�niI\�̼3�r�뱄F+Oq�ܖS�N�#���m���T?��3���le��D�`��!�/�#el%� ����afw��0���EV�ԹPl�
;��6�H�l�d��������,T�5����­Ɂ@�۪}�o՝��X��a����2푯�������>���m17q3͌�I��k�w4"�:���d�	��!s�����?e5��\|W�,	<�Cp�|�@pwwwYl��[��-�������w�}����TwW�Twf�)X�W<�v]�dw�]^�M��Hy���)�p�^��~	�XWݔvu��0>� K:r�3]��-�dڽj�(i���߱Q�tx�F��w��.��y�hX�V*-5���i>(ͱ�p��&(���"4*'�ņ0��(I�܃\N7[+��b54���zXr���j��?�k��8f����X���X�N�_}��M�'���t4#'��;r��k��Kђ��Xfc	�u��ل �xIGG�0E�3���>87�xޞ<��,����� Ҿ����Cnֶ2Vχ�V�W��6zp�t�:M��x,#
������k��_��!8�B�J���\f�٘�Ji~:��C�B�Z��}��-Dh۷]����x��߅n0��"�>��>t�b��TQ��@�� ���(�cT�Bs>�E�/۫I��2H�2���D�N>%ğF�ԇ���Z��\��t�rt�&`Ol���32��� Y�-�נ��0��(6p��nU�Z����&����#41N��r�T1�ʱ*J&t:߃��eH���κ1��s�joƦ���#d��%�=�<U8�������(�۲����yP��v(���,-,�^��A5 )�o��{D����6����q��;=�ΚJ�����=,�ܗ��y� W!B,,�C���Ws��
7�#�Kշ!vҢ�3D,EzS�8�u�]C�]�y;۞�a�w�L �k�,�*��-��M�{< V�|C�=z&]Ys���`y����,1u<#%���|�M5�J��d�m7ޘ�C=E`ٗ��8�%�@�V{�WX�l�fP�W��w5)_��
m"��H�~�װ�~U���s)>��QU�N��ew��=Vi�9.б6|��6�[�{!����r^�N�Q�t�%0���;6\FvLO��kZ29����(����ui��N�m(�h�\���K<����jj#ĠP�~}/���!5�v,�})K㝍�1�픔����kC�T���5�$B71X���W�>�� }�뼻G͈4���i�W	mC�W�uJVL��L�{��u=8 �����	�i�hh���}���H��_U3m�WǍ.����2���߼�tP�n�05(b�mI��_������xC��n8_��ˈ��|�`�V��-P��d�y�I3�K�HWUU�#�Ƴ�n�U��9qHO��ћ{�1gA�
�H��h�J�:�|x�V$�]�E�|3�&�3���-��`�
I����^Iw�<�b�*����1s1g0iK����)��k�+����":(��ʺ�{���DV�������,�$�������6�(ߋ���7�V��zVf�� &v�6� 밅[&0�Nk�/���c�v_U��)�\u�(N�|3uR�_�|��FT$w:�l�6��8�����#�=.B��7u�4�Q3?S�F'n�r& �?O� ̨w{�6�r]Տ�v�k��%���6:iҳ�/#.;B�K'��������.���T�L;���+niUM����g���"�޵<G9:Ɔ�I����j\�a�"���9�(���1��f���y��Bx�庖�Am��R�.���ݔ�a�37[��i6�ӊ`�6H����2�L+���E����y��ۦS�3��1'��K��)X����|�v��5hXEwn�$���ZǪp�%^J��$ �N[ȥo�I��V��}L���P��	?��j�O��s�?��N��=��������*���+�lb��I����B�/��a?|63����Q��:�M,���q(ǟoc�]�q��^V�nz��B���Ӿ�k��p�5�1���#3�N(������<4����k0�Aa}���G�O���_��ȁ��[���ҒhӒv����`C��N@�ْ�3�8t ��ջ��C�y�E��$V��{O��n��z�ׄ�<$5�B�`����őy׷&W�o��\b��e�k�̼���s�9GZDESMٲ������S�[1 ����2ZK+k�8Ľ�$��3�O��yD�+kx�����:���1��i�\}����483���]�E�w�[ -�e��q?�3��$w��ŸE�=���>���[Qâ��%  xȏqN0�o"���H~Hf�x��;��5S9���$0���ʱS1�.">��o�g�4w�>������k�/7 �4�L��5]��9<��Z����C��B�=��Y$/�Ab��ݜ,4���Kf��?7�#.��-�I��=�U��|�+�5j~~�؅$I��l8{����QɈ�ly���d��+|^��ru�"K��#ml�+g�?G�����ʄ�߿�E����# �p> h�?�U��pm��U��&�'���3�ٞ+�㛾ԍ���t�/68)� �X���1��N�Y��0�o���HͤҫZ8 �!�F|L�����߸&������Ja����&�x"קf��ٚ1].����	쬹]��9�,c��.��9��ՙK�?��7�[K;���w�=kY_$�ޞ`�z�_��C�5�4^i`�Q�Ja�f��`�cf2f ��e	d1���Θ��a;`�U_��Ȥ��y#��"��RM�u�����ݰ�L��
��0>�qE�]Խ�X$(]�m%���R�]"wXc�H�D�ͼ�F�ٙ��*ծ���v"����ZHP\�GGF8w=\�u7]�6�j3&8�͖4]笀�႙*�=1sS�.X�9��(F��V.�=H�i���]榋LDӶ->.��bI9]��x�'���u&��1HH�����<=�t0A�o%�j]#[���hm9H�;�촚m�lh�A77�*p�[��~\�a㡋<�r�:Z0O,I�����}?��S���$��p�y�|h��UU��97+��������� .��5����H��^=��h
� ����j�������1 t�J�d��G_���8O����n�}��Cb���l���d����z���nx8&����b����y�t�}����{�{�EӶ^���b�����Z�I:ͳ�� �,�䇊�۴��8#��,����7A��nש��Q؜�͂ށbus�|9!4��\x�ý�bqW� �039�)�Ɉ�X�#���iF�������^6�Y7�K��Gk���|^Ams,��Dv�Z����t��ó3�c�z[E�Y`knA��/���or�<����T�yq�i����|2���`5^]#�T#�k ��z��/��=��P��Ah}@�du��K&%-�JH����r��VG}�ܣ��7 i���p<6�O�GYY0��b(���Q�R۽+���)�X�(�
?W�XK�������34!�a1Y�>�G{�th��$��?}Э;Q�k(����4���t�=��q��̳Ҙ�cL�5����!Vmk�yst}ai�2�w��֠�!��|G���B1�+���/]��<Q&o�S�s7���|Aa^mA����|6}���md qt�ef�wd��i;겉l�Eӿ�qY&���!e3Lz���J_	C	��wlaM_�ܹ~6��`=z��_y\�`3�[t)�T��M~��"��:����!w�o��j[�z���=^mvV���>>�c��_nX\]y���������y�(�h&m׬.����g����:c���G3p~:�CLsk��ի��������]�u��R��FR��w.�X{6��74g�* ��פ����Վ���R��0�3��{��<�au2F�3�`G�􅃒���(6[�Y�m������ڍ#z�Ӹʽy������D
M MY���#t;� ��D���임���r�<���3KZa��ڻI���Ƕ���J���,�sI��U!_��ܕ�h�p����k���}�o%�Pc�$��<�4��rxE��f��Y��単�W���[�R�/��Q�;�GE��&����w�����?��	x�u�IM��gXD�7	�g��ZF;6���7��ۖ2��������b[yT��H��@M=��N=�mEt���&��<��c���ϯF�fJD�\�-��f	�v©��$qV�	���n?9����V:�)^k`��(lnN�"��,k}h�w[����������7 �.`@t��q�dN3��;�Ɉ�h�a��j�{��j��2�O�:g8���;MpS�B,��.����z��M�� �.%�P5��ƑA#����=%ñ��n���׻	mݾd��ρ^��9L��@�6���Ok�U0�Jo��N��#��L����+ߠ3��^Z¢�"X�F��iiR��q*;#v����$�H�&0����Xt[� �o�%[0i;����O�<�l]��v+��t� Y����,�>$�՟%!ҁ~"qE+Ǝ#�R�y+d՛[���o4���0��.@�X�E5:q�L���ը�}���yؕ�w`Wt ��,V��q?�9��ll��N�/)T�� �������������p|�����$�<��ۋ;�2ccb�=�.�.�b�T
J!�<7����$�������
�4�߻���5�e��h�Εh��n=Zdi2����xME���|�h�_̧4�Y�5��\p[��촩�����d�q���ʧ��V˧;��h�ڼs���(�������E�+ѥ�_�U{J18�91TY��3���\&�{䦱V�Ҭ/ﰙ��1Lhy{�[�<}f�0C�����f��ݦ�G��:	9u,�w�����(�w';���H��ר(����٬�ی*`��ń��BLOa�}���m*��(�Zy�W��,t�F�!?��mK�;9�{;��;Ok��������2�+(@}�`�p��?�E�4�����)���.��y;O\���D��+��~]p9:|k �a�C����5�"���n+�G�����5���F��uq��f��Ԓ-�4��-ߟ���������%]���p�a>cb"��N%����Q����%�,
h��"h�OCi���q�v��e�4%�h�`^w �oZ!�R;c�cfBN'.�}�֢P��=�A�t���ɋ�7��VU"ژ�@�D�lñQ�e�B�v&
�'B��.u�=��{!�X�|$���BAq���~����{�]�U��-�UC���va���?��j�L
�T�O>����&�@��� R��5'{[[E!�d�N͓�v gc+ȡ
�4�?��̡AE���ԗo���䒛��Onk���,�1�y��Rd,H�o9(��~Z��L	��#����V&B�w^��X��p���m5x.$�!)B�)��K��z�~�9��P �އ{k�"\�	�]�`)�ؽgW�˷��?=@�2�d�v�Ӡ�%��po��C1�ţ>��T�"��I_R�G�7�8X�~��Gůq�s�r��!�p��ĭl�;��� �]���a�ϒtB*���%ߎ�y?��my�#8)�����M�i	Ha��*�t�֤Y�3�_Ya�ZW���opUM��DI�m�l���8�}�6#��8d'ɩմc!�S`��얚��U�x����W᠓��6�E�T�o�ռ���늉����p3�jF4sC��ǆK�2q��֎�]��$X�����aIn����o���5�u���=)��?@����&B?W�������O�r��''-J�;� ��-!���퉍n����Q(����$�~Oi���0,��us<^�?ՐU��\��;�����;XbBmcA��F����"�
�o=���_���S��y���f�"�]";�n�k��<ob_i��\�"ݲ��ɦ�:�����b,a⭕�e<�&ǒ Ц����ڟ�&�Gf����BX�@�M��4�Lvh������[E�!Ͳ���nwn�9 ��-���J�b�r���,}[3��������9p�-)P�����X����Զ~���1�f�YSwC���_@�	���~�Y�b�m�3𑹻O��C�"��a�\H$Zo��g��y!��4jy�_��җY�	�=��ip&<ICF���i�֛ 7����~l#������V}$CU�_=�ͻ���j� �"J��B j��n�x���._x�@w�Z�	y/���v�XZ,��o�p�u�P��Wf�2f�%RRb�l�ʏ��(�����n��Cx�f���v�'�&TKR,M�d��*���tTU��v�g��]����ȤG�ͬK����%��w���I˂�2��6_ߧ��V����V�J�=MS�q�o�o���# �[����_	-m&�}𭊖���%"�q�F�U\A�4.�w�	X�_Înoή��q��)+���s�Q�(�b������q
��\|��g'��lφa�����JOu���]�#��3�{Z�E�Y)ѥ�CJ'���*��k�^�ZH�
e��"���}�q^G����E ���AZ�+�NՂ��!��m�X�$��:� �������$4鑵u���E���2����~U���un.�"D�%��WyD���w^e�0t����;�H?���zN�����y�]<���z�q)i��,�~R *�l������.��0G۶6��&����9��H*�M������]��]���)�6��M���{�LHd��`3�o���P޽�P%O������x~���������;�ݓ
>�j�ϸ��>D�Eb��
��zL����x�6��٩��=�bǩ�s��;�ȉ�@^$8�LҜu��$%���$�	,���J����!��$�]M�T��0��7��4�2����!ҿ����!um\*��+�5���;��7]&�G�r'�Ru�^$UF`ە��߇���M.�x������]�6A��n>��/�b�zZmvv~�f���+v~4Z�sm�Vc�U��XlE���>�yv����Ȭ[;��:F�I�jiGc��4s���3�b!EYj�͖��	�sߙ�X�f��15SF��Ci��Bd��5�C��N�UГ�{�_@�p*d2�m�����<.�z<����Կ�w�W��fY@Rdz��b�J5��C��^�f�7{���	h#�n�WIJ��@���ú*�w����x�u{�v����������z���^[+�ؼ�wok���C��⌾]��NG*�T���������@`��rmJ/&}^�ƀ\̬��bՓ�b�3�����YIj�2��F�:�^G���9��:��j&����J���{s?cD�P����@�ҹ ��O[E���������z��t��c�=RRo�8B�a�
Gz�ܷ���eJQ��U{��e4���:t�w��{�`��u�<7^������J��f��rm�iU��{��2}Al�����Z���2N�H`m���p6;�}[�t��k5�t0���[c�	,[�F����� �]=��67?]��yh�[��'q-�\D�j�;�b]�NOUXqL��
4R�˭�f������:�KE����J(Pb�KS��=oQnl�>��K(�RJ���=�U�Sm�����xI��ڮ�)�,������K����Lj��-�C�c����b�(I�Gݻ�M�r�w�mt���K]�9x��-w�Y^{�j��G�,W	=&'M�ws-�H��b�N�u��#SM�#Gkzp��3�"��oSqoI�$�Jktx�q�pr�sNDI����Ie�:#D~n[�}A���~EZ~R]���j��^�q�9j�_t����h6� \���I���%��YUy�8�P��u��w]�0����@����P1g��Y�kE�ƛ�"���86��?�ΐ�k�y>�͘�Su���gד��Xҵ���)�����鑓�P`��A������Z͜��Iٺ#�u��I*��w[��P��
*�3$�U'l!&\�9��q5N��q��f����*&E=a�Ȧ��z�L��`�Sa~�N	�Y2��9S�2VnO:c���0eC�Ev���3m��m� �"���,0bۙ��O�s5"7��/E���P�|d1V�wG���9-��][$?���k�aˇ�v]��=n���0�QY���K\��d .���F�{�9��&f��Zj���FSg�:�n���̆#M����Gl�Ā�!�j��[��ԡ":?G��wPlo����P�\ZH�VvX��X��\�w|Щ�o1lч=)�r�ϝ93�ɻWIl�/O��j��J������ �Ɩ�R/��jF����uf�` ��Z��,qG>�qaћS���txԕ/٢��56�~���&&[J�7�cՓ�0�WbZ����k���V�!B�?����$�t�[,�*�2�OVW�箩[
G/!�H�h�����U8�@FR��&:g���J`�&Bg�x#��9���G@�����0���ȨY�5��yj]R���}ʯ�m��R���s�_��7y�N�@0���kFl��n�d�e�v���Gٳ��z��{��=��R@�����rp���7!#�����Z��i+�`.+r[7/d�t�{҂���Z�7E@��	n\���x"p{k\c<m���-�������y�G����'������	� i�Dlǌ�ܹʙ)R��0�
e���ϔ�ې���k�3����%5��4Wi�U�H�]c{z���
"D/w��JX�2۸v�㙞c��ϫX@��p7\t[���@��0�����ė9��e��`�z��eZ'��NT�/v��Y��Ab%�&uJ����q��+5���]�<�`�?Q�CQ�|�ˊO޴��������-�Dc�ܐ��)M�;��<�*����>�r��^$�˳�X5@�j��IZ�A]Bv���[dB�)�Fu�s�kO�`�q��֬HnA��N����H7,��b�#���� ���6�Ȧ��?j<U\A k1E��.f����J�i���%�2��pB����'�L�����Z�ӿ�^,�Ws�X�g�ln9	J�w,���0F��h�1f�.v��eQ���%��ݑH7�&�f_�1�����VX�A׫��ô۵u�1-�-��DR�W3�yo)P]��C����o�_NYo��U+f�����J(�$�* *�,�����4�%��R@�[����4[3��l���{�ڪ��/I�?���}�H`x[�L
�L{sR+_N�"i;�7�jrLz���u��ϸ�j��I;�S�p��~o,�3�<u����tֆ���{T���o�X�{G��+�*A�9�Ñ���F)�
Y��@!=SG.�Pm<_�;�����d�wC^а!8q4m}"����fQ��ah�&�P��o�T,G���⣡�a���P�g�o����!�u�7���U�wԑ
����Lk�i�N�l#�H� ���Mn���i2*�g���gJ������HE��fc�V�s<R}����s�s��ֵY��� ŗ����#�^�� �b���0�Ĳ�:%�'NFߴrS��m8}Ȑak����
�:��r/>���UH �"����[������g��>���A�<�z���z�p�'����̖�1b�����m` �>�t���c��"pOl�cY���,~r_�O��Iw/G'�z���yK�5��:�)�=Fc�!Qak7b��*�X=��X��Xa8h/?	�R��#F=ǎ�쉟J��h���9�,�
��m���踻?+ʺ}�y�ﵷ���Z�b�=��4'��:�z�<��׀K^U鮢���?JIOg����:�U�J� �7�d�/ݦ%{���h�[S�?��_BNڠ��(%A����".a�[DL���).�h���l�1�,W�<��J���|�ؘ�>Fa]�y�+J����F��&)��K«���I�0��+&-a�b�K��n���>���ޜ|�ש�p�Gl.��d��;��besW:�1t�H�Ek�nZ�d@b���/�%vp��,�P�Q���,h�&9�b/�HV�#S2�7@�v�������~0^Ե?�CX�c��<�_ټR�!1~=y��I��b���(��eo�z*4���G�����߿�?~�B��G?�S�8>���#��YV��/U��s��zOx�?���ּy����w�Z>=�}P�KC�t��,%����l0����i�"�-1��ε�D�-�ϒ�o蠨��"�81�O+�gkj�����P��Y�!�!�{_�ڰ~��$�b������Ţ��]�m�tV>�BA�g"� �'n=ȿ!)�%e?!Qj��U2�y*jO�Z�(K�������C1
GIt,�N����#�kh/Ć�Ӽ�N@&���o�<R��{%�*��򤉱�Ur�Fk�|���4�6Xyh�`������[��P@��C�$��h��#t�H��m$��l4ArJ���ڐ����\]c!����'&����{���^	OV�T(O���G�������Ě�I��~��ç�%_���gT�i���+iQG�ҋ!�J���[^�Q�T�G�c���4�QI�9��9����ol_}��0��ъ���#'x�IaRQ��kv&��x@3%>ց	u��x���8�����LO��!|w�m�}�"O�z�D�r6!÷..�I�����xQ���5v�>��] �}}��ιOW����=/;���/�_R�W�L͇k�}S͇G��aj�5����ħ��4A�uw���m
��1`9H�JP4�b`�ذ�X�aFq<oHU���2��.W�s�C����1��W�ֶ*�ӌ+�V�Y#���Wc5�����v��#jZ}�D��jۤ�ul4���W�n��z,����B�壙\z�pW�l�	��H���z`�^}�~o��^�?7��}�>@��~����A{\��l�dVq�F�+;7 �D0ASp����+���S-���R��n�.K�G��g�=�`�st�q�rZs�l5mQ3����R���6}� �j=3v��_Ӏ�T�)<sUX���7�>�L_��]k�Ѧ�%D�|�0N�Uo�7h�S\�;5�9����uq.~ǧ�I����#3�Eܾ���J�E��<��L����,͜��He���j*rvÀ����؂���%�x JG=���O����K����F�DaS���X[��4q�0ߠ��օ�����+���F]���_�W�L�\�F�%�<��嚽�G�uܸ��^BR"WM%�%n_^&��V���̄9�_�z�\t=1�m7n~]/@�<3o�U�� �`s�}��nn�N�>�A��P����?�XOf���V��G�=����n�eQ(�z�vG|z���0� �����zA���$˶��輸��o��i��"�c|��gԔ��:�%~
D��R�g�а�lcW \:�<���@�M5�yyM_#��P�����#�Ņ��� ,j�E��eǙ���B3kD2����8����u�;�@Ʀ���m=sB�MI98�_��d讉G�w-�*!��,Ho�ZG/*��ي8+���w{�̿?�;*���w��"qw%��%"?��m|`k�>���l�$`�x���-�Ͱ���{e�����hx8��٭�~�'���#c���f����
�v�5�h7���F��֯/D�zZj����!���x�Z/����[��2_>c:�hH���n4�P��!S��|a���Y�\�{����������"D��+���f�3\D`ǯ�o9�8Pɍ.cU 6��_��D�����g����Mu�7��d�%�,1�-g$��Hm*1��^�C���G����o����P=߯?��?�I����x�P�P�s���B�����p�~��Y?z"�Q���.�3�j�ۊ�UH2���?�G�M�*��2v/P�?�*l�.o
��uwx֐����|�w�w�6��p}��"����b_� ��_cK���am�d�G��R]wSg�[�������N�ݣV�ŸJ1��W+�i1������QR_;��W��ru��.��_,mz�O�v�+^�g�����M�Om�KO��n'�>+����Шi?�:�8P��4���u�{K����%M���V�yӱ0eIv�lMv0�n}\�*��C��)ה�:I�g�
Nm�'t��ˉYn����^��H�[ V�*��-����&.Q��nB�#�u���7��؝&cy@;�E����:s%6&���sw'�i^uN�d�陿�S����x�6�����|ơ'"��T�w� ����׀x0�k��0��[
,�{� �&���.�;.��>��=I�C`st)HЬ��c����";���.,,ٷr{/�j�!��D��W(��`9���V��FW+&I����V�w�Z�O�ONGx����]E��E�_�c#�E���\3���Vר2A[/�����ε~|}B�D�>v��P�*�j��2x�3k�Ø,�7�9����z���M��{H��a���/5ZcjQ���'ޔ�#T��J�cun���w�(��h-��
�u�;o�,ٜ�qP�Τƫ8n-�.T�;d��%$o�x) �"��/>w1̸'���n��9�+v�n�>��\�"WY�P�rD���m�R�.f3!�'�3/�ۋ_�\'��c k��8&{�t{z<9<<����P��r�ǃ���$�<*�[^��Tt#��0oQ�bd+>ط�^n�����ݷY�o�����e>\i�&)�k�m�\%��׏/ϋգ����in>�`YmN{�휝LN���zޗ0=��ʦ(��l�b�8��IdEƟ�j9~�[�(G������i5v+��'-ip��}��A�v3|e��4�=�_����}�E9�O�{PR��.����Mw��'�j2���oLӲBc�
�Vƶٍ�]�+h�ͥ�1�;[�$�[^<�k����M
�1(���44����-�1껵d��Ο��M�ݗ�'W����)��֜} �C�ệK��-dj��O��퇩*6�9_�??o:����R���T�ӕ����^y�{nX�2���9��YA�n#D g�ޮ���ɴ�i�1�(�o��~���T��c%�u h�H���Ϛ��4�e����]<�lR���������Q����|3W
x�7K�e#�Q��B�w΍R�xo�M��Yil�[���E�q�����l^N2�h�g���}�*A2<�a]1_���.�P�ҲX�T���Q�E2���*OC��Py�����������5W̲-�%V�S�1#�9�tN����-�PT�F�F�5��O��T*��JΆ9
b��0Z�A~��v�k@�9�`e��Y֦��:�	;rAaH��S�(ن��Y��z�|"2������i1�͞�� V:�8�ȟZW�9{�T�Ҥ�l��x��2o�rG��O ���28�i�k���-dKe�A�8�Z��3�/s�c�s�����!�	�p������	x�4�uj��s�"^��o��°W]x�7�BQVOe�k�8��"�I��%:�: ��__`O�w6NK+��5��}k-4Qgv��ֱ�#��%�ߟ��v��5��ν����-�m��(�h�X=��;�1tSQ��<��yGx/�:.6��2���������g��X�Ȍ#V�u�uV��i�B�}��IN���F%�ۥ��'k�jr{C�7]���}� N��^Tc�s^<ZnID! ޶��$�3[��=1�۟��Hxa wGDs����o�y9�qr�#66�L^_������{��)�������Է5����ح�`��u)���=O���r.eW���,rkn�%K���&B����j���;�������DG��ƊRO���x��2��J�����\��:b�Ŷ� �<`v��_3ŷ�o�������*���¡�M��;�_�̀G��G�}��oW<���L[[.�H�Q�iS��q������n��a̜݊E'�0���p6J�A]
���ӈ��Uv�������U�s�I��o3������,^f��v�G�����Qcz ==X2�cH�r������$��	b��I�r���R�=���qEX�G<��+)� [{+r�a5����n)-$���!f�=���/�3�+:�[��1Xbv���S"���^��z�������h%�)Cf޻v�M)�Em�\7��Q�N��j������yժ;�ft���,Qv���t��������	�Ы�H6Z|���up��"���L���ţ����o��z��F*�n��5����̧6��{�V���[�bMA���Y�	e&�4��,E�7�1�� ˉ=j�DD�.��Vӱ��>��i)������� r^�G4J����k˥l���zj��|�'ڑ����k��|�?��
'��g���f�5�ߚ�w��x����yFCãQ��P�G���l�x��o���;�UHUe����-M$T��Vm�����D��.T			�u�SA��TJ1�܎�"�hoE��V/���|N���8�+̱�٬|JR�����9L2�C%���3�B��5E̯ɛ��a����x_��p|�>���t����ܨC�(�O��e�=B*�b^�Q����tSat���r�Ÿ'2?7�ς�E����b�`�k�!���2�@}�`��VE4�n�����O�Sb0E������v�_J���1��u�{���\m���A�jSY&�ʻ����u�����SGϭ�k2
�������(S�U��8~�M�ѹ|�#�э�,��9F�U��\d��Y��{����v�	�z3�ٲ }�M��Z�cϫ��~�����X��maݤ,���Kr��y�r˞�:-�#`�<:~�gY8,�\<8j����B�����7yo�����WHm�{��M��ئ�IK��{F��	���VܐA��o��������Ҫ����*G���0����Y��"�k7\	��q��p�1�4��7E�9uI��L���M����R�5�7k�����u	z�F~�ڷ ���ͳ��r˱*7��/���G8XT��7��������(�Bu��+M��e��0��o�yN?-{�Q��Qh՟�����fzs���,/�eU�J��*�ϭ~JAaԭ��1���;�	s��a>4�h���Y�O���d�}��*��I���� {{����J<���� E�u7���o�@rƇ+̛Sޟ,����Д5T�y�3|�j>�NF�8����I����\�b�R�ݷ�-�+�&���/om�sBC����a�m|������mO�t��'��l:��߮V�����O]�[/�PE)ջʎ����P!M�m09b(XooV�+)*
K�̔��T�T��;̀��m4B}�[�ڜޣ���g��]44뵋�x´?Ԑ"���(><��jNO�Q���I�����������kG!|,�+fB�g"��uM�k�ج��s��j6��ՎP,;��;��`�v!��`�P��~���l�n����p��X̊�a���'x�z���1���xo��\�Q�8�Z'�kK}߀D�˹��l�q�:i��#4?�Rf��O-����U��1\���1o��|kW��� ݵ?���d�OXρ��M�83E�D��^W���N��?rA=Gy��χ}z��Z����_k�x��	N635�{��HOE�nǞƯI�������������-�>]ȧ��.Ag�!��>\�FX�(󩕱�` ;�����?�?���[���>pF����O���k��HNRse)[:ĩ���S�=��	:�v��vF�?&�\0F�e���P�=Y"]��!(��D���˨SV3��ڿl~7�������*!b'�!�XߎWkM�b�説fEAńT�;�4����(��4r��]�7҅�����pݚ��K����p��SZdZ�D��o$9����9l����q�����YX���(O�3���;�i/�'!֪�nr)]��6��cw��K����]-���=���d�ef��21�~���TW2�>�:�
�5��m��c���}	5܃��>��+y{ㄥ�������v^wLͮ�wh��w�A��2sp�E�`w�&��^g�N�3�?U4}��L��=Q(�F2��kq!ŅOd�1�i�3j�^�n�·$x�1��i��`��՚� �F�ǰ����2z�-.���(A� ���/�X�pڟa�
�Z^Q��a�%jh�) �H���rcB8W�^�����o��]�v��$�ܑś�5��AJ�&���|0��IE��Cg 
<��<�(��I�q"�!�D���_�O������f!��r��Lr$h��}��>��X����+�]LX޶�_O�gj�v�r�9�sb��?��ku�0p.=y�<V�͹^���v&�	ٓ)�#�Y�S���{��ɝ>ko6乹ّ�B�0􃥴a�y蜄�U�T��f�\u=&J�e����r?\��e���8̧R&�݉�� �Z9��������m $�6�(�])��2^�o��o���F7��-��u�2�^Վ��KɆh�,� G@����>�֜H��j�йUm�8�c� �|���k�#=#�������m#Ҷmk|���W���)<����t>3��_��ĉS�����j4h���ϔ)��/SZZ���g�ӫ7�Oc�������w�RZiG1'r�Mmرy#�>[Ī�Kؽ�g��:�U�ճ3�D|�hߊ�߬���-|�:�Ĺ3'����v����_O�{�Ze��&�ٲi=OO{�˿$77��w�����}�^YC6dJ8DFj�<G�Y�z-=������{_
�<��3��ۇݻRVZ�*��)n��\F��Uede�PVd��B�����_�t�<��K�U��j����S!"�a�`��s]���t�4W	�G�d�.��Q6���O�k1��dċcžD�Ao�j�+R��ԩ߈����S�>��ߎJg��ś�v�Y�<��~��D#�=��[�b��ݴoۖ���;�>`�M4i׏���QP^��l���H��^%k���� E�&+^�}���F5j����l�_���zvN＜��=����׍�_rn �����9s&�ӥ_l�y�J�6�;P/;aäQ��*�"�i��k��=��Z����b��_�&j���6���_�w�H�?_,��^��1c�#�=6��x3���={����F�:�����$�gss�Qh�M>��4���{�mdg&���CUe%i�i��.�-VJ�����/��I�<��+6�T�(:�*oC���a�4<e��߹��ͦwSX�@mN�LxQ j�@(�w�r�>}��?�
��Gjz�$b�3�7�ό�p����b"59��d+�M� ES�-[Ƶ�b��s�̫�лv��W^���S���� ';K����ʫra�촧9{�
�l�Z�nj�#�Ƕ��9�U�%$�����>E7a�r�8.�Siw���F�Fu�>���"�4�3��#j�
���L��NN=D�F��ؾ�4�����_/�۟��g�^Ǝ�MfZ�lŻo�%Y��Y,\��)?Ğ}X��|�A?�N� D�}����Fj�J�Y���Z��9�����w�A�Q�F5��˥�N$��i�3�j���?j���6>	v��K�p����|Q���k���^CH�Feb� u��hU��Ū��0'i��o���~Y"�D��-	��'��痣|���k|���ؗ�M�1u�x���Y��\PH����VV�^͵�J>�j5C�=�>!?aY�}�m6t�<�PP���������z�s_������$��衮���e��q�k䮺��[���Ǹ���gn ���^��WRTt��¬�[N�x�y��wl�jR'���}�|��\��]�۰�ˣgη8��b ��J�	�֠yK����)�p}(B�.�8{t7aO%�^
�8�.�&�JNreU�T����6Cј�z�Y���Ɋ��ɟe��H�j�z\N��q
��h��p� �~K��Bx&��m#Pu��//=q?��BiZ�W����#F�*>�F���3h0��<:y<��ë3^�Å����&��L&#� ܭk*nܞ���>p�]�mL��y�Ժ(�nݺ�=aC��m~~�p�N��|]��K�ֻ��x�3�@��'�ãS&�h�<~�	�����W������R�^�zQ�	Q�t�7@�֭���E\+(f���MqTV8eZ0����IzZ"-Z��/�L������-,��kv��۶0|�`�.���Y\�\���ןM�7SZ^��%�s��C�;��{Z�kp��9�n;-Z7�����������Q�|�t�[6㻍�	�}2Z*��8k�$�"¤D�@' Y|�H]���ZU���R��0G�g�{��_��e���P拂|̪V�\�(��?����E�H鉶G��B|z�nFDk�^�h2I���-ӣCK>��6�F�'}TJ�
@x6���t�x�u�L��ښ��U��2�Æ*�E�SK@�K�&լ�8���M��Ͻ?s�G����t��3�|�M�z��l]���=���ÓG�������77 ��wO��+���5���ް�bic\"搃&5s�uk���[��_��\���Ǜ-�j���u�^�����*�Bf�EK��0�->*
����i\=��We�$B	&�� �P!�������JI�v�������=r�\8�Z���:=O@�Z�	��*#����%�ra�J���ʂ�4�3���_�&'T�l�b�f.�W�
�	h�����e5�;K�����ڳ+~0�Ͽ���'�����رY�n��'U7aѲ����1|0?��)�d��%5�ϝ;'{��F3�=�G�C���CbR<�׮�d�G�>$%R=a���^z����瓏>d�(s�	VW�������+����\�VJX��R0��2��GO����9y�\�u�0q��a���ٱc];wc߾2����\)�Ξ}{�N��n�
q�;v��YPP@��&ebE_�&MX�f�L�6��}{�.�FFjə����-^J��:�W�>�=��%e\8{�S�K�wq/T�,$��B贆(��ty�K���u��iv!���qȱ�5�Puu�}��6�J��V�EA��M��á�T��l"�/ljU�Oz��D���Z*�AN]* .55UXfO�%�ٰb	��Ge��y���T�==���"	I|��j��Kz^}�B�^��u<��*�>I$jū���̴x��uU�)q��hd߾��������yמ�5�u�۶}��
�{����]���<pc�����@���=�>��g�\�ӹ����Bn��L4��+�_=���;7]\;�v��z��7_�mǌ��5�Z\��!�2�*R7<@��;r��%ij5�p������h݄3�l�U�<:�k��-����>�ٳ�d�p�2��݄˧�� �Fy=E\��+���ڵ�	�5d�gIv���HKL������6���,�	|��"�>z�U��<�Qg���a��M\+���o�Ƣ/P���ˆ����5��ڶ9i�\�x���6QG[�D���&Q^^���[��K $z�5t�ҁ�8+Uv�����}�&mڴ��p�r�
^��d0����f����o��!E֭k��ŠSa�����s���h���n�B^~=|D�xy�>�qF��3�ͭAE��_�'!)��'O��#z��^�����&$�S�.�=Q���J�y!
SW��f�I�I�]v;NG%V��aĐ�����Y��d��<��[��8�m枻'R37���ߒ�.�-gZ=ހ�,�l�	� �1"�Ѻ���^�.�[�q8$,K�G��>�P�T��
�y5�*�>�K�8�' TD�¦7�դ�ǎO�$����I̮E�=�����T�
���a�{1nX�|4�xM�p�EJ��S7�{p���k֒�m��c�8̩��n�\��}n�U%r��B+NQG��Z�~��I���s�S���_��yiu�˛�:jh���O�>��¥s������]�.Resa���0f�S�����q� ����[����]/�������F�*G�u���@��42��g���6�[�`ZB�i��+춬+���_.����˽����%2�Tk-8\^�-��WVҼ�Mx�!��_�g��j�^E�JM˼L.��M�ӵcΝ;M ����i�N,���g砊��D����J��z���"E�����������A�f����^aCR���p5�U]�rѽC{t�
�-_D���گ��JMie�l��u+7m���Q��Q|x�KI3���H�(�ӡ ׋�0X��E-7>�,���n/N��ΌJ�}�Z�f��n -�UU�Q-"��E�X\\,���^Ѻ$��D�X���D-T�[m���Q'�#Z���T9�ęM2�$�  c����X�b�:�J��d����AFv6����$�J+�9�Ig���,��(\+����M�8�f'@6>!���2y�ɂ��F�;j\�2�]���9L�0�z5��}֤Zuh�<4��m�FeY	�f�O��s"�"���B�O�0��qM��T�Qc��	�3�	�d_�XP�"�Fڊ��5u���<��<��:���V3ee�v�]��ՊVF�҅-�G�F���X	�0��BmM���lA)�U�݅5p���iN�UOŵ˄�v
���_�nm��8u�<��v��~��oA���O�`w�P�
f��p�-��������G%�7"��9^�q���඘�F�ޫ����$^��d
չ��b��Q�S��~���!S��1d�>3����67 ��vG�����[_o/��p����6B�J�A�D���Bj��"&׈$��VS\RA �P\i�җA��'�Je !���P�A}�ť(�8��H��0(aRU�Y��]:@�Q�=�~��^-[ݾ�j5ks?_J�Q�d7��U�F"�H2�w^���I�In�l�6�q���� ?���}nE�$�l�~�O�v��آ9Mr3X�Ϋԭ����%���
|/,��'�˳�3���$fV#ͤ�FZ
�F�!�Q�h�_��l�P˫^�x�Y���<u�/ʼ�%Pc� *E� ��-LN�Z��(��FD�)Z�D,���o��V)	�q.2 ~q?���V Y@���q��e�*�!�D�)t�x��Dj�,�P��9�Ӡ�t�Ɩ��!�����T�L"(���3dff�(�p�[�&v6����D4��FNz"��BB�JFD�z)$';��J+�<S\�.�Ҋ*y�׭�������%T��`2���zQ�d|{\��d�˲� �UUUI}��Tjծ!e��"9YH�8��Qv��Me�CT�q;�r�E�\δoך!CȌ��� �������?�N���@�e�崓�� �5=��:�c��%�t)��	Tz#TZ�Z%�A	�/�N�Q&k�S&�E�:����G�N]�/)&�n��?Ŝ�Ftx�E[��V<X�o3��>��g.j!��0�A:���x�,%��(�x�!|A��Cx�
�E�1��<tט�;`�_`J�q��bn �_�Ѹ}���ۮ9o��L"AB;���@�~|.fa�)@-�O�� ��p��p��z�	�V�L�b5Q^i��s�Ҏ�d�Z�l�Ue(�6�e$Qr� �;�$'+��k��Ġ5k�1x�����ڂC�Gc��z�&H��Ǳ�[�v�
�}�.�P�ƍ�
��kiX�)�l9~���M�(��Y���KO�����i�)ڷlIvz:��Q��9.��>��C�P�^=����&1�w/��:-6[%���H骑J`Մ�5�����g$�J��5	�dE$/ ������K���t�e��&�.R�⍤R�4�Hˋ�R���'��Kؗ
@�,n��7 �l�"�uy���^7o�~���1>�'HRb^���ߏY�P^r��G���2�IN��B �f߁�|��v��D��J�~bRnG���Czqϝ�	z*Q+vU��A]�>�'D&蒤%l �c�{�P^VƂ��Q#'�ʲb~a<h/5�%Q�z&f��Z+;��_�Y��L���I�T�p��ت\���ә��B���%�FCYy�|�-Vn�Ո�J�^�9Lv��(eg�F��Q)�*��
5��s�8��%ݡ�'lH�+�8�,f-��^xm����F0��^\<{��]��j�Z>��3�������D�JH-�XK$(�o���_�_�/���D��S	�d5Z4�#b�"���)a颇V�/����t�ӛ4T,!/��c��[�����x�����/��d[�c�]ѡ�	{<(��`�ۍ�����eGo6��5Rg]�5`Pkqڝ����Tku��&��d��\�3C�OW���L=x6�.��S(8w �N�Ly�����gN��ǝ�HʬN�7�:1G�,'+=A2�Z�6*��#/7�vZs��X��wnێNcD1�(�Hϫ+��۵jJ����}4�M��r�z�!�=/��_s�r>k
����^�O�g�}�Z��Ԇ���ONZ*A�[���m��Ir� �̴TIhzIwao*��D] �H��~em�I[����R����Z��T�KM����o�n~�z�\<dee���ș3g$����㓀D{��+�����"�E,*�]����&#u7f��-z��7L�=���Cpb/�L��K��Z*+�����h�	T��Z��E�m".����sԪ����QqU؅�8��K$�B����JL	�����~���4�ٳk7߮�@b����Fj�����IO1�񔓚����e�����%M���zY�Z�JX-�f�����rE��7=3=U�siI	qq�v�K�\��rqͪDH�F4��k�m�8���p\5�6&`�����̚0AGj�����O<>�	w���?B��2{�<�,����ǓY����V!5Aa�����񸜄�I�Ө���h�%y�`�BK��8g���J'3gE�V�#�b�B�.����>2��ҿ�Lw��oD��g`���>�}� �    IDATr�j|yD�F���z�Ho�Մ���M؍ޠ��fG�7���Ъ��<>	�n������ ެ%⯤n�\�?E�e\�^N�.]���F��fpI5�q�^�_��dV���ųD�����S!�f=���M� k��d�n;�0	!7珲a�֮[)�V�6k�Y��[,���1�瑔]���M͛R=��WK��y�{�h�����g/�����ڵ����u��=r,M���[��hb�'�L-�%���"j2��٫$�fgdbQ��GQiIT�D�}F�� ���).*���v;e�)D\D��VQ)�.�$& ]ԅE�B�/� /~' ���V�I�_��b�n�^�7^����łBԔ�zj��~���h���8tz����жE]�y�)��A>[4�������V�c*�EF�*���+��bR����g�.^w%h�XQkrq�,:��
qi<��dW�c��[Y��*�j5��R�zMT#ު���@^Ge��K/D9��^d=T�t
���t�*W�c�A������)�F躋L� ���ע�x� �$�A��&$$Ȓ�x���k�p��5̩��3|�����@�ϡ2�&��˚�����r��ZlŅ�~��tm��G�H��9s�%�z.�v�g�$!�!uD.���Z.�P�х�h��ylH%;��.�(�R�Z����JMX��?�F-�|�
.��*e⨁㟺s�Վ����R�x���{���,�z�jB�H�	U-o�ڈZ������
��!1���V����W�dn4X$8	G.u�K�t+���W�6L�0�>�o�~�&\*�g���h۸���[{�h�z�"f��������D�;��*5���+gN�j�S͢��8��ﻗ�+�a0�Re̠���+E�h2HͭE��O��]��l��wf�����^}q�},�fFK"ղj�����3r������Sv�Vo�YQ�I��g��V���ĚG(�ZV6��J�ŋ��iXR��& BHז����������
�ɿ|EF��?��ɓr{��ԌL�Zw8llRRҸv횘��q<n����)�-�".�1u4q����ވJ�q�]|��k\^�J�����ۇ��w��go����кY:>�y�R�8i�"i��Ë�d���ZB�L��Y�D�.�� �Ȓ��|�>�����3e<��L0&s����̮Cy������{ �ʴ��wN��izr$gPDD��L��9G0gE1�a]]Úִ��3���4�����9������z�z���}�y�ٕ��f:�s�p�����6�"�����s��S�DQ����(M����&R�T:�r��� �K��dȐ!J�P[�@sS�P����Қ�Xm�%G�F"�QZT�H�҂w9��TW)ЌG�8]Vex�$��w'�}-#��H�Y�;kQ]#!:��E��3)y������F�!���_�0�P'ɜ�SA<��_\�n��s�"[�٤�e�u��͙d�$���+��>@�a���A�&cC�+_z1ͱ����=���l��O9���Λ���`I���[��{�ܥw������,N�ٸ�%e�i�����XrX2��AL�}jV4�O��m�Pld��#�¦뤻;��h�}˵���Ӭ^��^x��o���N(؅I3�W5�h+]�X<nb�#j�Mgs�*ٴ����M����<�cAj��-ă�$�m`�)H*C�1���]�m��-{M�����瞍�H7R�wFh��{�p��:TkS���_T��bG�9GL��_�'	]�N,%�	�\q��,�M��`˖-��mfs��L	�C߾}ɤ�=V��hO��6I]�]Z��B��� ���:�sL��VT* ������$�H�2G�*pp����c����簉L�Hc^�0n������L����x��'P�KP��S�]z��Mx�b� �e�}�V������%�[�����rani9�X,����D���<��r��8|������y�y7�Q�{3�W!En������Z����H�q�Nd��[��ѴYI(�G/Ns�XJI5�\��HDU蒈&�T"�X�}kz�q9qجx�N�bn���PX��U�:��.aܑ��qU������"���j=��d�D����k�|D�qJ~�VM����=�a��&	k6u�2��%U\lNȥ��awc�2J� ^����ɒy��Wִ���m���n$��'�kX�]~<v'2�?s��K-���w����+���=p�mK���1t^$oGOd�'L܆�"�͌��c�p���������A<�"����j&�%������:��f�?�T����(��o�x�~f;�T"�����O⛯V��LB�#�C@.������p��#�1ge����dJ
<��g�m��֍�,lՒ�<t,�6���X��x�_j�q�ln �T�˞��vPZRA$�!�ż��)��i�0�	z,�{ٲ�g�>�*�SJȂ��բSSVFaA@�A���&S�5��E��d�) m�F�����Ѕ �R�2&6�CI������V�+�jjj��󨖾$�E�q��}>���s��i�0���9/՜��:����2o�[��s_|�^��͆��8hh5����wY�i�*�ib�*�l%��+�e#���uF���e]66r=V�"�%��"RF�!�i?{	{[3��槜yލ,��>���(x������y��ٲ�G���^��
�M4����s�UPf�^�]i�e3v����y�L��R�����l��*Xω����bS��σ�aWպ�Ӊi��.�
�;�W��y2����y���V5m��i��� �Վ�I���p����dg�.;n��G�f����L'p	��Wy����dr�~M����2�E���S^���2=�]W���%�f�I�N���'a��#����3���k��������?�����1qNG(����`&S��*Uz"\�3��L:�N�~C9��E$�EtD c��}~l�"ipn5O,
�;f��By�ν�B�}��L3��y�g�1�p�M�����`�TZ�����IkG�/_͡��9G���'����r��ש�^��U�Z�EU�ƻٶu�~�3�<�$�X����}��uQtw!�x�Pk3�x���J|5��#D��1��JcIg1L[:Ju �$ik�%��a�Qmf��)9T>�ݰP��(�Jz��]�y)�T��0�{
�*6��c�"1�RAoPf�� %�2=���ck���/�n�@��gr\=�t�$+i�M��&E&����˓/`s�1,643ũ�f0"̝>��b�V�c"]'Z֋UW��\͈AN \ Ī��\F�9+��������]���:�$L�|���gs��7Sի����N�;���[n��ֱc�V�>'�D�8����u5����9z:��M��)�/	;�(W�YdL��>_�ekK�v�)��\����QVZ������ҹ'���a#���+�ǂ�e��s�xz�*Dk0�fH�Aê'�%�hW�|�\�d�y��8ٶ ��l~1�`٬�;�*�=�2qy|��$�idt��cGǐU8���0Hf�dE�`8��v�(���p9�$'�6�:q���W6ŝ�pڱ3n������,i�Oq���{�{�M/}Q:��ȡC^S��'C�Mt��f�BJ|a�z�h"KSc�{�~���	���G��
kފn�OY�sS��hY2>��n��VΘ3����p�M�;f6w�xu��Ȋ�H>�����U-~B�9�E�7��.:����g���[o���B�[�F�hee�b=���G������X�j5�?�[�:���2���h6

K1�~�Z��]�Y,�ם�`O�Gpf;�]�!�ZO:�L�&;3lJ&%�����V-ۼ�cg�4y4%c��P@V�z��zf��1���J' ݣM�g3m��*�G�b|��w������=��9�d�ݣ0��%nB&�j�--٬��!�b��5=�5�N&⌓f3���1�p�B�Y͇�I���.�M"х՞°tSp�U�:�E�3�T���x�J8l��V��ɋ��lh�����'�Y�����bsi\r����Ow��U^��͛	E:�H;]��r�8=NE�hk����G���"�ݩ6�mm��	��ٞ�l���B���+N@Ks�-[w�����W�|ڦa�B�*�W��9|E����7�RL{����t�D�o$1��O����腸%d,&v	pF���js�
x�n�pډw�Ԩ�mbW �#P@kG��"2�8EŴ7֫9zqe��H�g&��c��g3XB��(�|�/@&*����U:|�8n��[�����+��3�_���3o���O��w���7��'�f�q�����.����ڢ$�A����]���x�5��]1��z�����w(��!d>�xq�	'��s1�M͐�2n_��>��̛=�%��+�s�H�j�������������;)--e�9
��͐����,W�q	�uI$�
���'��~�׮a�Mw�=d%��G�ۣ�jw!��ЈYR��)�,�Lb�X7�X�+K�H�C�D�פ���ىvK"V�j�
y��=t�b���������ֆ��U,�}�d�.�K�-@�N��ɊP.(葩��$MZ�{��U;�^��9PD�x��+��4��2�H��q�Ӫ�/��3~*���T����2g�xfN�ءn��]�� ����|���J�]Q'Mq�h�3ح.�W�ki��뚝h�Z������ha��*J��*���,$g+㹗>cμk���{�i&����E<��C�p�tB�m4��������]v\'��6��-4r��S�3�kt�	��,V�&�❭ab���ށ�aU�?Q�Bav��MSs;�pC�:(��ֽH ��g�@/�\t�1{{Íi��b�sX�	Hv��/��p��kd�q�KE���qE$�M�8f�0�nb��uz�f��"� (n|�	n�]�n���Zte�[TX�a�H%���gu��[t���hohR��f`�cH9��)�>p��w�������B�}��|^��λW��i����=��1���6�/�A�r�DԼO7�8ܥt��F��������{��ޣ�|�46�e��*�~�av5%z,ał3���̂xO=�$�>�=����aӦ��Ң�a:���h���ıǝ��)9`�HfL���bg�����d[t�_�Y*�c���[��[����,Zr/���pU�J��ߋ5��������y�R]a┹|<M�+�4�#��5�OG�$#�ܶM�˧<ǥB����[U�Z�R��۫R�lv'n�K��1ɢ^\\��[g�ڧCW�/���U
����.�[S�ȆF�o����W�˿�eS �&�.�!�wi�+��dJ�#�L�9��Sx��7qz}d̸2��z�������"�B6�J>c#����?���Ƭ���q�LJJȫt��P��ș膃x,CSC7��W��J/��B��B�V���+�s�����V��D�9�t�T:��1zxo~��{>[�����{H���PG>gꔉ���M0b��z*��P�k �T��֮a��݄;D������95ϖ����}�ۻJ͜���{w-�~بd��U���{����J,*�˼��b�	����T�
?�[���b�CKc>kq��bjYe#R=ql3�)2��l=�?qS�+:�X�Ds;�����EL5v]6m2�ɛ�\v�^�K�ꛔ���립��b�
�ӥTF���>��n\t��s���r�W����ASS��^]�쫯��9�`�D-"SˠeӐ��fԂ�E����j�v5Ö�9.���,}��;w��r�9)�Տ�}ga%	���E8�I�,�+��_U���^��N*��Q.s"���Å��e���L�8�O:N��/��2����+/娣���8���SJ;�����BKs'^r�X�}O�ۃ$4VL�-��ҧ�����f�����<;� �!-^"�-W������ןb�N�UW�i�ŰŤ��3���0@�߫Hh;k�0���SY^��|RA�u�
] [lL�('�/�$af�^f��s{��	�0K�����.ϗ�ľֻ<^���sy��aW2�}3�������2�8��pyt�'����з��q3G`׷�4�e���io�Vnf��6����'��3j���6Eȓ����8����x�HmXl1,Sɴ91k)��e���o"M�)�{�5f�8��ʹ�yh�N�9{�ٗH$���=�i��8b"���n�h�[Ϗ�70�y�"&o���nbf�������W����\]�ۻC��<V���9�Ѓp�zR�:ں���rY+���6[6{�P,BU��\���G�F�VL�[B,o!!�p݊5oǁ���F�������������d�Ø�S�]�B�r{ˋJ#��j�H�)�(Ô�T	��d��\�U�a7Hf������X(��_��[�������%O&k�Y�zlx�a�:l�����+�͗�����\����o~{�
����_���]SE��U�T��R]���ćJ�w&�����M�Ĳ.���x�v^}�\�)'��֭��?d O����c=�3���t�&g��rݍ��d���c&{�x:�4���LVT�[p.No���U�5}�����3~�裴��)�g�^�|��:�p.��Z>��[.��~~���IzW�PS#��M��"�b�aϢ�R$Z��F���"]t��l��3�>�����ۿ�J-r�1s�}�r�8%�E
tٲ���'������P�@���k�Ke-�2J^��*��}a-چfQոH��R�Ku�#}����o���U[^� ����tΰY�J���MЭ�j�������LFGك��0';�CG�Q8���1�d��2�yɛ����e��(Ua���aq�y�)�x��r�p��Q#	�W#���J:��]0�'����J8���k+�Y�p��<�o��8����5�DS�a������x�HJ�<�#!v���G��ݭ|�v=I�Jw2E�j�[���n�鰪�8��IZ[Ȧ#:()qs�ac���6L�sG=1�9�5%>�'PRޛS/����/�R6����D�4�8��4���hX�{8
H��y�@�?y�6�����ID"d���T�ײ��� �y��.!۹�<%D�q��Ie��F�d2N��O2��a�b��Y3�S�n\��2d��3��ѓ�>��]�^�o���?������v�
��x剏?�����/>�#G$�Y�I�2�P%Le����b�wV'�1��=��V~�i��s�Տ2�ٜs�����g0?�w6��IY�� �g3����[�x��֯7��������N��0��޵c'����;w��1a��̜9�ѣ�r��CU�y�X��7>�P������q��~'��{/�R6���5�~�鋯gSP-
0��
�K�B`���E0G�g1�Qb��9���R�8�:� Z궰���T�c�MF��/�6�4����Ś/>#SVR�*�M۶#�n%#33j�/_"?�0�`���Q�T��*my� ��H%�k�.��T�آi�����H�/�+_R�����(.)Ssb���*�l���;�"�H���<`� �N=��?��^����o�8�dS�D��y5+7Xm=<	�Ѱ���b�K�YK��tNm8Z;�q�
05'�\�L��g_x��ʦM����^y Kn^̖-_ѫƥ�w֬�@��:Z��̜>�>5�j����1cƑēYV��P���/�;�!n��x���ۉD�t��I�M�6N���U�5~���}˘4�`e���a��Zvl�S>�"k��}�Vp��L��G�b�:�9�Yf�FΎ#�a��H�����I�v,v�R/��,�B:P"�4cqR�Ң'�B2�$����ƚ5����(�(���/��\�h1O?�4���^y�a�r�Y���Op�Wp��ת���0,y����ژ3y�s�~广��n����������G����/��fܝ7����p��'�V�N<)���LP-��beKǱ���^��a{���H�    IDAT~�Ҋ�DÍ�w�}��v��g�$�(#��csX��:8{�$���~n}�$�!f̝�7��H8砑#��˯�������æLf��8���8�ؓ�6q �U^�rｻ���ǳ�~��ֶY\��a�\��|��w�fly�TW�|w���jR.?�dÑ'���o�m�(*U�ǱCk(rk|���x��L��r;���Q������Iy���8U����BBTh�D73=�2#W5�M=Fi���|/ /����L�K����+S�����	n�LM^W�]�\~�O�&����$PPDCC�bۋ�O��:BݔT�������[t�����qd3<��L<��'��e'�RNs"3S2���vى�ġΦ�ǥM-:q��V�������)=�f�U��0]쪋sϽ�0邏(,�{������ﾓ�"+����H���e˿e�����k5b��*�j��|�"����kXlNr�M�
�����Q�ڛ�[WO.�����ʦĤ�����b���¢gH�"4�ե�6��+��*\P65}z3j�Q�~��s%���y+�|NٮZr�\["J6֍f�������݅�n'�H�7t��Vi��rd�Q��.�=��/��f�w���F����Xr�-̘~4�~�=\t1�w�vl��k�U��V��[�,�ȣg�N��r�֮��'�\��
�G6f?������������+�/��]�]�G����Ͽ���;o8���$��{	v����
J�+��mW�.��ێ�e#�uS����-q����0r7ߴ�];��sg;[j��rSyg1`1�̟>��3Ρ��'j�i�P\SMqE5�\���{�lnV�-��:��o��G�v�9���-�&S����Rı��:�!�H��-{�%>����b%k�8�&�f�J�
K�͉!�.b���\N��"4Rk��	��F�İ���4Mu-��䲔(�a�Knx$��&R5���z�i�&��xU��Ţ~�����%�'u���j"�k�m�Y�
���k�׾t7ѳ[�����s\jk�D,Pt���hR�z�R�83����.�q�z�o\ɈAVƍ���7*	�r��D��Pճʓ���d�d�ҳAz-zR%��2��e'�y����-��o}IE�Xj���;�\i����g���l��C,��Jl����૵?PU���fSYYL��դ5��������+,�v��[@(�$��MM-�z	�Q���tѷO/�k�q�,4�瑩v'6N;�4e�#�������;ҦHm�7��ǟ��W��/71]�f4��`�[����p�\��|ޤ���\^��r'e]dw*�E��R	<6��fL2d�I�.��~�]|�����'w�u��w7{�En�m)���_ˑG���e�����Q�O>��1����q�c�)�z-���GOy�ޛ.��_|����W`?��?\����A�u�c�w7�{�+8л�"#BkS���~�'৺��"a'�q�D�{�h�<���M;s����'W��<�=�0�����K���b	��XO3�A��x鉇hnꦬ���m[))�n!�]]�K3�ѩb#�*1j��_���w�!�2v{���
���vZ[�j�,.��.����?��������1����L����=8E�TPD.PB�~;�F��1�(��P�)�����my��I������!�L� ��sO')-.T��ή�d�l.�4�� T@���Z����[e.� J^ ���ޣ?W�ߴ����}����9����;!���7B�r8�$	,��*|y�d�g4'�X���ǥ{bf8|���1��.?��"x��p�IŚՌ<��(��l��4���n�ў+/�ӵ�� J�.0��L�-�Wc��]�%%NNZp:�B��ws���{���%�6����R�-�>c������1w�Te��sG-4��>���l����Mr����B�k��f�,6�ѓ�#�5����c�ٹ���݊	^�+C��cG)�6}ks3����Jx���!�8b�|vv���X��Ӟ��HS��d"���|��������\���\^"��b���CX�:yR�%�DB����R�G]S=���C<��|e���(��d"�dm�!(�~Gg���a*�	T�U>��r_0��������
���c���������yխ�[�y���?���	�/��	!<�B]RIZ���$�%�X����P-w����6v6X��Η�5w>�z3v�h�n�Ec0Ɠ���*R%��)c9ﴅ��қd�I>Pٗ���g� ��-Ic}$�������pʂ����䠃��^'���j��qQTRLBR�t�J�ڹs�bv��7��۷r�K�j��|�7B����$��[���QVYC��!�RR衽n��Fn%�z�3h� ����d��Z^�,���Q9�^�S�R-�ʆ�bq�h��e�)U�*z����d~�d�T%.D:�PO���LJ�j=���&@*�}v����6�>���L�l>�:�� B�'�]��1�8��Sit���O1{�$��y���7x���0���h%�c5ܤR=����B��G�ұ�
]6'*3F���|]���QΉ�]B$fㅗV��ۘ>�X

�L�6���Ɛl�E펯������_SUُ��6��g�0��~�=Xi�;�Q~8/����FyU)�1�.���V2�,V-���	v�����X]�ں�*<'�);ڢ�b�.t�C����G�0L���{��nPuq����S6�t�8)�l�&B��9
�\KG0��y畿��ǉ��TW*�m���t���>444�u;յ�G#t��0f�p����	SP]�Y看�4�j�E��t�ˏ��bu�ŵMX�ٸ�@�+�8���))������ǖ�`���wÅW��Y|����������[ZZ�w=�����~>���e�P#V��[P��-�H��)�����U�T.��F'��N_�(g�s���n��{��WT��O�����b(s��GN��J.��*|?�L\%��W�+*&�L��Ј�ˣg��,9&r0W_q9��ɼy���L�R⿥HX��W6��-�M=Nj��0o��wy�eַg�V��$��왬
:�{���^��Hs��6�!(��Ku�D7fw;nR�ۛT���o�Jw,�.9�yS�$\��3�}�TȺ�U�2��*����O��<O���M@P���U <�������^i��i�o����<G'$wݰ�*�Ff�}{����Cu$�,f�I�I�׃�K�����y�q�LL��[�	�EG����T�,b����FE�겫��p_|����o�<��� �H�[%>Cé���*����`N=�l�æ/�SQ��c�����3�q|�u#?���!�˙p�(��鴎�[͇��_XLEu�%��I�}�{��k+��+NGg7�x���V����B:"��� �����,i�n�GT���۷+�E� ����9��ٺF�X��9?Q�`��\�l<H�����������҆�Em�"f���88�ǭ���~�\#	Z�v�J���w9��sPџ�n�	�mQ~�CHu6qSy�7u�)R]q����%4��Rv�5���%�Kz���#����S�r�5.��]a�����+���'}��":�?���?���)�s,'�r�uo�j����b5�3�\�9����
���4uxc�F�y�s,�B�x���६��k��Q�KJ�I<��i�8���5u
]|���`�T�����Š���-��҂�f�:���c)�bN]x���nim���\���<N�`JB���I+:I�j��w^�����n��FC�q��]P�VV�ڡF.���hlU����5d�g���&�Z���>�҂r٭K��-(�~6���W^����e�}�7߭���+���3<��?+p��O�}�/W_}5p k����_~YU�R]���_������[���Ӆ�>g�n���z�e��*O62���k0` �?�<+W����K��G�9�������jN=�Z;�t��r��������yGMLUa��eA
\ar)�l�H��8�^��4V�X�D���r蓖���������FV�r�g��������V��;{�nc�L�K�a���减�bp//f��5���Q��Fv������8p --Mjv���a�6��n�tEZU�ؠ���V�cS=�w��"�m{]� ����K$^.솝d��j1(�9�Y��
��M��~�i�m]�>`�r��|̙���,��!>[���!.���6<�<�7���W9u��8�p���	�A��3)*{U��J�u��g�;�$�	�A����k>�ȣ���?dgK︓%w-������{�K>@FΥ�`"�H��.a-i���+�����O_�����,�;�o�\s�����������_���=�;v������y�����Y�{��|�C���DK�!W��$I�$6�����?>���3��ꥏ��W���Ȧ3=1�+]���C�U�������~�/+�Yp�1|��J�����`ӦM��v3ä����+�0f�f͒p��9�8eZr�E�y�/L�2��ӧ��)��_��Ĭ���������p�C|ל´{U�ޱw��k/��"[TB,�F7�8�)���*G�קZyck���;�;�P��q�Ջ��۵����q��W�'��u'��駞�7_'
f͚Esk#�>���o]�`�F�R�.�"���|�~�a�/_�F�&Mbǎ����J�6{�l�W/U�^ȫ���'�|�_|��ŋզA���{����|���7nܨ�lӦMcŊ��~�T��ӧb�h�8�eJ��t�C-L?�	#ʙ6���f,f�bcK�Z6�W�T��S�6���]�\���˒
]Z�F6�#yT� k�Hw#%%���	ʑ����6���/��.$g��ç�S��o?e�o5r<{�r��q�&���<��m���o ]�,���drV��~k(-+Q���;j�����o%�2U����e�\RR��v��স�ɸ��^S]��'	:��iv�٭��m�A�TV��q��S(�=�w?���>Cs�F��'���gS���x�N8�$�Uܬ�K#�;y-�����Q�8��n�Sy������x������1}�L$�������NQ��]3���*�;,�C�GA�k�Wyg��\|�ʹ�DN�aKv�`ִ�����k�����_��������g�������3fM;��Fz�WN=i�H���Z�,�\3��"�8[1�?�Ľ���|,g_v;�x;y��n�0��Z�?{�u��>�1�&�������7��x�MwRQV��S�5{&C:��;w���ҫ��-?�����P\^�Yg�Na��sθXU�W]��s�;Km�x$�Z�m��j_��+^z�5�y�|�����p��l64(c��>��{��f���Q����E��W���_�s�s	6�r�������p�
$ϲw�>���w,��|�z������s�Yg�ᗟ8��S�Ỵ�>�$^�&�0a����1���
�6mQ <y�dV�Z��p�����W�~]�y����_��E��
]�]y�;j3|�p&N�Ȳe�X�n���8X=���������[4w�h�L�-�����%�����[�̝ڏ�s'VZUvx&i!v��jv�6C�8�	wA}i9��U����cY��c�J{]����pJԷ�9j�X�~�EY��&�ȗ-��5k�:u{:�l޹�qc�0�%;�m��ݴw�q�).�������F~��W��6(|2	9Å���*�dz
�Ǧ��<'>����J�
*�6����?��6>t���~޼���69�f�@���i	����'Y�f3Y���i�Ț�Zv����0�8��Cku�����gL���J9P(&��V	ہ>}�s�-��|����Ex
��+��֥�����l��Vq�3I"�:Ł"ZZ�C�����*�o������Ţ }�i������o����������[�X�Ֆ�G:��t-����g���p�N���Hg������fmo����X)G�|Kz����-�0h��XW'.��ۀ�>��3O_���_��9�s(/�`���).."��t��xCϡ���74q�57N������ES\r�e�5�[���3N��ϿRȡ�J"gǎ_)).��-�	����;������#GRw��qe,cO����/� &�:u�cQsf���#�w�'"d�Z�1� "-uq����n���+ǵ��2:��7�l:�f�[6������뵟q�q�ID#���GR�x�g=vm�-�1T��}�j5�D�>���ŤC�SSS������	GR�z�lk��C��w�ǫ�E��\TUUҧ��Q#������?#��aj�,}މs�S�{+�g��ZB9|E�X/�p�a3�)U3�T����4b������)1��n�j3).�Qpc��X%+1v
 U,l\��#Owg�T\��4��Ng�SL�mdt�j��<�l�+��%���_e����Y����ʸq��4u~��3��Ӧ��PK�����Ҋ~6�Q��6lT�q�.��ɓL�0�����i5c�z-�Wѻw5U�#���u?Q_WK����}��ۧ��ɞ�z�n�A�j4��#O^Ha��Dr�|����^IG�F:k�s���Ț��3�B�nFП����3���?�����e�֭��w���)/��no=n��g�}��?^��g�A�a��`��3UǦOi�z�ۡ��T��@�r�;e���~�R,6��>[Ōy'��T�t��gO{����?�w���?����迃[�ۗ��uۧ��	L��s@u�fL3���U�2������y{���v^z��q*W��9G!��IN�]i~�nl�㏛��/=��O����?<���x񅿩
WHS'�x��!�9LݞM:��n�wA1'�~����c撊DXt�y��W��{��E��5��������ѣ��ǟQ����~���Y%1ri�w��g��T���{N3�p��-Xu��C��#�&Դ�"=�y���C���&��λij����Ey��g�f4�����%�b��;�����߱��/��@IM�I>��SVS���pݍKI���<0�矸���7�y�n{�E"I~��)��Χn�n���w��h
�6�;m>�|����|�BQ�+;>r Ko��֭e٪l�U�ގ$eUC�47Ii�ƺ�5i������
�Mz��}uY�ذ��XԤ����*q838]�Wf�ndT�.�=3m#�i#�PG�iS'��w����qz��d��7�og��ٌ?�h!��ˏ=��eo���w0z�!��4{��2i�!*�v��j�PVZMsk����%؝V���%mi?�,v

��,��s�1%�>N�>Uҟ���.��-lۼ���e���3p@5�z�����o~������*�C�L�1��α��Vn��m��Vb2���7���O?���qŸ�Pa0�r�c+)*R�����j�ذ�,V;�@۶�d���嶥���F�?�D%ż��9v��nK�Z�{o�c�r��cf��?��k�p�u׳�{�U�qڅ�ўw)�_G�Kdk��u�y~K��S���{@��n|��U���u��ic�a�(���&<;b��J%@��Ƥ��4��@�He��������ʁt�S*��)S�b_Y^��3���og�c)+*��ۖ2�_j�+T�ʴ#�c�{2��b���_�l�/�1s�	x��T����I.�``E9}�����8�J��?�@Me�?��#�?>��W}čw?¶n+I�A"�D���
g1�*�iOCZ�Htao�N.��x�x�V�x���;R�ܧs֙�PW��������0C^Y]�̣�p�G�f��<��g�Z�|�����ZD�����=�/�[���sgM��Oa�'�����Nd1�&�2�C���Oxw�g�5|n�|�~�名���?��9����;��8���������ޡ#�Ewب�*�֛.e�>�t�m|���d�%�r4�CFr�Cm̛9�>�1�͖@3��$�h�t<Ϯ�46�Aޤ��Iy�O��%:�j���<C�F�
6�l���R���Sߺ�^�J�Y2$M��7�W|Ű!�<�(�U��f������V��H�    IDATq�vFҒ����i��RZ\Dc���ر����0]!���J߯[�����P�	"˳{l���0�7���w���آ�{ZΎ�� ��8XIr2�~������|�'�7wQV\BU�ތ8t<%��Ԓ櫟ڸ��W	g
�Xm�&�u�P�i=�F�'�NqШ��t�w(�^�*�\'�fT�W��`1t��>��y�5_~�E�+���/��%��I���JE��'�zR���f&˙g����x��g��s���;\۽4�Eȓ�����x��k/<�����?k5����@>��^|��+�޸yڥ��e��v\�ZU5f3)�_�,ֆ�g2,6�����ش[c��%��QЋp:IF�qټ�0�#�h�3{
o��'̝���駝����g������W�Oaa1����5��6����w����<J[0ȕW,��*��U=Ju��Dg�Cc}�5��ٗ�p�g���O���o��CW�X{���Z�$�U5�KK�Ȝ��$�لѲ[�΋��V�+�N瞝�r�>�G�K��]t���FU�N��K/?�Q#G`�噿�t2��j������#[~���W���>���G*gr�e�p`�rZX��j6l�AR��v���<�ަW�\q�ͤ�(����٧���~�W���������R��o���+��������H��:���cYp�LU]KW���9��*��(!�FKt�p�$F��2v����Z��%M.�#����ޅݞW)h>��T:��p+��k�,#>�:�E�$�Q,F�t.�'�"+.u�̼�W__Iqas������+�S�����y���6�pv���q��ۻMM�t�X��[?���]aVQ_�h���A/�%^Vݗ²"�>�Ɉ灤��y���
���M��G���j�_9��>�덕�2y|.N���N�UZC}g�����߶��)�x��"��3��OX�բ1���6���Ib�#]�}Cy���iV�]ݬ[��G��o���_u5N���︇/ZL2�͘�8e���}�y�u�dYx�O$����˯�7l���{�q�Dm��a�Ut賦.�㍗���^����v������)��=q�u_|��Cn��T��i&�4���L�Ѭ�;�Q�fS�c���,�z!�-.�}��wV�&d��x��Ri�qK6OMQ!ӧL��
V�X��1ƌŽw��u�\��QÔc��7�� �H\i�;;4h w�qE�9o�5�T�0k�z��p��W�p�x"IJ���p��N������7�ֲ�<��k����h��hd3a�Ar���2~iɛ�:I�7�m�U����;��H�鮯UN[��7��;7�8r���^l6��_y��^��2�b�w�����ڏ3�ċ�=�ѳ���G��(����??� �?�0w-]�S�oۡ|�K��X���3�(���znY���ٳ��t�%�T�ч�����G�)x������Wl�.�����f9j�d�L;��^���f��'_�%���9��.�n���̟=�c���c7�������#:1�4�ėI�HgbX�y���N��KKYHs9t��ck�1�bB#ĭ,�h���dƅ�ۛ�^Y����^R����v�]9wWwu��Y2�(��8��� "aT�1b�4F�9 
�������]9�����}��u�]��B��jŖ�]{�>��"}揞p4���hJ�h��^�ࡣ�+.6m�ACM�Ǎ�)o�B�/�\φ{p��2��dV�lf�.��NuU%յ5ҽ�`kM��-�(>�Z �PY!�_�4܏U����&䥼�-�b���;��*B�rjz3a��q�֚����t�������o��Uo�����GM��1å���K��BO�d"Eɤ��e�;�'RTWײ��Y��C.8�"a1�>ƌS�$pӳ�͈�����{��BU�rBr˭7��u^zo%���f�Zν�Z&����i�>�o�է���^���m�/���	�?�S!�e�}ꩯ>߸n�5WNႣ]�{0�|�;c�
)��d��'��$N��A4����Ư;��x��؃�Ɋ�-�)^1�q�x�I>_����GQ,����*;�����}Xx��Ȥ�473n�x:Z�d~����Q,&�gYT���`�g�P�2nX_<N���0�P-�5�r؉�lش��m]�2�D�N��A�8��[K�^�B B-��)�PJ*�\�d�n�F���% �t��][!����W�ȣr�gP����*�2v�y?W^})��>������{��XZFfV�}����\y��9�w�_�n�0+K/��0��Y��Gtt�Idu,v;o��&����\~�E<��S�4;�b�)�&0b� ���
E�~��bI�@u̱���xnų��e�᨜�8-
�y:��t27��V���bt���݌/����?�?C�|<r�=�+��=��b�C��h�sٔ|TE������a�R�P��_KB�^*�u�YS�{-�drv�F��_X=��_�1q�X��{��������k(h����^+�O��R�T������'Ғ�b���;��I�^UT�%AO�;v����X$��f��,$G�G��$1r�&Qx���WGy�M�^�|���|��O��j+B�4��c&��9���������
�EM���䨰�X0�rP$2�v�/<_�����N�R91zO�3�S�d���Iv��#�g~��]�8��.��7߆�n��܎��b�қ���QR��c��f�\y�9��^���7Ҫ;1��;��N���=7\9�d���ïC�8����n�n��?�oܳq�U������<�>�`-n��;63��)��<.��[C�Jd�N�����p�#8+���Y��=法/��W�-��ϵs�c��;�I��`ܸ#�j��`����-�d�J*���/�ɱ�����K[s#�q.<�d��-a�%�L��x,�a*�}�n6l����M����类��������>]��jeD&9sN'ִWfTz�jVJ���Fj|�`f�)Se�����tFH�ø}v�#wQ�.Ǣ9H
ҁ�nV�?}��e�M7K&� y9a�x��}��/^������co��Y\Ƹ1cY�n5/<�,%C��z�z�1{�������QM9v�tE�a��;Ѕ�TQ�����N�����Y��@�(�7	iY�����g�L���ǖ݌){�>u%V,��h�rD,��b?-���c�vM:���%z�n=z��̆���u����4�����G�m�_ϿW�F8�N��,Zp%�7}°�!��|�U=�g}|��&�B����j�j����M���A���PU�PP'9=KKK��aIЌ%�x���,I�����#O*ىb�ӻw�jj����yw�67�v	y�TT�����xٓ|�a)��$"g]���p)%�U8z섣a9���c�������K�x"&�t��XeR^2���P�f��������b���v�X�!�C8�
m�2�l��r�8b�^yo%Ɍ��<��o��ւUH)nꤷ�ኳ���P��\�a@������}���|�WG̻�D���ʵa.Y�ŷ8?��S�N!�K��h�f�A�R��+o~��7W�&��;��0G-e�#,�n6?�/�Ɔ���Lf�ׯO&N��K��Ti�Oz^�B<%������{	�F{X��X��M=
���-�����Zz��][G+[�o��+���7o%ᮄLS-R�x,G�_��h��hTJ����(��VP8�{+6S��r�J"��δt���l2s���C�lgJX-�%]���^���f��%	���q�]�	ǰX2ٸM��`��FD���E�mM��ҹ�`�4��$S8m2����U��7O�W�bBb�𕕑H�ɤr=�v�����_d���=���X�L:�S'ɝ7^C&�Ă9�s֌�t�n� (t�"<F�,Bz�w3�Ũ�;%N�}7���( DW�ɉ�]IYy~��΂E�RU[G���:r �vo�/���Cwn�D����j�bs����ˍ��y�9��#��~�x,L$%�	�U��3̴�w���N����NW$���6T/��B�/�F�27�l�H� ���ѣ������$bQ^�}��&���
���c&a�ʙW,�Tփ�nF��7���0�T٠G����&�9r����i�.<a�*>?1�;u�@|��}�[@�� �����"S���d�R�l���W��������e]5|�Ѭ\��W^|��/�M��G��W�~�7�Yp�_�����a@?to� �{���'�=r��Әu�F�c.k�[v�Dٽg�Gє����j�Omlw�-�ڿ/G��$S2Iz>SB��t�yT�|�����H�ע ?J��@u��-5��U1�6��gP��F�+f���+6��E������1G��>��%@DS�8ݐ���f6��]���,�n>�P5�>��tkj	�ͩ�Du����ԕw;��G��V�`���ln�m�0�X�f���cT��JA�Ĕ)����,��=M�`g�]����@s3��.,'C�%�ɒ�0|�H�"	�(�>�I�H�ض����Z�d1���ǌ��^��[%��e�Ӽs�����4?��;q,�t֫��U��3٤����${�1U�12"覨3e�0.8m2�޷�%7�è!"�v3���v�T!�rEY@a#�b��O�� (��ҋ"q-/�����E���x��MK�s���q>=�7�폭����:�8.��	���9#U�|�m{���ێ!��J9���4E���ni�۷� ���a����	���j��]�������nqR��岘�V��<�	��ؓ�r7VA�SU�l�̇k����i�`1L�x�9�p�lk)�sV�LN��fQ�9j�.��{�%�(���,R�Q����ج����%+_Q%���^y�b�.^�vV��Mfz*]Ġ*�(&�c`V����8��?�EI1�,���5�aΒ[h.j��"Hq�2�]�r?ܡ�����O~��{m��u�m�:��s�����Xһ(�3h��ۥYJA!*yIz�l�ֳD�d��x��S�[L��Ț ݣ�l<̻�=��s8��s6�Hn��.l���SVڅ�!&����jvH�p�gLt��ofok�3$w�V���^U�LXJf��WU���tXT2���J����Ń?��S���死Y��V2)���.L.+n�ƪ����n�#O���MQVVA)�'��J$�̕��U�~��=��ݾ�Y�����=�z���sIٍ5T�I s�݄������9��+y��gٱ�76|�-�M�2�]v��v�!��5�=���̤7��sfN���O���3p0�LV���{<�2��f0w�"f]~�*H��8�F*ӝ�.�O-&IR3)��ȧ�84V�N!�E)��gN����a�BiLz#vS�٠Xa��.S�J� ��bJ�^���n(r
!��%�LU͒ճ�ĳ�����=�����l��EE}����޻��=X<�"��B�hV��c���vʼ�|>+��>�=;����(���v!<{�6�̔d�z1�$�)`skrZ�N��@���f.��Y��n�^XU�����a��X��#b�,6w��J��i3/�����)��!��ɗҘM��N�b��e'�ӞK�6@$r�x���b�$�E���r�;pG|n^@�慳�\t+&��y\�ƟdH�hf�p,EI�Я�P�n�.͘z��ͯ�w�	9a�	��l�M�����&|�ϥsg�?��~�C?to�a�e7��ێ����9�(7F����l%gn��F�"��L<���,�h�����w�yٳ��T���P��J���믢w���q
��3ϼB{[T�'M�EMC1)�(�Y�eE�.B]���>�����N)����e��I�cW-rd�"úU&�9]V	"���o7p��w2���r~�i�_�H�� �Au���,����?����<h8�h�����s��f_ͦ�h<�A˞f�FM��w�{�C%c-YI'�23^��ʃ���[L=�,�Zv�}��;��R5*�+em�k��cfM��ң�HV���T���SW�f��O$0X�nA١���>�&޷W�Կ�GBs��N�������B�/A�0�*f�-=2Ij�R������1A����-X��z"6�;"U�#��*��B�&�d�
��ꪅ��M9��B��{�����Ϊ�t%so|�U&M;����8�cF�1�ٳ}N���������E��Y����7z�h���G�P��H���H�͈�z39=C"�$�J��-8�\+u�U���C��c�I��t�v�~��l޴��MA��.l��1��G�gwX!o� ������ J&M�E�W������d�\A'����nÛL=���.&A�31)���M<�GN�(}���+>ہ�����*��gM�x"L{4���C�z���ݡa�,$DL�Hx�q�6L��x�$��6e�{/�w����{������^x�/|ද?Z���KgMeΌ
�(QMY���Y#[H��l��Iq��V|��<��:���r��n⺛neʴc�u�9,��&���L7��3g`s����<��+��bb��aح"��� 6�F&�=�T4E���f�~؄��>��,'7�d�N���sY9"U�
�h�E���t6O���:H{4��K2t�0n��.�b׼�]f����y�[L?a2�|V��9�F�ƛ�<'�>^��)�㩬筷Wo�q�%�vp�W�����3O/'|��T2��egђ��p�x��78~�i���;,�s5��vpXY��K>��k�~���Ϳac&��QG��O����d��������-A��o��N��q?�͝�e�]@4����1i�h�d�#�tZM.�B�(R]����,� G�f��粔9����"hod@mS��a'��1�"���+�W���|�{="�dO)�jy�p4a2r���;#�d�/z���|�n;#'���_�q���ǔ��3���|��5�����Zxw��hf�|���,'O=�^=k�e�45���QU�_.
M�d�L<�%�����ew�9��PMu�]�5rt�[Ȧ�T�W[6n�̆���͔�ժ�&����CFO����NG��ȗ'��<J6�O3S�v𹈤�F�0Wr�<���Y�=���(l�}�ŒaH���\��k*��+�3j�X������À#F�T�y�^:¢h��ѻe!
�BI��)0i�4C���ڃ7]{8��O~���.�0���o�p��~٭���m¤qGpLC�cG�(��*)���WI���9���b/���dˎ<g_��'_����_�Mw,aٲ�1�,�4�D>�h5�/����/�;�|��ΰ�b��PEC��\2�"��E�j(fM�dK��/��F�fgw2�
�O=�\� J1#u�FA�Q�� �y\r���h�eظ����:©0z� �þPf�O�=r�p+�y��g����L�<��.����{�.:9�y4���v7��$9�I}^xa9�=C\;�j~X�5�\���&4�������o3���x�ͷ�i����݉צq���s���?��s�����1���k,6;#��pD�:��>z�Ts�G�ݱ��$�_��]�ys��L9cf��+�ID"�0�DE����G��nWt������?��4�!&�4S�>��%�10	Ȓ��"�f�
�( dVl��%��%]���K&2�f����6�"'=Vg%�bϿ���8����*��`�ϹgLcǦo��ܓ��?����ǟ�+�����n>�s��x\6Z����F{��AY������-�3��l�*H�ģ9�6�ӭ$Y�D������H��1�Kv�^� ���,6&��UD���r�Ћ)9�WY���J��M�=��{�>���%�	0?[����/ll�W��3�C�U|�ط�2i��Ȣ���Ï�0a�H��}��\���<���9p�l>�Ⱦ��e�+_�E
%��ơv�iS&�x��9�ɏ�×wx�~h?s�X���GƏܗy��/�f�I)�؅7����h�eݱ���_w���M�~9!!    IDAT��n�'O����8��í7�"3�W�x�p<���F&?�k��g���RI�B����b�u��e2�q�,�,�����,i+C����>���߳;�\Q�hf�Ѥ�	\�B���66����� س/�R	��&�,��,��9�8�kho>�{O>��睍��t��9u�̷޿g/���w7s�W�7c�o�kle�q�p*%>Z�6��A���A���b��6Q^�5嶻��s.��ݷ����0����% G�m�ҷ}��T�;�ﯕ{�!=�1�7/.�i�M6���R�͗����!�)���p鼅d�.2�*�Ndu���������X"��n�vxK'S����fΝ9�1܌d'���V�<u̚���Z�����Ԥ嫰z�d1;e�P�K�%5�� t�4h%�q�=�`�;E4G�D��bȪ��Q�wϿ����|6ͬӧ���W��%r��٧k�.��& ��z>��f%��ѣ.De��L>B8�&�U�K��IkT=/��G�3*F�b��H��Fc��c[6o�n�`�9)Lr�ಫ���	�1fҩ̻�i�v�ș<d���P�`�9��V��.�v�mm$�)������IF�4�T/�"B��xn������9����o�lZ����7��w<�cO���N����p�w3w�R���Oe%��PU<��s �r��Pհ�K�Xf攉��k���!|�����?�m߬Y�w��3�0�����V����DO�$x�8�(F��tV�R�m;�x���5��������^�w���^��VVV#u��6�R (��L"N�mg�Q�%�J̈��Q��Y���NX��@2gPV�KN��P�sr�������e�!���4(1J9"nm��Ӗ���r��z��g�˚�6�b��	��P����/^~��N8�X&Ʋ�n��g���s��1��#,��!Ɵp*ކ�|��WD��tֹ$���x�{��<��}G�ǁ={��k ���?��o��!�������w�z���`��Q,��6��3�L�}9�܋�p���v:�x�q,V�z�`Xߞ���r.>g&�\��}(;���L?�|k9|�'�uf��D����!�،����<@�
�b�薒����(��@2�m�s����>w՞Nj�M�
�r+V,[~��nqOm�8V
2���խKׄ[� �"��N>gE��	�|�-=���,�8��K���;�61a������~��9v��X��_}95^v���o���a�0	� ���&����]-��(ᰙ	U{i�YI]����5)ta�&�e�"E���od��]l޴���Vҙ���]n��	��"��Lyy WY�������n�)��&���J��Vj��v-a9�]v>/8'NY�	���$�� �,v��1�b�1l�0���+��rP]ӓL����C�輿��[n抹��o�Q�M8��vrT�� ���n�Gd����n@�<��r�y���v����a@?��w,���-m㏟8�Eg�Ēي��T�H�Vq�-��a�_�^�]Fy�?�m�Йr��G��t�Tҙ$kWl�t`w�	]�%�H�I�Ȧ�Tz]9b �RS� egEE�,���y9��}�:����C���젪<���Z�<vy�R�.��;O��'2$�
�m�I�j%У/y[9��p��ij�]����Ъ��F:y��e,�}){wrӢ9��5�V�|�7���`Б�ɻ<���DKG���~���e��k�w��qةo���w?����xb�s�:�r*�ըf�H T@��{�����t��f#G�{���J����З\�H��l��ݗ�bH�
���T�����	OY�~�=bYO��.�_���É�t��f)$�h�$�Ab�<��NA��00r���G1���SL%9�䣘q� ��*�V~�cϐ�	���]��ٷ����$P�GCYw����R4kI���w� �|�C6�����}�ӫ
����c�v�b/�[��QG���mX��
�ͬs�c���7��ʋ�����ߐ��$�qs�]��cӜ��Vr�n�]��QR�����D6�EuR*u�ĳ������9��,���dZ�,��]D�J{XM����T��˂ؼ<u��z�h��	���Řر��">�J�C�n5�vK*�Az�H��.���3g�Ncc#7n��.��3f̠���+V�k�N�n�l�����s%T�_�f����Gk����Nw" �_��륐)�D?ݬbŖ`�O���7_{x�~����K<��͟����>��#Ϙz4�NB��'l��b���
&�j�޽�#A3��*�t셫�>Dm�1|�������\�"��F/�8��38�)\q�%��Q#]��+82z��Q �K���Ύ�w���}�Q���^s5�~?��w.=jj�A(�)\n�L�{��w�����ǟ�ԋ/������͏ݰѾ�R�fB	�)�����IN�����"<j�BN���_w���0�7`
Tʈ�\"I��[��&ȃj��ￍT�U&w�/��6�D'g��܂��g��f��N�}	%!�R̸�̾���~O9��:0��wEHw�`7R]y�o��E �%�c+V3<��2��ɘLd
y�^��va�B�
b��T�-���!��0�{���v�Y��b�`Nu/N5�Ihؓvmkf��tt�S�1|D̊X���,&�jA���ê��v����D��u
-U��N�X)*�ذ)B�T��]�ߗ�&��Ŵf��+��:ԯ�X��}v�mE��k�,{]��R��(��u�Բ�׆�i���BV��\�D<�͔�=%3�j'�d����Yvi�*�7���8��Q-N�� }�Ɍ��E��E�EԊ��9�N��Q�H�aWW1�A1b_n��e� ���a��}�w����z;�֭�ӈ����{�-�y�f��@e{�c�3�tRx���*k(�]�Hkm�S	M�To��TG�p.��ӏ?���8����|�����tÖ	�>�K&����)&P��R;+�PĘVS�l#�ߢ#o���_���_�T5T��)d��V���Yᖥ)�	�;�E�_��O�Ygr���i���1�]D^fS�.�v;������{\��q�?$��e����q9�ح�27i�y`?�u�ضs��{9K�Z�+k>��O�h�i�N�������)�P.fJ�0&�̽�\j�r�I���-��v'w=Ċ&�"�;�ř��5��3�<��~l��Vvp�#O���[|8�U��mً��*w�x�x"MsX���r
�ʾ(U���ڕOݿ�r�A�M�;���u�bQ4w%�=��������YQ�I��T1��!�Ĕ��)����LQ��c�s&6v��hsdS����Y�9vd/�uA�=��؄Uɐ��3���f�	Y�h����MT�̂/b�l�lh�3l�,��{�s�V]�"�@?���*F9����}�?,���@��M)�dܘA�W�2����=�a��n�:N�S&�YT+�l�p��p���.��� G�SM0ntwȆ�.��
bw��e2�9p@��9���	Vֲl�#�u3-I���444p�Uc��Ŵ��`�JG?1ʗ�q!K�o���#�r��\��Ȧ2ilV�,�E0�QG%%l=���W^�����	���h�/^���˻�J:��d�>A�T�P"�Ձ�jCu8P�R�J:+�J��U�J$C�;�[�z����w-��?���?ܡ��o�`�ϻ��o�o�~�%gǕ���;Ŭ�X<.cM�l
�Sq�p�]2;�(�M<�Ŝ�����~���]D�>��D����K��rzA��N8n�M�=����#�`�q��l**�
U���7�ѱ�����?�Au�M7I����/;���<���ZI��r��s9y���9~��g>]�%���O����vwR���m���RB�Χ���(�j$��&���,Yp�RF>���廍����YBxB}�iv�V�����¿����c�/�m�V$�<�����������1�_ov�����&�k�棘MX����rr�S�'�r݀�%��	�t��A;K^��]�Q����#o�c_� w�`=%�'w�^k��Ɲ2)z��O�PI�M�Yz��Ck{��@�I_!�B��>�7s/?��O?�#�2��,���;dי��$J52'^t�h6��&F�%���)�CA7��ktE2�l�s����x�j������a��x�?�P��T(ѷg�����ee
��2��*�d'Z���?�ć�}���eܘQ4��U�6��وF�R�!��.�Ϧ@��#
a���Dhi��m�^�563h�p��:��=1�<���;�xl]����l�c�9���]ω'���)���H�D��H��S�m�t��Akk�m���_��Kz}�,?��c���лOٙϟ?�>��MM\~��<��t��a���8�M��
f	��>X�@4�-��q�Z"#'@ZyE�*��Ӝ����>~��O޹��?��v�����g@����s�u��>o�Df�Ա�;��߶�x��\.��a��g��{��U�
�
���)�{p���y��wX��7���&n��nN>�|���"84+yF�)�޷-��	cF��GϺZ�N1��6�WBJ�U����[�~�]ˤ�ל�s%cx㨭�¢�0]���"a)�Ɠx<>^{�Mz�a������7���K�c6��Tɑ�̗ξ��z�Ύ0󯽈��
-{~�b��a�V���J�7�P� ���R%�Q#�2������ �N��Kӎ��w�be�`	�3o���r����x�����m��k�@�Sd�IR���_MQ�1���x惯$8ѻ��=jx�g��pq���9��7H'�U�����a��~�m�[r5�Q2cQ2d��r�^UWKN�K�	x�e����u�T�t���&r�4W^u	'=�'��݄CKp��9q�:Z�%(��� �Tn�]��E�RM��2��ɬ��ps{
�d��ZNm� *�zq����g�����`[3�߰ �ņ��A�䱫vR����,�q������w�	��I�V���)���޳Wա**�!م[�6PJdsI��[ٽk�MʹR��Ŵ�g0�c�U�O�0Y�lܲ��/���^����=���A��Ü9s���+H�%
���X����SA3r=6)c�(�|F��(��ʵ���3�=zp�i�q��E���=�o�z��hh��+��Y����s�u��)ѳ����V�A,�>�[z"�KI@�V��K�k@�Z(��S��C�:q��O�y�ه�iw��w��30�>�����͜�5'��E�cq6���/����5ҿO�lNn+y�%�t9������_��`܄q|�f-�`[v5��*��TH��Kг.���?�Θ1���]t�7S]Q�����0˃�<d�#��륯�˯���[�s�]wKW�N��5�\��i�����~�U��C�5TWW���m̞=��~�97�E�l ����H��BFWp��$$�x����os��|̹�|lF3�h+��r֬��?��cN��j����?S�T������{��aܸhׯ#������9�ēQ�A^_�1SO=�{ﻇ�|��>Y�C�����%��I'������3h�x^X�%9����j��ewK�X��u6��5��f&L����u^��^{�#f]<G�?�b'�����(��`9Q��㯐ni�7��R_Q�9���q/bB>r�p&�e��(U�v�%��+C��0��)<��1�͜8��.W�ghli�N�>�FXĔ�u��ʱ�5�i����ǟ���(�R]ӗX*OK['[��ƅ�]ȸ�c��^<#��d�bN'�ODط��~�*��=6\N�a�ii6�ƾ��ٹ�w�2mo���[�њm*�lZ#����?��Ï����9�{9��y���} B�~#1Y�2�M���p�)��ٵ��];W���J�d��m*��B���C���.:t�,be��x_���2�<�L֯_ώ;����k���3�0j�(�y�]9f�����]��$����LK�z�BG/� V����0%*���USGA1K_�^S�N,��S���c�Xp�!p����,�C�X��΍o�4b��q\5�M�}'�b9k?���p�d5�ng�9�٢H��bq�������/}�7�M�޽p�*X��:���ր�-����ZcȀ:.��|�]}�L�9=�m[7q�3(�:�d��`���:��4�_LSK;��_���g�IN׹�+�?�'N>���h�Y2�CU�|�r�|������_��naCx���� #�FM6��$z���^~���\C$U"p1�����)�˯[�u��������ٗ^#PU�q����e��������`��}��m�f�Y�!���;���3�7w�^_���d�x��2z�v��,_�4}{�����,{�YLBf��8�SX�Ŀ�T���>HFd��{�m{[����򺥤�
r��M#렐�P^�k��'Me�����m1�jm%�J "Tʫ�$\��s�����	��'k>&�QS��gg�PmN�z�yg3v���z🧖��*���'��v��9��3�S������;R�<�'���w����.��uY��m&v��������k*C�ʤ{�܇E�	�������m�i��Bȭ��!�L���n7H��2�Ld�o�}w.Jfk ��##KE0@��=t�wH���hh�2����.�d��I�N���g��N;�Na�X�Z5�;2�{ｗ/��&bWL�:�x*I}}=�z��FC�׋/�(Q������,����)�$����]���mR�':t���Z	�bU&��&�M��@�9��/���~������?��;~��-�Ϙ>��gVS�܎͍"T8se�Ѭ�+��.X���O[��D�˜��p��O�܋/���;g!�w
w%�����$n���d�Ё,^���P˖�Lφzz6�%��+sI�٬2m�b7��q��뤱��7�����9�̳Y��c&�ƌ����f��'�`��s�%���Y���<��J�X�<!�!?�R���T4�ߢ�i?ȧ�Ȣ���`��C�R�]W�]�vKy���&ƌO2���%�Z�>c���|���Pӣ�PE�4��lm!�NK&�J<���̺�
^y�E��f~��$I	��~}����}�}�*��;�{}�h2�ؑ�9�,�{N�o�OM��j���[6I괅�|��wL>�<��@�F�o@��s!-�ۮP-�\Q�JE��Iϧ)�E|h'��G��V��E!/s�I���T�TSA��s3�L�b�K&�勂na�?G m"��A��G1i�V��'�V9Nȶ����)v���o���璸]��4nO����� ���a]��zFD�
�y:�I6х��f�I��˄	<��S�3>c�Y��e+;�6S��d��	B�г:͍M$�E��}<%��N�(3x=6�]��y]�sYi c�B�E�ʑ�*�^
	�e;M�ϲ�*��'�G ���|�����PQQ!��`K�ԟ;~��G9����_U��lk�I@z2.\�t~?%�CF�Z�Yi�#v��aQLb�NyCy��O9��o�s�!p�������,��o���y���j���a�#[�
�Q�(ܫ]ʗ0�Ĩ�Iыv��M&Z�T���V�?�
�DUMe�j.�j.��\J�Db��ia���㶛�>�d�ψQ���l��	J�R"���M&������g���hjf���rW>i��̛$�������Ɵ���5���S�8(��;}��,��>���$��}g��D���۾4����X�����q���j�ZYP4�y��ӦK��o���:;n$��T��+��NU�C�~��b6�ɧN���Ob2)���JN9}K�,a�7����52����g��m8a���FJ���x|��x�~��q�̓��楄��8vʉX5ѿ�D��g_x�}Mm���'�u�\,�I�Dd�A6څ��b�[1�+��$M�r���b8��{{�$�e3._@(�)
EUA��X�g{�;�$�Ma�[0�YF�R1Gg4!���b��MIQ�XlҵO�K���	�1��]M�ݤH3�=@�    IDATkN�[fϻ��ڛ���Ţ`��19�h��-�~�-��vEt�J�b6N:��QGc�U���g�a�u�qۭL�q
;���^�_���#�E�f���1K�T�l�LV(2l�TMz���,J�=#�190Y��Egl��ی<A��]C���[8�	%�������źHL)�^��(��T�K�L���#Vb�$8	B���ǎ��t���.������vɈckJ|��,�nR$��#w39	�g�t��-���C��;|�;�C�Xp�]�~�u���O�<kz;F�E�Z-B����&r"2S�KR֊�V�}�ɨ1�p��E�z��;�X4���}��Mmt;�Սa	���.ȃ����3Ϡ��O*Ӊ��XPd�G����m�)��e�$:-\r#v���.�T�6����cǌ�Y�n��Ͽ�T�*eT�������W�]×�6��!�4�N�d��E�[s>�+���Σ�#��T�X�Q*dp�\�cq�{6p�ig��켿j-m�$SO��Ǟ��".eCfT�۱N�p;���kX�ҫ7�t�.����|���Z��떦.�/�����t��2��������ı��� /���^Cׁ?x����;\ĳ���7��v&��]qH�a��G6��f�QUOg"�IH-�����C<*IU��@e5�t��It��)����&j=)w��d���8��ߘ4b�(j!'�T�*(
���t��$�	�ʤD��Ev��dF�zw��!�R����.�J���=h�2r(�t��\ds�6'�B	SI�k��I��2��ξ�9W_��իx���9�����#h�z��JTo��^ U����:VE����{ϩ�`�<F�(	o�X���.%�C����1���',��e.+����Fgg��ob�!�K��BS\��<rz^^� }э��f�Ν��)V�K~�������(�� ���)�p���z*������*�М.�C��젼�V���,�9��c��l����#��%���g��{��\����g�u"��TZ�8z\%��A��t<��pVU��p�cPƽ��Ć_��_���Ϳ�7�]Ɍ3���Xy���8~�)��5�d�,l8�Yf�8�3O;���Ȏ,�	K�P�����.�({!�� �P9��\rٕ���Y����?؈U����J���C0���=n2ٔ<L��*H�<��;����|��n�f�����(bRu��4�x+W<GM�KAtS^��V��uU!v�ه3X�����O�i�^rEcF�5�̠" :�.I
�UUKs�A�e,���0]�4Kn_�ٳ��'�Yؽ{'��\"BgG���cq��$����w?��b��i�헞d믿QUU�ju	�Ӳ�w��%zOS钙�w<Hvo�L�%Com�9���	�rJ&銦Y=K1#��P&~�����a��$�옅�N&�X���^�DDz����;[��I��_/R��'��$S]r$l���Z<RN&���+�ўy=#���յ2%ܕ��:�'���
��~�NNX��44�"�L�d`��B����T��ܸ�:jB�v��L?�$Ǝμ��8�p{Ȏ�3���u��5�6V�D�E>�¢�P�"�|RN�y��a�M�l�������3�j�kR*Ih�KQ�$�"%[D��V�5�J�E��E�B�N�/c̾�}?���_����]����5׌1f�}�����~��E���k"x����Q:=fG��G�,"�2Sd&ە��7��nڴi��ˊ��mۦ&�a#��b���o��������{�q��1�{����ٶc��Х��}Q�F=�������.����Q�����d0S�Q�����X�ZA��g��+�6�ׁ{`�wV�:W605#�~w_G}g%-�{хJф�d��*�1����Z.\��r[��Nf��s<z�5?l`��s���3��I�u�=htI�V"83��ya4�Z���_�@�ZeMuv***q:�
S�4!0�ZJ*KY���\��Z���3����P��$�]M�EWԴ/ӯ?ę�Me>��Nc����h�M�-Z\�
��3�����P?���aCX�f%��gꔉ<t����3j�$�Y^��):/%�.��ҥ+4iЈ�?Ŗ�~f�?��h�#|�շ�4�o0D�Iˋ/<��FF���wv��铬��3�zX��˾]K�:㒜�xWI>�IF��*B1=����Z���t�ы��lV����%�����S��g�f�3��(��Q�	�����
|y�X�o�������7�������v�{�8v�w�ёӧ����
�6Ė���i�_������iiܠ�b�_)8�o5�ωc�ɫ�N�_��L��u�sg�ٻ� �V�W�NQ��j5Ңes�?HZF=2�r9y���� ������քVIkK�	�k ����$�<<�`w�n����]wv����];������S�hs��Դl�k�{�<^2R�\>O�ì|��~�nK�i�QQr�ߵ�D��љ�����fG�)B���51*�*d.f6�ǏW܎�c���/2�|�صS��E�.���x����7o�"|
In�ȑ<?b8m����҈rؓ��4������l-f��6L>�ڔ4%[��.���⤠�����~��3'�x�i�.�ڄ^w���O��j���,?ƺ��JN�bO��	q��1n���Ӣ��_z��;�b05�l�&����3.����_XD"!��:�4j�,`O<:��%@C���D̨��]m�d4Ek��J����Q�������i�$%+R��H��� �>��׀����lD�&iN�����q���X��D�TAI��5��篗�t�BÞ���W2s�\��z���Df5�G�?�Β�6������o���Mt���,�O��8w��;u�^Fg2��Oyo�LF����^��~���m�k�>f�"��?u�/7��Κ�!!TU��?����8l�}���O୷g�l�����&�Og��;����?�]d��,�`!52uc�=>R3�	�ʲ4�_v�믿N�zв͍��ȯ[���k���(Sy�Y�idg�r�����?��}ƌǕr}�>JӜL�,��]�����Bȁ>222����cO�bUUUÂ�p�|�^���9���O@�ª�k���n���]M�Z��xԇ�o#7�iEVz�P�KVI*dEV$���*8���2i�jMT^�!95�-�~����)q�(�X�'��رcس�7�6�C$�Ӿx��;;�����D�\����o�����Ђ���%��#~U�3�ڂ^Q��Bt����,]������+c�U��޷o_5���+�s�ؗ/_���g�y��S&Ӱ�/�M1$b��n.�ш�� 
��h߀%;W��5�Z�A��tQ�C�{��&WwO�kW~mB������f�r�l"�t�%�D+���K��|kv����>\J0�UZzv��������}�_���S�/���`Щ���C���+NI�JMXُ͚����Q��m�b����j�fe�FBaL}b5j�ݳG���2��gK+߳�%S�	��Hn�<�ф���f*.B� I�u�yU�Z�w4�v�΀���B���پ�7{�/k�]·/f���D�e�6�g��ÒSIk�i�̝9��^�����c�9(+�&59���.���U��/gշ_��������F^{�5��5���ᆛn��}1���h-I	��&V.�G��eێ}� �咅Lzy����v�X�y'�"�L��#����ϩ�t�w��g���i|�d�k���C��T�BB6�����ыV7܈���o����އA'73S���VU����(*.f��7�N_,�!�Qx�kW�TE���*f����~��%4jB��=��؟J1��6�q�����vj]�EHNM���s\)f׮��~�1j\~���2�4n�A�뚨��p@V	Fn��vR2�ƵVTѰA.	5'�PE�n��r����^�H"�U9�n��Q�_�̙Sl��#�W1��4P�}Ea1	б�:b$.�Kr&�`D1�����N���ĕ�,�Ү�������?н{w�����֛��>x�`�f9p� �ϟW?��'Oү_?���[�7��������).��*R��ք�����g���e�ר�Bk�(c)��{�3��a/Ձ#��%^����=0�݅o�?Q�ZuĈCgD�)#Zz�f�%�"DAa9>��HL��S����P:qq��lܴZ�]%+=��$�mh�6��ؒ�N6�	KT3&�C%s�c���P�ɬ�<
�h�jW(�*�6���D�#�>����U����2I��XE~�]O�H�4*�s�h���6�\#r�PH�uf���!��f"e%��l1[7��o�~��Ճ��NVP�ޒ��Sgy�ɾ<���h��#Ay�Þ�ýeޜ����/�a�h��m���G�֫�:�&M������t�֍�����]M��6o��]�M�~������H(H���M+?�ܩ�2u����z/�π���^:�ѝ�G��^���s�E�>�����D�����0�u{�};w��3�X��;E�����|��w��?�7܈���-?�@�;o#�捉/���*��ѿqd����=���K}�)GO\���è,��w+>'3+��/����և����@$΋c����WHNMQ��7�2|�r��Y�`.?m�D��0Y�l��#������x��Q*W���4v����d�4��҅��8q�#�.p�J�̆����t��QE�m��d�:�ۻ�UU;�7e�.��u��VG��=).������l�N�v�n���R�eƌ�#9�g��۳��̨OD�#�РID0DBd��U��6��R�ףt�ܙ����Ox�ؼy���N����~�S�ӧOs��aU쥸������+�L��N]�s�T�ܓ�9-+U֯"[��M��5��}*�8OH$�u�G������^w�yu��&�:pL��x���Ͻ��[�B�v���qJ���E<� ��@��Հ���H���\ٵ�CnUxu;f��P�6�$��;�*�E����ګۜU�����j���"
*����P�eMe�2by�p)�F��p0��Fq�
�"$�g�$)]q�pT5r��b**3��0��q5�D�q����4�1��Xg�}شmE����r)nW���?���?RTVNB����j���	��D�����ӧX�~+�Q1��׬#���E���z�7l���<��`�����v��ݻ���ª�?����k�[�
x����]��䬖��1Z4���߇�ܩ#�Z�e��}T��x&�8%%�x�γd�[<��S<гi�ɴhP����͉3�Պo�r��qS^g��Shڪ�����~-O�C�EKۦ�4��PD���TA)���-o��_������@U1�|�)w�s;񈛖MsHMJ��}�)(�$�~SF�σ�����A4b��	̝5��om���&M�@n�l6o��m;~��ߧ�TP�흻���V��6ױ~�r*�
x�L�����L��.k~�{v���%b�<��J.�v��%�Y��������X���Jj����Gw%s,/. �abλ3��￉`dч�,$:���_aʛ��XRU�4��st� 9i��&%c��!�N��T��1c�0m�4fϞ��� ={>��q!�	�.q��B�dZ�ን�S\\c�W]��(�,(,w��IAR��`R��d'
K��Nq���{�	�'ԁ#��%^����=0nڂ�Ϟ�[�A�~%j|������<eD�	[U�é��QVd>ژ���R�� &�u�����֠�;$�M�v�Q{�6���0�Eh��(��Q�P�g,V�NZ�N��� C�ҥ���-&��팵{8�=9���z�#q�<陊�p{�[�H� �����^o����h�ϯ4�&-TՔb�S�Ή"΀Ř�P���H�}�jLL�(�p�-C�^W>��5S�D��79��9IQ�q��Ju�[��"��Z�H,���)&����L<C�`�U���Ky�����QZMD��$/>���Dl����"A��ъ�|q_�]:2r�`��v+��8��nf���,^��M����!�I�k���gX��2Ǝ���1b�4�J������<��o�c���jB�t���O�"�,�����<���6�5HS�Ņ�����(U� �ƿ�Ӄ�����A�c�Kc���<��!�^߂��{+HZ$^?l������y�N�4�� ���=�3��W!�V}M�6�Q�V<��p�8|���ȯ����pZ�ث�IJ�y�Q��љ�W,�~�\:u��7�6�Μ�Ì��2����v�i�,��n��Fl�il���Jts8�yi�Tƽ�iZ�������G��Kw*�>U��D"��e/��^�\/Y���y���W�V]��"[K�Q:)��^�Д���U���mEW
�'�1'%6��*����S���P]�y��������e��k;��{�_����s���_�p�܂�X����c�3����ƙ��#��*O��-U:�/��t�˖j�v��t�	
3�R�)]ZZ��a"--�Ѧv�z����4�+ܪ@;�m
2ٚ��|^���iOb���d�婠��l֤)&���e�!�:u
�3���\.�_&%+�3���*eV�0�	�ϫ���*���%/<5�;B�%#Iv�q\�%$';�&Y�T���b�aO����3����~"� 1�O@��1�;ވA��䦛{���Ji嵺�B."�R�H(G1��D��å�W� �GJ�b�G\5U؜��ב�(��r�|/�)D0���[R09)
�Ռ.��r���Q�9���^9��$3�H�8	���3g��I���U�K<e�����]�mހ'{�GV����pB���������,��kv8��^�u��.��Cta��g0�'9-��E,�vǎ�f�˯�҄WT�&&4/�Ô)�x�띌3R�Is'�˗_~�Ɵ��b����VbOMV��О	cGҴA^~�#G��U�W����`o|~��8�%d�k��*=�	�ܗ�7�e��?y{�,f��!߮�LqY%����B�{��w�<'��]�&��QPXĸ����}�i>_�sJ���k�Ft�t���Ms��.�xq�nH8,&9F��=��=d�`5����e�g�gѲ�u�8v�@X��Z��Uմjہ�gKW"�l���_8HRvz�]9j�2��1fd�0�����H�A�|�E��h��͝2jt�8ծ]�����ׁ�����z�`�5%���άW&�.�TS��H���A��,�6�A/*1��T-���r���V�fI�R6�f�򨾻KW6n��4�.�i��VV�N���T���hPdD����tR�M�F�KS f'I�z�D�a�4�`X�`Lt���d�����9�^!?iٙT�x�AŒ��h�(f�|�>�ћ��M�R�Lur�Rٴ�{U�qW��\�L���������0a�8�%��hMq�Z>e��G�s��E&LxYEfFcA�̛Gn^=k*!3�/_a��w	b�5㰘��ig�;o(ƶ0��8;��c���Č������㠷���Q��)�t��$׷h��74��Щ�u�����s�;$�͆V�ǪOp��~:�nB�U�&�S;��g�SP^ŹK�X�hm��
q�������*+�N��}�N"Ҥ�u�c2%����1L$��`�����<v��<ξ}���x�&��:�OĜ�?�%řL��Ms�<n8Vk�޽�����v���&��>�1�!�zG*�P [M��8v�Ȅ�#شa=��;3g�֌�l޺�ʊjzv���"��C���̞<�����U���X��;1O<7���#��`T��8�D��4vSBy��B
�.�����7�&7--���2��H\幇꽐@e� ���5ٜ*_>�q+NT(��]������ɨ�����x1�$Р�os#��lKe%>��rhW3��=�Ϝ4�l�����K�V����?s��ѫ��~_���e�qU֨=^8'!@�u\
v�X
��4���YX���MyPkuj'��9w)��E���HL�x�_$��hR6�Z�^hٍk�h�ŕ\Mc0��D+�;��=�ڣ���&�P�v�5�&�bJ�6���X    IDAT&!�:f2�_�pt�j �!I��x,����谘��j�#�Wi3��%Ӻq=���XX�g	�9�)΀��ʮ�Ŕي��Y�Dc1�^ai��{��A�s�N,Y�1ZC���~�.]�p��	��T�˪x���Lw.�~�nܯ$Q�6��fLPQ^���#�1����R�%���[	��f6)u�ـ��
���&L�&yt���jZ��c-�o�w��#�w`Ϲ���F\���{<@�T���;;�¥q��i
˪1;Rpf7��qb����O9��i�)�����/�c���(��"�b0ڕ�@��f3����.�٢�avy��������3e��Ty�DE���4�L��[�p�.�ж	�=�,��6[R6o�����X�$�ᒤ7ȧ<�����.��<�_����{ye�$f�[����RU�&�i�Z�l�
�1������`a�כ)q�1$gS��b��%�Ѣ� �����P='7�@ ���H�KB����2�X\�¡�Z1ɛ�Ǫ	g9ijmfu��<j<a�����B	����&d4cNr`7[��"#��NX���k�J��5�UAwD\�qϼw&}�i�.�����o�]0n����W3������%uC�|���D�����d�b#5,�ZY*��X�o�	�o8F�_�2���(S	���рQ�hm"�U&�V#�2��UX��G	t)�R~���Ҁ���W?���Xm�C�������y��sÉ�j�8���T+]~:�b�41l�(ao��Sh���a�	x<�*r�4.B̓ݾ�>_��λ�R�㒍-�貏��������	�ԫ��������e<��A:r����`�'ѰqN�:�ݤa�7x��^��o6���7�-��d"Z3�b��7)����4�0��M�K�����DV�]��j0���ͧ_~NPc!a�O0��h3�z\4�r`҅��}��˥�m�v��\>�\��5ǣKV�L��"v*��e�*4Gv�6m�����K�ĴF�z!>��"EY�jqno��L�0�gOs���<p�/�''9-�ތM��������}h�4�=���Ң��<�Rw�ـ��$7`�jщ[����t�/Y��}����̜7��s�Ǯ㔗U�b6�_pC��D��;/�B���Gu|��.V#��	�sz�`m\�Y�UMS�MGf��#/���������T�o)�B��n6׆��cQu�HA��Y��J�Rs(��2�㥸}!U�.B�
�KR]Mq��IF=E��f�>�*m����nw-�5������X�u�e��q�.��g������|0�5�n��������QX2���be�i4����������֘p��r�[nc�[j�qƵ��T��dB��t
��B�M�|S��-�{Bb"�'���O5	y��ZT!���Z�٘"ę����<k�$�E�
�W�;�3���p��I�!�#�i�yn�2qHR��oո�.��bz"�����AL���v�x����EU�o�|��g���*^��o�Q�4�ٿ� �3��I�˭ ��t'��z�NzY5�Y�)����g�XTE\k�l%�V=�B�34<�p7~X�-���4��$�`��C�:�u<5�y.��������&eன������ן��i=�	/�;ݢ���U?l����AC���(i��6��9���;y��;()�H��9���{(*.'I��~|��*b	�*L�;�租��{���I�<�W�OYU%{��Ee���O?�7߮�`�)�N7�f���XF�I�^���0�~jE5��R�[��rUa3B� b@��zN>Y4��kV)�������i�_�;u���pć'�&5����Ԩd�h�ė�7P\�����NH�O5��$"�	{h���E�o�^*�U�&Y�����}m�J-�a�{C�y���+�TH#�Rqa�G)��ܻK>�`ub��)/� �Б�[�^���#A1�S�*�1����l6�	`�WЧkǏ����:q�]����#pr�7��sǭ?q�=�pmX4�y�O���\A�n��Ք��}�jWEU&������+�[>Q|���y��k�p���-�LD'y�0�Mz%͑���� �1�P.\R�#* CHB2I�'��b1G��V �h���8�D�쯥��n_#�/r�
��tL�k���zq�����J"�-�3�p�.N�_C�QC��Lۦ�	Ք�`M���,�W Vӿ���q !Li��бcg���Jrw��Q�0�y�f��{T��;�Y&��/M`��e���� �i2Y�Ѫy3�8�h�'h�V�<�4/�:�]{���'���F���J�����|�t1��M��qc����=U�ף����_}ʹ����WH���SS��߷�D�Ghۺ%%g��,"=9�6:�d����̘=��O���e����B6�\N���Pt�j��� u&�����ǌc��qL�� ��x�צN���]�t�8�P����Z�l�q��QΜ9K��j�4ڢa#G�����?�������1x�Pʫjx♧ٽ� ��^��H�������	�>��w�}�v�o�x���}ˆ��	�⤉ul�K�����Z���[�Ք�h���<|����Ӵ%�K�	�M�T�l���C#�a��(�jj:��/)[�^�je��ו�T�Y
{�U�ɼv����LQ�����p	�S\r�C#`����K L$�#��c�m�Fo��
�1$9Մn���ۖ,��Ұ:p�]��k�{ݽ��[4b��S��w�{3�d�4�U�Z�n$��߽y����.���f�ګ{u)b�'�Z0ڒ8y���ށ?nU��l#)-]�ϒ�%�m)Вb%�B��M����G��,�����贄bq4&�h��h�uZ��*��a��!	���'�F\�섀�
DH����"Q1����#!������ �#	ɺ6hH�h�(����NR�Db�o�)�`$���\�"���ڑz$��JFz*_��H4D�&�2d��k��M7�¾���:B�,!�ɵ4oޜ�n�|�e*�AR�p&�O�"VXZ�t�V�h�c��˙9y<3�x��������0�*C��q��9�|�˾Yó�'���IyI>߭X�ȡ��(/�1c�(׀��`��'K����Y�z�|��ߎ�g�c��|�o>�����#�'���\���g�:}&OEfv=4�0s�}���@�^=��a���j�*����V�l�����<7�|a�qG�v�9�'9z�z���MZ�ႏ�"��iV���~��~}e���|��cƎy��{wg���9u�47�����ΰz��a#�����?�f�S����FX�Z*|~R3�������i�L��K���%#D��=>̱�3���1z���̜l�ѐ����j��>X���L�*]M����"�e��Ңr�V�S;�ǏW���f)�j���C4�܆�L6���BjԢ�a	T���^+�u��WW~mB�7��w�<��|�gR�d��d�tU�ej����}��suW}u"�)��.��C��r��D�A�ՙ��3��j�h-��?7���hBT�jծ\����4��+�VX�t����-v��)n��qG�j�F�A�A��ъ�5qܞJ�;��uxF5:�c�@HeB��i�h�>�a�j�q�3���d����!;�J��t��*�g��M�%3I1W�r�[���Z΁VoTY�����e�*����CJ�&^�!�������ŋ��/�<)�6"S�X�*��ʕ
�I#KFoM&�������ύ>fʋØ5mY��]�{?��2����f-�g������&�:K��|��s�:�وͬ��mmi׶[~���_#��2�V�a����z���%�b���4o�G�F�U���+WX�f����՚Ƙ�Sx~�x22����_0��c����.�\8ǫ�'q��%�v��Q�ʪرc7��{RI����%Kr��1�ӋV�@vF6_|�%��cŚ�H��ą�,Y��G��?��>��"�a#Z���?m�^^�����d���q��?l޹�;:�B�>ʝo#b�s!��];����|�1����J1Ʌ ���N�;͐�l��Cݔ}�˥�B��b.�KZrZm4�٬P)�'���T�����Ev������2�}�}��$�����0ڝJ�y����1`��#.,�D-jd0[�����t��fLQ��k�xmB����[s�����	�����bь��./��e��Ϯ��e��}�2���T!�79��k$>T�������3�"ZlI��ufB�	�� Q�Z�C�$��M�jJ�� e?Qr8)�1���N왙T�z\��2�G<n��.�����^����Q@JNn�X
��'� �F��)I�NoTs��Q�����ɱU�<|�U�8�����+�>9�����o�%��,:�4���.?SUU�&{�~��'r&�>��߽�������}$%%)��/ Zc�Ҵ�u<?j��Ƒg�&�)�F�Sρ�qU�Ӻt��r4�����G�c��׸�i����}'N�������d7mN�œ9|���P^Z�#�O�&8�o77���M�6q��9�þ��ݜ(t�XX�E�~���~}z�)�����&���ѨA+���SCG�p�tyy���,���5m@����
����o���Sg.p��9���n�A��$�z����]:�m�V���kd呙����3hu�uL?�%-�g�^��pKR]8̼>!�QD��m��&��e��<������뚱�m82�hѪ-G����gx~��O}S�wv�Ӛ�:��dF���r����~�f�j�)h]�1cR���c�"����ZU�����ua6Y���RZ�f��Mx�~Om�թ"\%�@���F�iل$�H�_Ebj�`����[��K�̞2��t׮�ڄ^�,|b�ѳ�
���G�l��J��x��+�����+��8��d!ӸF2�K������']�l�Vϥ˅<1pk6l��܅9%���%�%7u�I�Fh=	�e��}�8���S��]���Z}��Rq�c$,V24"a���JBn�` ]<���6�S�Wk֮�dMR>�I�T�D�T��UcHD�ܴj�Bi��_��ACLi���fR/'S��z���堖�M�m�A\�"�� '��f3�9����˼>��*�N���s�1���l�m�vU�9�T��J+/�2)�2�_��YmI���."q�~܊��Dg4"U$�&�P��Es_c���d�6�U˦thی���F�9|�|�����;���c���J���zV�tv�r'>O%fX-��߿�5k�0w�R�T3`�S�\E|��<�2�x��t��N�I.f�?o�F<f`�����?���L�,6�c'��Q��]��APYU�r��u������0=��ڗPDJY��	��ކysޑ]!��4�M��y���4^>�U+����8�R�RD-k�	����};�h�D�:�/ĥ����}����·�d���6ΥA�f,Y��߮孙�ya�$,ii�DވY0�� NS��:�v�jJć?!�K!g���5#ϫ _�G��vI1�Zm�q���m�Fב�������_�z}�L&ek�̩GT#tN�Z�ăAL�t4�����ӊE��R}��I�
z8��_�x��ׁ'_
��#g�kW)�/��
�uD���@@�����yT���Uor@Ɂuu�]v�M�6e�K�HNϠ��K�'�h������tǐa�ƨ.)P�(�x�Z4�[n���������c���:u����əLfvϟ�T1�d0�d�~�\V�qѸ7jҌ�W|GT�_0������|�j�� �\ߊ&������LMYw5��]]gN^M�6F�/iI���J�����DB���Oh�M��ޠS|��d�/*��&G�Д�����Z�sr���NqI)1����T�JI���HD��j7Æ�a�����s?K�8�Y�ؓ�A_^t��>z�ǌ��HS(@�]�Y%�l��Y��G���ٸ���������j
**J���Jk-{t1��ݼ��9r�k~�ǃ��Q��鯾����n�	��Kzf/����Ezf#{r0�����h%;5�wߙ΋�F��b%� �3���>5m�����6n�������=��+Gc!lv=N�����ۅ��
v��)��%3������g�~��̹�bZ�hC�'B�e\Xr�߇�b'��?}{��V����y�����$)6�����gK��Ͻyq�Df-���4n:�h�ம��K`ք�I�ѲY}��R��(%/'�d�T��>����;Yq�kE���W$mM��닊����1&eR$!2{*���v{
e��'&S�l�,Y��(9wr���тIU����nY�጗������~����'�����?vn�@�>~OA�W.��Sv��C]yj�0
R�hT*//�ez��[�Q���b���I��L�2EA�Rpz?6�2o�����с/�b!��	V��p�X�>ޏ_��mV�6i��-?)�+���|'.]NL��T�JS�����&������i�F2R�k���#�z�zJk���Fv�F=<x�=^:��K�վ:5#�K�.)��֭[s��u w��3��H��
�DB�[�TMT�B�D;�V�lN3�Y� j� MSQ��8JL�����Kr΅Y/��z9j��r�k�y��P@5R"��f�a�_���1l���ik�ubA7o�{��߅ޒLfV��¾�e�p����z���\�n@�@�ʯ0c��t&�8����L�a$����II
�֩�fQ�M��u�y�ow�����RּW	��<��T@n�V�:x���Ӥu�:3�{v#;=�^��/qC�fW��xhٲ%W**��$X�n+��O@Cff�"F~%74�ǿ��`i!]��s������������Lxc&GO]"3`M�%�O��(�&�Q�AЮy���g��))*#\^CVJ2�嗔2�jI�^�&��1��W0��(�FcA/��ϥt�ե�l޴�AO�d�Ѿ�u\ߺ�j�T�O\�P����� ^>o@5ξ`�ŋ3o�{Ly�MjB�I\���rr��(_�Un�U\��n�b���ND!Q�F�������{:|4��G�ᣮ�_��	�������ą�R��)n��S(̿��]�Е�ڿ{?����g�`��]����N���|�`��JX�EW���0V���o{c�iDe0NXgEk�)HZO������H���ts+�mF�nT?�����{���s�<��f��	L}s:i�j
��H�^�9��^��҉��Kqa�Tv��E̘3�Q�&a��,�c�[��<�]�yㆤ���DI���C
>����ҕ+�p�͔��au&)�lir�xٌV�K(��(:U�c�p�cXZZ���m�2��vq���Z}�N�|���.�s�/���Ap2���*��<�r���{̋/�g�6��+n_�ف�`!$��	�.J�d-oO����P�to�6���Ñ}�E¬ݴ��CG0��9�e�b���
��ý�0~���e������+��mԨQ*=�w���sU�1����MY0�
.�z�{�1=�/O~�7g-���AN��q�C��aFW.�Ep3�����Ճ�l$-7�%˖Ѭ͍T"�=~��>�9U���<0�a�%p�!\V��UA^����e��-�?yB5B#ƿ£�%�^S�I��a'�7ӈB!�Q� ޢ�DB~R4$=-�`iM��Hy�7�kNYyU^7Z���������PG���_]J�_��72���}�|}s�3N�8Iχz(v��l���+��xB���v���=]����+���ULz�N\($n�әH�Ȑ�Z��*J<b��������4*9f4&���dl�[l����w~<�Ց�t�u�L�6���'�͹�Y��:	�R���KKԄ��k��]FU�x]��򹫅^>/EG��W?'r�hB��h��`�%��ۘ
_� &�z�"�u���W]:K�]�]ap��)+:K�[o���7�{��U��5�7q���,\�)C�A-����+9|�~}{�����N��u�\.5l��'hд%��l���j<�?�,����n�ޣ~�@�m��đÇC�I�F�	8H    IDAT�N��:���j����N����7!:�eB���I&�$�J;{�.WF��V�o0q��1��.V�Y��ɱ���&"� ��Y4!a��O>��Od��M�ڽ8LY��#��ቁOs�rz��٪v��Љ[X��C�ۖ���֠�k))-��+�ۻ,ZH�N����e�;Hɬ�3٦u>�=���|]ɻ����1i�K4����׆���������b<;�)6�R�^����
���)xt&e!��І���A\E��ph?�<؍F�5!��K�����{���AR&,D�QV+q}H��Y�x�}�\8�Ô`�/k��th�a��?n��[3��L�ŔT��>	<ABx���*&�����kf��)�+]�ں����f��M�;���|���h�N,�T���k<�*�q5x��X��;�>;D,��խ+F���/a0�(-)�i�&
b�]Y�0����^Z�h���
��/O��$��b�CH����ʈ�������f!f�(�f����C��a̎$Q߿Nq]>������QW�/�ڄ^n�i�>��d�bֲn�L>z�M�.ֲ�C1e�q�,��q+�S&[岦��F��(ӫ�2�����"�3�w�b���5؈���*�B��i1��RLa�x��3^'��g�{�%j4�\�F�MEE5>_�^�� ?�
�wZ/�*���ߣ�����*��Pr����7ȿp�*q^�[ɨ߄�W�R����ᑞ�����4q��%Ξ>M�f�X��J2��QZQ�՞DeM-�\&�Zc�ZG8�#�"����Dsl�XTQ�H�@Ч�&iH�?z�������f�2n�h�S�#�����iX-��{Oy�ҪF���=%��۶���)�R����uFz�A1��>c�<�ͭ[Һek���{�<�G�s�!6n��'�c��Wy���4��F5���5�~n�7b����rs[�zm
C��xo�=�#F��w�4�ue��+��}�oę��2�-[���[Oł���g���i:ҲK?�RSZ�Ӧ��s`������B�[3f�X�ӟ#�Y����Z���߈]�$�E���1�Sx�&J�^���wU����8p���������)D�)0�A�M(U�]�u�d-��T<�/�g/d�;�����'�������G9GZ���tf��1��n��O?�eʤɜ:��6�X-�%���V*��j}�M"Y��7Uj�4�>����t�,YJ��}	h�$��b4ەIRyeI��+�Ù���hAc2�HTk�ւ�lQѺ�p����r��]�Κ4��:p�]����#p��ׁ[�������ϥ��S�·_U;t)��X�K�L�Rȯ��%P�U_w���?���jQ�����qv�;�+�P����LPcT)�tڭD}n-�������ؽ������������4��^�J�����־#~��w5�l���#*�2|��s6h@���)6��ɓ9w����<��şb0�p�|��.����p��A>[�s��ɓ'�5k��yjw�י��xqڜ�R#���j�`b��P��������F�z3&���x��,�C~����vl�y+i��*�M�˗/QVZ��b ����A{v0n��S�/���e�������/,U+�S'�*�xI<��!��y1�A�>�f����冶*o��;;�v�X,v��^�d!�>9��w?�M������]U���c(�|�[nlK��|Z�hFiI����R&�ɯ�ذ��WTa�x�;���N�0{��宻��a�O5���CcK"l�Mh(:y�S�b!rS��b_|�!�����
�k�iԊM��˕[��RԤ��"8������TԨf/=/��I8I0�!�R�nU� ��[48���A0�ѠG}�K���pЃ�nV�sM�e��_Ū�?�y��̞1�-����e��=9{KJ���HY�e�,:t	/��O�,��g����`��U'��*�HB�Ĵ)*ϓ�0��!�i ���Μ5�3����*E�(�J��B��Y,Ne�d����AkQ�B\/�A���!U��w���;���C�g�5Ƚ?���{����6x�~~\<���(�{Tda��E����:e\ݕ_5������QX�f���*4�Z�$4������-� f�ډ�X�8z���ط_~� �&F��<~\��CCeY1^��3gO��0O�{~������ҢJ�5m�o���v�kXM�6-�t异3�a<I<�a^}~�u;�F�f�s��j�w��X��|�=�u��
(������T:��3�����P����KN��F4V��8ĉ]���[��`BӐ����b����&Fii)��׬�Jq&���C�mf�oӒ�o�AFz�j��_��Wߜ��զ�t�B1�p\�K:�N��e<�_�&�Q׵h@�zل�^v��IF�Z�j��_W��ojI0�LA%[
	��X8��l��LΞ<ũ�O���[Tðsϟ4n�D����{7)��{�twu��g�II�ADAQ���Y׸~֜�,F@\ATL�� Q� "*Y����9Uw�<�����ݿ`��g����ꮷj�{��s�8��h	]s:�D���!�?n݆�����=�c���8| F=��68x���x����8�0�q�}fo��%�V�3�1Z�e��R&���͖,�j^��H�X��:�vxKJ�&��pB���*V�J�!fq#�Rf�dh5*�#�X�q�a�|N���`�'ЫS;�6�j8�L̜�$N�s�y�]�8�;����p	���DaL�Q��ѐ��d����b��_����P�Qt8�PS[%U�7'�`��2�9p𹘿�+#�� a�����T�-��H:��E�@3O"�C�U��,b˚V���#ݚMaܥC���C���Л�^�R�7�����o_�t�o�{]��K�ro�l`��,��2�;��T5-D7�۫�M�|M>�4����YX�t��X��CB~ܾaՎ�)G,1#i����L6!��P}9�Nz	����
�6�+�|�8Tz k֭F8��{0~��عs��o�v�{�^Q.#���ҥ�ڵ��t���kR�U�(�U�^�[��w,^�5��蓸��;E���y���ޥ��āC�����&׻wol޴V$W��\.��^
��&0D,�V���X3�Ӛ�����A`jꓓ�JFq��a���,�~~;R�	�P���`V3Ǝ�RF�"�:��ݾ���kϤ���l�ɬ�d��z(^&
�S�0��,� �$Ie��rf����	���܅p������EAM�	�f�HB1Y�p��]*���bDc�Q���"�x1d3	�T�K�j��_%h�f#��x�K��HI�@BW~Ik�h�cP4�4}eR�u�U��5Ҹp[l��n�M�L���8j����儧�I�3�z*���I$�h���^���=�^JVE��	�{��ͅ!��>��g��䖭[��#G���(~��Uoqb"dBce�������j�����<�����f��:c�uc��va��_c���r�WT���g�������K�dI�dD�1�lH�p�h�jb����$�m�����4RH��{�nvH�bO��ڑ�gMz��ۚ���r�-�{��{���=��p1��ｍ�ߏ�T�=N����t� ����n"�i�3�r�� �\��L��̶�,E0� c�G4c�#��$�>�0U�8��#�@�	�	x3V,^��m\���9P~���
\u�U�={F��իW� �Mt����ܹ��?��cGPU[���*th�
o��_}���y7��vLzk2�(~ܲ��
Pv䠌��سW<�����nC4�^��j0*�!8�4Ơ�mV�߬8	y��Ng7�1(��/��2`���9�/�Y�=WD��Ր���J�	����G��ӧ���PQ���[�D6���h�D�j(ٔtZǊ�M�(��T	����b6�@N1�ߤLf�#���&���78���DF��#��F�T:��,P,��aȘ4��tB�ߩ�@�L*Ҳ�[�$c�&�h���9}Q�� ނbd�	�q��X���#�hD���B<�M��e`HdD�'�n5	��i�#���ӶB���C�܆J�*�yPԦ�դ��Ռ�*x���W~�Y���x��.Uo�#�CB�#�s;!��Lv�UT��rBqؐ�zƤ���ٝYT��1��[R� �ꆻn�7��V��9���sϣo�A���e��#Oc͆-���a���,��Y�ɌblV$�Id�u`"������ב����Q1�����@��{�_w�@��w�o�ro����_�l�o���!,��&�zG��!�d6I@ߵs�T����!3@rTL����V�k�kB�C�5���u��U3��<�26(�<��L�z�����0����o�.X�ͧ�����-�ܹsO�ݿ?�;�A��W_-BuM�/_)sÆ�(.,�*x��E�������e�_�������sp����)�
�����yF'���Wy�o��I�ܭ[7��m+�IMv�aXlNC��Uz���Ui�b�@�o��J=��i���g��-p*�ڡf�����w�CYM�[����n��Уk�9�u����]��OT ��->mڵEy8����A8��9G�����*<[:�eaRi/k@�i�� KS����kxN+'�,�JJ$�3�&Cp*��ّ��Ӻ��.�td��~r|�UU��D�b)�3�p�ߘV��	�ΘUaS8�h���;�'�)�|y��ZOi������T��3Y
.ŎL*	�����
��E��'y�:��z$��)�����f�����Q\��pv�"Hi�ba��j������2�8�5p��p��}�n@�1(����Kz�! 5��0
G7��`0+��fеC<��=��%�A,^8L��e+V��y�KFն���܆�)�ؠ�]p��d��y��#�ȩ��9>���t�)%�L#�AL���_���4�=����
�@�������o��z��e�h_��V����j�g&lv~��Ȕ^�F�11*�q܆�X1>ib{�""�B�����u?��>����u�#cu �1�HUCNc���kT�g7b�E��U������	մn��&��� �8�V�¶_vয়YIG���E�ؾ-<�}�v�[v�={t�Uc��/[Ƅ�o�]�>��|0K��6�C��|�ݵ�'����1	�E�سg
�
�󼦦&z��pe4"�	��`FX��m?���	C6-?4F�� 	�~�T�LF��A<��k8R���Jg.5��^L��n��V	���}�[n������sυ�n���"��i���"�7��bҠmt�e��V�HHԢ��f��j�#���5D1�6�����*8�~�
����F�`��aG���2:h�i�ݺ��&kjE"�Yь|���Ȣ��	���V��;t�"�g�yrQ��5��q��x�ʦ����������i���D<�d85�K���=����3��`=�t���M�`��M������&�Fu��K�ӊ�Vm`J��hR<��Ƃ\Y�L(�pc@Z�m[��Z�6�+��eb�,<9>4pج���qZ$i�8n���P������|���>Z�n���VX��\q��x�9��0���p+���᭼���H&���9+�,�.�N'/E��rv'2�􉣇���?om	��`Oo!�5���ԩ���R���P�=y/6-]�[w����f��aŦ�?4�Ci��R͋�8�tyK~�!rcuu�l��X�a6��p�B��d=D�p�n�	G�Ò��φ��F^��p �W-C�v�DXf��a�!(;Q�/.Ɩm��Dy�H�N�6��j"�ێ���0��ѳg9v�_8
#F_����H0��7p����mmղ%ؿ�ؖ���	��J�hw:����ѽg/��b	��
�-�������#//�S���A�ng���	����׍��s>ȝ�{D#���Q��Y���m��}8xX���>X�
�i���A�R�� �50�qn��e���;�lƀ�t#̬�Ʌ6�Eq��ʏZ���_���,�o���
��*3�4����ĉCȦb04���2;�����Җ�M��X
�A8cN[\Ή[-�X�����	�J%tw�n�X�FbQy=���\t
��Y����3���Edޝ$BV��wQlvt��PT�`�d��"�P��(L�6-V������A�ϋ�ʒI�p�ʞF$#q����eQ�v����O�l3���
��e`s8���Ĵ���łPc=���	��z��!~۷[�.]O�?�"�t�3�FUC'j됆i��,��&8�.�^��}d6�o3�I���Љ<�8^���$���",3q��I/=|ǣ�x�k���R�7�[��7;ʗq�j������8��h���i��77?�yqk��|F55V�J�>�͟sL���?�0�9>a�^:�4&�F��$�dB`7e��?C��p5>�1�'��IE'�FY�a�w�P�Lvl��J�Ua�{3�ڌ���v��Q8� 清ݧOo�ao�w�3����x葧U-8x�\�k����+A�%�}zg!�Q ����}�@�_H�c_���۟I���5���l����m/��2�Cg�w��8��~H$� �"�������p#^���Ci��fM��!.@�6Ep�������:׻�Y(=R�P$,ۚ_�������D��
q!��(/V�Y�j�0I5΀N�@5d�1d�����#�ϟJ#�!"�u	,��Nu�ǡdcb�ѯgO;|��Y|��u���d�v�M1��HI�G�oG���x<B�N�P\T�-[~��{�	��H4��alذA֬sǎ5�BTVVbɷ�`��`�1|�j����v�BU����>/v���d�V���h�J%|�t��H��1���s;j���Q/ߗ��n����_��l�����'1�/����ǋ�� |���ظ~�8���{&n��N,X� ��o D��}����P���K���*?��_�h�[���֭KPUU��'�K�x�W�����\px���f�kc�[��a19�&��H��<�%�F�o�,�&Al5���BX��4	��p�y�^{�EX�l���[z3��OM�t鷻�����ݜ�����h��#樌*f![~�*���bo�r�x|'�N�ӡXڃ2�=����}�h�q帉�	g�4:�:�X=�:�
��z�#�iD�ǌ�_��C�q�U�aȤ����ƍ�e6w��Q�]0�<Bd�y���Ubڛ�bղE�p���{��U�Va�[q���y����P�Ђ_&���y��^}�Y�<	�+�[���}�.�uCMm��ۻ��S�T�i���'U�E�3]\�}��&������/@0ĞzN�"��w݋��:���B��H�>=0�oĂ��W;]v������0Y̢ڶd�f�[u�v%A��J:	^b#k҂���D����S�)@��S>6���-*��}�t!�sh �I1��d��F6Q�;o�͂3:w�;o����r\z�e�hӮ#JK˰z�j�޹=�x�>��q�>|0srs��a�X��AAvy�Q��;K$ѭ{���"��nD�~g���
��/�/�w�ʫ�b��i��?�������ħ��� ���I�a��7b��h�`�|n�O4�W/�m۶�9��B�j��}�D$�vm���G��M�ϧǐ�C�˖�����ǳ>��^�w��~��7�ɿ���ɃE�|�k�]�7�x#/�׍��B�Z�j�g�zƌ	O>�8���
�\y��Ӹt�hL{�L<���?�SD��r��x%ePNh�7��mf72���7dA�#�B�`��i�� +��&A��"K�BI�tX�֮�x�{o<~w)���-�{3�ȯO�~ٜ�{�%Kh����w>E��m-�&��瓀N�5+Ɯ����[�n+A��K�VO:��L%��x�q�|�m���E���8�� �a�B:k��Mä���5 �P�Vnxm�=�H�    IDAT���!��i,�v9~����QfۏT�!����,�ِ��~g�٧��-n~�m\��gc��C�ڼ����l2K��w�p����)�Y5r����Q���{
#/�T*tYB�o��r�Q��d��x�sM8�׫ϙ��U�"�Re/}�c�`�
���(�v���G�����
��Ϳ���۷G2���=��ҵ+^x���7�"���B�A��a2PD�(]��c$8s��Lt�r;��n���SF#|��H�x�5!��>Q���ө��r�#UX��<��m(����ߏ5k�Ⱨ�����B������<p�]x��[E���:\y�58�O/t�������_/���F���{�������C=$B>_���9��������������`̘1�-��޽{���O�6�}�ރ@]�@�w�s7^x�|�t)�>�N�:ʚ�ڱ�[�����E�xӍb�tɷ0e32��|�J���$|��l����H5UU��;E���;�����e�]��}�b��������k?|��r_0q����}�=��~�+��B�.]��'�qƌx�71v��%�ع�#.���6p� O�h�.{cF�:^G�����i2���D�c
����=����4�yоؚ����u#O��Ռ��f�-z3��{��K�z|)Il+?|s�����I�!���(��m�+tJ�rf���EE%�ۘ�,�����1�N�~�G+k��ˇ��5⪂x��B�T2����L�����nL"�Ƣ/�``����8g��g�GiY�׊�u�?���;��6z4P��'��3O>���rڏ?l��^�u�ݹ�������t2�d,�d�cF]��S�t�r�F6b���ܥ�$+<GZ�R!Nw�� aw����سs�T��zg��C��B �ۚMQ��ܽGo|��b�F9Sf��h���oa���9,� O���1 ��Fc0$��WN���ӑ6ؐ���٨�~��K&�Y	���өꀛH�c"�C��T2	M\rr�1[œ���i5O��̈Ǔ���x�,]�ل�EE���$̜=_���֣ϙH$�]��b����3O��k/E4�?���c�C��]1s�����w�)��o��@�{��{���M���O[%yRL&L�23f~�w�N���_�D(���:~��;�/�PZ*Jր����ߞ�>����v�D�.]������ǟ`����Q\\��/�cǏ�c�v�UW���ɘ<m*ޛ���ф�K�����'N�?z G���5v�X�~zWq���N۶mqN�r��;~��s�=׏��[6��o
�_RR��o������c���O=�h<�/}���RP�U�:��̈���'� �"]y�Ŧ�ߢ&�0��K$�͉��kN2b��>��L�h��d������>���-z3��o̘1����	�,��~UG�a5[Pﯗ*���Z{�Hc�Q\�JS�k��˨��*"mW��~�F��=@#�Pm�:|�{V2��%�S�b@:�@2� AC�^l\���8�بΞ�	�m��k�8�`������p8�@]%�z�q�x�}fQQ�L-�O����է���Z�}*�g{b@�m�8�=
���"�����m"��M�C��h�%2~Ơ�D��j�JI1�=�$�3��B���XgD8�����Ed_y����TT�	����ǰf�:�ti�
�N��O?}��̚�9��^��-�Un������T��*	�|tѐ�8D��l�hK
�}7��p�QSS�ݎ���ڽ]�w��j����Х]'����pyܰY=8Vv ˿�W_6/<�$6�Y��a������q��kp��_|1�V|�A����/<���:,_�_|�@��'�|��
j��OJ�p�"��\�S�.J��۶m۶m۶m۶m������m��s��g"&�n�22����V&�粹T�����n�ȥ[�}#Wm֍O(��3�`DC��n3
&�����eq����T�~x�S>���o�*į��`��3�v�ݑݼ�@��Z���p�h&���RjY ���v�HA �H��h7����s�����3)�h����h�������e~��������Tϝ�ޛ��w+�!�l^�V A����E\�Ñg����cx>��_7�d*4�����-n]�Xu������sa{z�T��Q��NH� ����4|�
�k��h�b��^��PUߗY�/uu���a�B x������T���o����}O����9q�O�*a��H�Jj�:����	~��6�|�>��R#�[h�۶)�-/�����Z*6m3�v���m&�ģ�Dov�k̤��@Y�8��Ⱥ�R�)��%T�o8��jqԤU.j0@�ɨO�2n�����5��¥h"���zԞCn8&2F������vT���K�n�&��F�$�9r$er�D�2�A���h���,�9��s,)(}��"�8�g�oy(���q6�G~_i�Ԩ�yP��v;�RȎe�y���kÓ	ý&�RX�߭��	��b���b�+���F�|٣l'(ہ��o�ۥ��azI�ZEҐ8�a̌���#��rU&�(	����xσ�
�����	�>2 �ҟ� Q]1�|A����1d�O��ʮ�R+��c��3������4�-[��n��{JXt0��[��x=��$z�!A>�iK�hv����Y11�0R���F=���»"-�l2���ǐ%������|y��>�V��&|T�T���e(���D<q��Х{ɑ��7����w�c伱H�`���N�r��@@)�>OA$0����RQUG��Ī��~� y$U�4��"�h�t�.&�1[���r��r����,��%���&YE(����4r�(]<�\�.D\�7�ԉ��S�;4��?B��Rrfh��qdFz�S���?Y��3t~T ���'�v:�:��?']�����&���u���~�,��f���7���̦��)�{�I����󼚇�����̮��׼�cQ�l�������DMCE�����ٳ�6:a������aGB��*�!�MjOy��-�Ù��K0��HIp�8� �A"f��3��ɖ��!��aVwƓ�FLEjF�����Yd(���Qeu5zS� +�ZS�!T
Tt_�,be��q#�bh�b��t�.&41B��(0L�#��,�>���_wk?ܮh�2��OD�	S3Se޼q������S�FN������Lvu�/x��@�� ����0�.�G��l?�`���d�)(_t3��B��ES�g#��Ř��YG�@��f�"���tE$��z�u��E���z�1za����!sF�#����K�C/�(���;���W�s)y����{=�\s�'�N���?3�s�NrU�6���5�Q��}�d������	��q�j��o߽D!b��'8���g���]^b8>�lg�W�M0x�����FRL�T��}=���p�M��T�r١d!��1^t��m�w?�T/#�X*0��og�
N�u����5���z���^ȎǷ������_ݎp�}��k�z1�y[G-^�gE#�'�
�n�I���V�i�zD�cFb��!c7�S��b$΀EZ�:�'�s?¨�����S������
�����K��|)X���V)��X5HV�xt�����Nqw�W��&�Wɋ�_����Ϟ[FK=.����`��R��D���r�� a?:���`���]]<O7��j���!2�\��zǔ
SL�6�D$@�^8r�����2��mI�Y�r�����2ǌ�QM�Y�Y7EJB�ɐ5�K��Ы'�˝��J��9��ǫ�����@K=O��t��VOd��}�"^DҎ;�j���K�`�J�
3VCZT}�7b���p�j����J���|����]j�h��+Enw�T����\h���	
�e��dD�G�>���"
��	[�~;.�b ��$����a,e�d�R�i�|V�p�C@P�'�h�� F�B/�{���e$��φ+z�4�4:ʄa,�E��裱���逖sB��	'�{˛�W_�L#'x��9�ؤ�x<:c,|*�9�S;�贀b=�.����6ˢ�w�S�]v�ml*��V�G-���n�F�v0A�;T��=B�{Q7���v=�O��
��Z�y���y�
y�����+��}��h���t������A������Ku{��y��Ͷ�g�`�s;!g�J@#a'�&�n4/` )�o�j$�M���Y�q��Q�^���2R��c�󻵾�}����w�0�9����y/��J���e���RO�0�8�L�ub#�y�-E|�8a�� ��p��-5T.���>�R�b���c?��`���>1/���drOwR3�\��PZ&YΖ��i�T�x�����	zݝ:R��������Mb��ɵ	�r�u|�Q�ߏekEW��\ı糿����|���������0K�\�*,޸!rJ>�Ė5A�C�rv��������̚BS� .lw�}eeU�Z��Gl�58E��>�q�?�X����ES-¶R�')a�l�Dyq�W4��y��v����[�����6 �!�o;^{��	�d���?~�5�)NH�9�dТ�o=r��E�я���?���x��Rٿ]�"��Q�>��{x��Ǌ��@�A<t�b;��DA؍j�c�X5E5�]w\>���Zb]ae���|{_O��&�vZ3�K�0DO��L���v�\[9v�4�:Q�w%�ǥ�D���k�Y�a�=�C͌"K!nFN�-<v'�G�
O4񐺳@�����>�\�N����&�e>��(5%���I�'#Y��7�F�;�9�܅PQK�%�O;+u�	��Ys�Ꮺ@a�p�+*+K���5�	����7�J#��d�eHW#���*�j��C�2J��6��K�|n�����9ՃD��\��}�����8͙o܉�H4o#&vH�M������H�I��D��q��3���!�5q�2.~�-����:���ׁ̣[s,�kN:��Z��U2�!��d���ZVZ�T
��[�!
ڙ�zܱ��2�9l"��`B��LVO���}�d5�y�<�=מ�-v lq�c{�!��:9ٿ����`)6y��'oC2���J�n���f��^���)��s;�;)�*Y~��宁���� .*TmP^Eo���*�&4W���B-M�ڰ�W�!�������]��IK��B�!�R�� �I&)L������gz3!��$��9i�VjLIE-j�2�N�ڃ��ڶ�`�W��'i��H<��@��i�zߣ9��}��p����ZXzT�0)�1����V?��lU��g&�M�[5�V�7��"Bᰕ^���ӡ�u�����4~�M�i+�%$Y"�{Rx���T�_"�=�	sįM�������Z.�A�W�g���AS�a��S( w�\��\]M�;kY���j'.��͟tU:�oac?b�0t>%�1�J��\42�2:>쫭~�I����Em�'�������-n�82�8�PS+���Мx�O�49�F�\�r�#o|���g/�����5�w@�
�*
pSe�O�z�*��_M�L�9�<+�+z�ja#���\S�!�6�|e$�HV�D�ViJ+�v#�f<��J:�p�
7q)�Zsw�=";�bIUs���O	Ȳ����V��lB���o����y}�
f,M���AS�h��M�U_0`���e�7�ߏ�ɡr� �g���IMg�'tE�~YL�\&�q���K���*�U9�|w;����;��]�ֲ~�V�z`J�CE�ϑ61��Z"�%�ת`ϼ���)����H��r4�2����9����n�Q"d��A��w���tl����HJgj��#Q35c�Z#r٩�_�&#Nʿ+C��w�޸^��Q�4j[�
 �����?�{�b�'��Y�Ê�����5���0B����RE+3W3w2���|DosW;U5�!��c�P'�)�'�<��+�>R�%�P�+p�=1�]a�¥k��1���߾�'������<�懮iB�#Q��`}�D٬��>K1��@�DT/eO(���	�����x[!�bb��'8��۷��1��D��O����_��q���8��"~"q���1�`��ȖHe��o���5gh�|�o8�HѠ�g�*��o���؊J�a�y=����cu:PB]ۊ�� ����f��S�%���^ݵ�(sN|4;��eȈ
*.��F����ڴf!�D�$�6�O�:�6�P�H#��.$��<�����D5�e�$��̲lqZ�ԗ���$i#{g*�v[f�y#Y+`��`]����v!?;������#q�D��d]-==� ��Oܻ$_8�L�I�g�)LP/����ּ��=3.�JG�ۈ�S.M\x�<�94��Ѥ�܄EC~Bč�z&�bJg��be������J8����gt���z�>G�:?5���o�R
���p7��&�dUP[@�)��ՉiK �~�2D�tؼT�H�Ԫ�kj�MK�O&�,�b ��Z��B��𾧞!�&��ӫ�(+��rk-������`�K*9�ꔜ��,ʙ1,��k���F�T͌�OqY��|]�.�֓�US�r�[��N�ߢ�4eZz�qM�3��y����v�|\ޟ�mh������ŉ���ٌ6����]|�M�	��8v�B��HT5����h�]�=��I&����A��DR�8r�tZj�^$F�m���L�<~�Y�w�=DG7�D<y'ɡ��na�u��IrB���3Q�=�(��*2G���(ŕH$�h$�;OT?Zn�|B��%�VBV%GS��1�$�Z��ϫ&��@�M���R&�w�`]�']
g���<��-��֥��JeH*FɅ�HH'(�s����aɆiJL�� p#T�Rf=�B�-l��,����g�6�}b�b��'+q���'/X7/�視���o��?��G�V�E��qOu��B�!�L��B����A	(��$�OP��¤�q���͊��;���ѭ�8����9�r�3آÌ�D���~����	F�� ��	;�x� [�;Mo�{?l��B����+���V+�����C���
��XE��T�"���K���4������W��f4y�u�U��G��[��0�:�Ν&���o��&L�,���Y�G�n��:�g1������XGZ���{��:�C��X
`����S�s��S^w}�~�@��.�
V[AO�Z2w��q.�����(	���"k����^�M/^̀N��"���Tu���؛���ݪř��Ϭ:;��A�Y��O"@�n�$�d���CK4q<w�PW/N�/.񌙝��39��f�]T��1;����� �d����^�,�N�֊p1`�x�ʔK'e��<	��!������Q��Ȍ�u���V�-eԬ�ǐ9�n��)�kw`��UHm*�T��V�T�y��
��!5�_Zc����|'F&��]zjO�E����T1�8U��dc�%T��J�vLVKD�\��V�
է�=��_�}�%5%Ve�b���>~��$�BA������;^���ӡ ��ff�b%"������A�d�z�����&%,O1�����x�^��U��f�ߚ�7|�}��p�6TN���j���A�L����A���~�Jg�[�|�Ӫ~����r�~�<O�)�򢭭�<%y��И���7���\L�Zz��n�p`�m��g*���8��]R��g�t[LV1`�O*!���Ow¸�T�.�l�#�Da��7��7y�AC>և����S�����^�;8�;l�]k��E�l����O�^/�@
&�cne�ܯqY��^��kXw&���c���c�N�}��qp��2?U���F����C ^��L��:� C�l�B{n�Lꇚ��4�;0=������ސ�K���LUc��Q��p"0�C��zC�]A�c�=l���M�J&�ÐM	��@�."*��'�f�����t�}w����l��������ӣ�rV��Ҥ�_"��щ J�����Ճ�hi����R���C�mQ�� �Z�W�,�0���
��;�P$�����`�::$p�^�&<�2!E�´?��\N��c�ۚ�!�L
���L60N
\>	ӭ�K�&QAHݭ� �o"���4�3�VٶRJ�1m���ԝ��W���P$B0l�(��]O)�9�"#�d'#j=}s�7���El�ltZ��7<���_��F�!�f>F�l��? 	K�~&wvJC�ht?���nI�����������?v�֍`��䝵Y��>�@i�]�E7n*
v�j�!�p�*�#�����AN�'�t#� ��q�ڷB��w��,���|�;Uy��+l�	|�`�M�mJx�US�ˠ�$���.�k��Vy��Z��6��%�#c+��23s�IIex4fi�d�_<��%H�2�ΦF��j�e�خ�`������s��nC_���a�1YW[ߏ�G���8�F&��5���ty0��X�@�Yo9��>����LY���K��Ǌ�������ʾ(�t�2�岈�(���8/��nù�����m�-kk'��a���K;��1ML���G�q���ai{"SS0� �Y������3Hg���k�U1�_̮�҇A*��挡"���5Fm��5M��JLS��W��b"�"%1���:�C�M~�lY*M��+r��a���A
���%z�O�C�J�2ۛ���S([�
,Z�Y�HJ:A)���g�";.@A�}�X]�Wp:��޿���W��IŦ:�*U�+��qh���'@�ٱ6v���T��y��CE��-������[���� G�x��O���E���v֣�1�kd^!��#Gf��'��D0���B�M*4_y�6%ZDu�=lh��8i��j+��;.8o|�T�N�P�� Z���w�Z��}$�R�Z��:H/�Ƴa������o�̳�K`t�2�3��L*R���������y�=W5Z��*���`������bgP��:̓sM��<I��Lؠ�(�Iy	����j���*�zKZ��N����ݜI?�	}*>��R������.!�h"a��C��˓��K�߂�P����� �����i���h��/� q������=���Hy��5x�0�)#�ԓ8Enhܒ}�SU��\1"T�U�P��l�,̡�bjT�OT��V����o�yA
E4��I]��W�Tt�S��+�Ҫ�̤����6�(�e�:0-xH�:?��hA������A4�!�P����_tx��`��:{�K��Ed_D�	�M�w^��&G4%��QH6�)b��ğ7��:�lq6~ޢl�G����6��V�p�-iD1����2pMh43e&Z�F��5d!2d�]�"�/x�M�i�_�
����.���L�A 2{�q���3�W��b��a(#� ����=��K�S�\���lCE�z��0�����qo	�b~!t�|��%$8�-FU�R1�,\1|��'�ezK|/U祐>�xwV|��t=�.��n�KA�
K �����i�1ӓ;w��dP>噐VD�[�����d)����ҞH�T�eT���;s>/%N��Du4xa{�x��d���J(���C���ȗ?��L����(*���r���;θ���'=�'W�MM�q�����q�,�D�W�S[�g,z�����P
� ��f�!��+PI8°���AՄMC_0�� �*zO��X�#��s��Y��"&`Wn��Pz�&q��HHE��7��A*��+l�{��oaҮ��";�_~��x�;�EIQ�4�v��Oj�P�s�	cI`�Ͷ�SA�z� _rD�s:�Y���(�ZTeFj𷭎�[� ��je;)�l4$:d�^KU~�8�佡~���B���:0�8��"�/��T�U�2Bn���g�["�:�b(T���'U
7����hmZb:�w��Ѥ����qmP\�a<�����Z���u9�.��;4X-��螣��#����`cɑ�9����c��>�����5�?�6�<v��S���G���H�?X�=���>+e�ż���'�v�:���z�9�����vr�]9�R}��՚]�U;��K>۾h�gd�|��b��U�������S��ݜu�߾��8}	�'�~�����/��lI�ϻg�������F�VC��<�] t��ٺ^ �	�~�ȳT钸g����?XB[w�h���>�b�}ͧYdV�q$hV��買��1�>�Q5��1�Ph˂�����HƁsn�Q/LoΏg4��L6�n׫X`���0_{pw��g%��F�!��5xP��4J/Km/�RN�C.��WK�H�&*6�
ѮΘ�\y#�A�Q{�6�(S���6b�`��c�͒c(��G~i�c�`�:l̄5�!�Q���OJL��eQ�XFsE��-z(�Qc�iBSP*��儬�9�[w{����	��}�]�TJG���~c����|��������w%��!���G�׬�#F��+��oY���Nʁ��G���%�3�@�94��r�I�n�2C�l�^�d3{��{v�z+�`O��T-�#Y��ѳ�-D :�!1௹\�e����@�N|z��>֯�P�fT�n�-�l�jZ����e��h88У��pA��{��W�܄+����v?ܰu;�d��IO��'n����z��M�|P���1G�,uBe6�55Rj�C�-�Ɩ�����O�QRgC��5���^Pa���O�Ļ��t�E[l���+�	�-<IS������� �}��c�>��b~�&/%z�Ƞ$�N��ǎ��4�N����%{����n���"vfh�C�]���Ҿ⥇qg�;�p�Zϟ�3?������#�
�K�����	*�C{_iP�@��d�B+��@�y�)_7[�ʜ�!J�ǒ�$i�ZkRp%�F�S��_R�,�3��]�C���WH.g/��5II�҅i�)&�fȕz� 2�$5�(T�6b�;*��|UaƢ��������Ǘ{n��-ܢ��/w���1�,}s�Q0���� �� �v��&H�/ߚ͵�'��րqu�j�B�'ڂ�s�K��l��NX7揚B�>�L;*���a1��C�����}���u4{,p�鿥W���1��o�"��ì�;���_\e�/����!���`���vw�8�j���"���\��*�����Pg�Y8��lι�{b=����Nu��r�*�/�e�\�y�QӝPL���ɋ"sxB.�{��SNY�R�a�Bl���kՅ���H�s3�ꐲ�`�Թ��z�Ϸ��C�ބ�>Oޫ�N	C�9k�ਙR$t@~�7�����1 Q[Ծϛ��?����Y��%^��+�����n�GE��c�!��JТL����Wh�$8����G�FWK�k�qMg�x�$}7 QOQ�o����;_	�܏��6�x����'��6J[��vhmhaڥ(F���܀@Y_�NN����Z%v�����k������{+�p W��D����΁��e2k��RƁ�-`s�m	7m���(��w�
�~�6��9�% �)J�R�?��n^&v�cC&�`�T��[7[�<�Oƶ�I'��JwL�WG�a�wJf��/���u��
�$SU�*�A(��c��Y�E�k4�8�F���O�p�$#Ǜ2��p����� �w*L6�(���?������{��Tc��l��l6h�#áy�~�gB?:q��1F6J�	IEu�{	��ޗ��z�Y����'����[.J_�u���(U�\�WE����NfF/9"�ސ�4m�)�¹[�t���w���� �WZ�G��|kox�.%�*(A���` �꩛� oibo*��|�}KK���'�rqdy�_�uk<�蒔��w��tE�}z|������I�V�q���Ë�SL�/�l'��@��sg29Ռ��NQn�F��9i��f����!�ǃ�#��]��Ѷף��X�ѩ��qa�u
�g3��t�v9Q�K����c��O������G>��nE��#��&V�p!R�]�\vĳ�ru0c WLfD����g�C
��j�G�v�P��'����[�p��_�ЃӠ��$`@�>�T�lʻ���=\��.]0�������U�4a��\AV�{�
AE=�{��,>C^�cuM��w_�Դ:�Hv����3�5��۪����?����!�ş/ ��y�������f�����8Ȗ�m���~i�M��3�qjY192^�1�@����<G������}q�n�v�w�c#�q�/��ba!��@��9����O!����8��j:��������EA��g�.&V'v�x� ���*���󔫞j�v���$�'\�>"���;�&`�B��t��w��NO��mD�������q�A;�py�����^wbT퉾����YAc�MX�m����G�,�&2���3
{��z���,(���4;\��q9'4���	�ƛ��7(8�aY�+�셓�++T��&��)Z���+���U�� �~����#V�u~ɪ,��ޜY�{F�wB�G/9�J��4в�6� �r�U�@c�53��6{�o^lnC�,�35^��a��2�aw����`��R=��7q���r��d!#̯.�����H�vjW�М�d�0J�YD���zJ��׽��ݼ`�it����Wi���&�e��:�`bjr�8������}�`��kP����34`����q�Un�.a�ݏUD��?@pܱ��)?=H%��]�>}g��"#�d��٩�"kIR�b8? ����!2 �{��"I,XuY��R�Ĵ�@�7�����>��W��BH;���"g��xx�9ϰ�Z2���*P~�`"�g/	dxl�-�^�}<2�axM��]��J������ç��A���i����c�%����G����F������rY�Ѵ�ʱ���`M/0ZT-%5M�N�0TaL&_Hry��:E%��,��a.�9�"�����S���ս�����pJ^+�X�̘�� F�(}r-b����80i>�������_�@-Ӏo�Q�y� ʰP *2�/�dRC�eSIVR��35\��p���ڒ.�v���ww&]]}�-EbmD�9�?�|ȟ���C�9ZN�jl5��Y�Ò����bY
}������J8��������OAπ��*ׇ���h{�_�;_����؉���^�Q7�[n�</����;���`�L�t�0k����YО�����/ �����_?���� 2cO*~����A{��)��z�,`\i?
r�C�jСm,�����ɏ5��e�\hʫ�+ �m/EfG6اH�n�^�U>�M�![��}��"d�����}?,~W��܅l
A8/UBR�_��O�u(Pf��d����r�w�B���,�*�������c����h��`�r"�z��&�]��������2��0*B:�3��j��������5�̛�H-�QA�O�jwO.��?"e"�ڽ�%�Q+7yg�L��֡����'j)�5�I�����ZS�A�X�
�~6}�u?�'��m��u����}b�&�<�%���OY3���g���H����j��������HJ���h��ҷ����`B���b�K<����߿}{��"�_Ok
�3�;8��3��.k=��6vc?��.���Un�ܹ�֬�LH�3��E���Ӧ��;���z���6Gz�q�4v2z	��C�1�ð
�@aJZ�S�9��t��(��ܝ�_�����a�ˠB� T��p.]OUWM42D�eW�lF�Ծ�[����@���o���w�������@d��b���Ֆ,X�v%����9!9-.�^N��8��7\�z���=�|��S��~�ͱD��ϓT$c����;�B��:d�)qf#�g3u� 7�)���Pc��R}C�t
� �ne4��C���u���j_���� ���_:���Az�V�ozBOP꽨���U�U =ZS��I�t�k��u��������-��y���*��U�Q��7�1����h���}_WV�1�o�#���F��'<F�cm�a���ܓp����xL��VU#q������C-N r��Q>=�:������^q�xB�1D��

:�[Ϛ�W���	�`��V�12
l�,��,P��٩����X1�̲0~~dM*���.���t���~ada71
9�&h �;s�R9怃4�YCD���5 Mg�v��SH�=_���L(��� >�HM�k��Ĳ�`W������,�Kz�,^��*B�ǚ�3���b�cv�Φ�#F�Q�5�]t���AD�r)�ϥ���D� jǮ�����`3�A��Wx&�3��C�|��n�my{�m���0�[�Z�r�(sJI�(��F"����(H2:)��5�0�A��3e7z*��8���fRj`������c��{�Wf2>�M�'r�)�;~i���s�0��,J�=C��R�yj��Z�s�D�9yk_���k�J#�M�e����I��?~�X|f�ա|<�`t�Brb��%�� ���<Ѿ�6E��,	�42�@���ۜ�S�-~������a�\�]t���CR�<ƃ���ԎӺ��0w�1�7�݁?�*>�щ��8ذ&$��L�'N��9�{4Æf�����]g���YX#0���� s	���@PVΈ)���N�r	�����H�R���#f!P5�?�p1zLC�Ԅ��y2���x�Ər����ҩׯV�~����#e=v���*JgTH�.�TX�B:h�ii���>=aT�ݛV��Z:"k��q0w�I��DC��i���4V/�!�5�p�r�q|�[2�[U����ņ���x�x�Z��7�͝X����M��b�0%U|y�9qG6	mZOs�ԝ)ME���âE���@�r��6�Y��~��2�O��O����C��EM �x��w��ϒ�mP2�{��;�S�nf��Ե�"��X��~a�J}�W��ikznR6ԪVq��~}@	E��#��(��+���'� 'X�,��S���ݎ��x�����n~�]�X����>�ڛ;����B�c1�_��~���~?�B�5r��$��2y�G�ď�D��ӎ�)Y�a���UI�Q�K��2a�d���e܂���`y�wZSK�S��<U�7�P����R=y����z`4i������)]�u/�F�H`���G �{�Ƥg�����u�S�HI��˦Thy���j+P�L
[�Z6!P��!����;�[7p#��Y!�\���lmLG�\�Q�4��?�8b��Q�˯�@ꚏY*P�d���xW�t�d���:�Jew�F/��xQ����DRAAd��N�I�.j"*���w���Zg�}�z�!�R/����g�����yQ�:ݞ�p���:l(���w��x$�ND�N���CQ9-���p2 �J��H^Kݧ�N.%����.F#���F�sD"��P=�(:=k�R�; �f��>��-���P�|�Ӫ��w+y0�a���ߋ�u������tI_ ��j%����p&�"�E+��>>���&ˮ�B�fi�����dΧ�C]��!����t����c��]��c�6���FM2
J»D5�U�<o�:��j��4�o���{�����p�y�ңx7�mZ'���X�D�N"�Z�m܌�Δ5Mک�[��Z�)��j���0Z�7,��P�� �s�yn�s�~�Y���鄐�:05�\�բ�e��[7:� ���EC�2f
�<��G�'4�����E`��K��@�=�A��%k;۟c(4:24�-��S��<6����j�G'�mt˔Mh����c�ʔ�\h�fjCp��6���ߓ�|j���o���䀿,��O7m�כ�^�[_��cfe�V$��y���l�Z�ۥ�G9��k�S�Ш���ܪ�tC|��gķ��y:�|�u�h�������i��G�iȄQ^Ri�m�8��Y=����:9�V7u�{�{ɯ
�]�An~ �dX���]��T���ƥaKT�-w4�s�s7�M�Z�F�-"|^g s\z�d)[eH)������	�:��
jb����9H�lt��Ƶ�q��k�^�s|_mTz�A�.Y�B*/��0S��f�a���r���s�Xq�Uըz�|n�IJ����m�CIA�zCe.�]�l˷�e���r�>�>�P��3���A+'l���` �Wt�����IM�n��g���
�|���Ǿ⥒:�z,�D�(����-O+�9o��\��_��J���~��oet,~2� ���[��{	��8�&�	�Z�.L�8@[�Q��A�,Da�l 93�{�I%(�B̀�]�F����П��� �����!f���Mอ��I!L�+�9g����(�4�UPU��A̅j�:j�x����:h���_�pR+[*G�4��j�c�>�F����0gP����9H�<�.�9�
�]g��C����2�ndy�4n���	�V�3
&������9D�(��?1`q��#HGEa��lx������<����c�}���[�J���E6����m�z���|s����WB�	����&�O�L�TD�b^\g�~>��\��x<߁~=�<����k�clv<E��?¨7� ��`�2x�H��s�Q�j5bKZd�.c�w^Y�Nb��j5�\(b�<�sPf>��JK�_�����UF��г	�MS�9�����Ȃ=�DM�1S!������~�VF��s�y��� .$��+��M>�쵚��$!Vd�uz���V��c���Y�{o��xW�|���'[���w� ���:���3t�����L٩E0���"�=��'b�b�V�� ��d��ֶ�/�9�4�X{A�)"5|�2G%l���;jM��'��b_���^T*��T�?4�T.�tޱ�(�9D���8XJ2�R�AyW���Ū�K8��|��fS�w��Ԑ����)�bxw�]%��Efۗ�f���� �k������P-쁀�	b�М�p8l��N����v�8���-��}�j����}w�@+�
é�uH��qK������$p�Ԕ���ŷ#!���|��"g��N9\�V��c�`�T� @�?�+����~��l�p5���Y{�&ԯbf.�fm��c>�nE�F�%�h��,�"�1�Ce�t�HW���ap�.)��|�(G�FLF7�L�_��<�u[���v�:�h�ZB�q����˃<�}�Ι���O7P�z������0�)�	�_�do?��t���)�5U��[�7b,d�� U�f�8J��h�j�߭y�����Q�TC�i�)�����'�\�yb�<1�3k�h�?Tz3��E��s)��^�K�����R$^��@��;�������s]ɚ��&�\յe�$�|�i_�v!�g��ϗ��M�wL��ީ�p6N�rx���U)�)1_�)^}�"��1%�� �oS�p?t�����8/����VX�}�������J�:�������P���(��F�S���6���m�rٰ�1W�В(��;fcVVLQ���D� � e���k�k|سb�Z��0���Qz��B�>Jk��r"�.���Lǝ��#G�*X �&��[�g�/xf�o膅��9y�1i��|\4vYO7Zr���U�`2������᪖
F��e�33{�E��*}a{%0n=����M��	���L����u�\���C9	vtT�=�L�3��{�xV3��X`2!>��L�haÉ?�i!�}��tB%H������w��.�����z�Q��<t�թ�jO�c&ѯ���!un�����I��I���ct5^P��4X�e/<�]��P�A� ��*�@(���*$\]I�d����=F7�pmw�a���k�h��:z$�U9�F��Z�,���cs��w{���0�^r�*��bq��O�Fk���6~.�a�@[�A~�����e
!���5�����A�q�oc;v�aW�p����шip#�S�d���(!F#�h��T�^��2O��=�˝5a*�՜�����Y����g�a�d�uy�]�,�(Z/��MБ��!�
͛���]K7,�a�_)��Q�� �@k���ťxu�hL�:+W,5��S����Fl޲�ϕ�Y�8]X�������3�_5��.�P���/�!@����?���_No�!����#���,T�S��!!��2�@'Ee��!*JH��V�MY�B	����R'n���gKZ\3������B��������r��Y���Iuοӈ���1��N,�T��Ŏ��Ź"�������N�f��b���8q.N�.�Ӧ���=�p���3xt�������u��8y�4��\�Ą$��0�.[�>>���(tZ�8�-�
��n�-G�.�a����v�]���]놗_~����+*�+�2�4�n(1�~�lP���Q��JpWz���o���z��"�T��w�E�������t>��vF������F�>ZxplLe�� \#%�W��K��r�
x}N�c���ʸq�y�|��ǈ�&VM��&����Y⠋M���$�ez�MSG<�%%%�^nk�C��z�XPR���G79�.�/>�Ic�Q��C�D2�]l�X*}����A�sY�ʑ�ҷ.���t���ɹ�T���[�ݴ+�v��W��T��ˊY.��΀� �`��u�40���U��4��J����%[���1�/�r�</l�SS��_�`4#�e�������5���st���>�ݻ�ô��_���Bx�,_��<���*����r>g^����P7%��t=R�q��=(+���#�x�Idt":];n���~�mD[�l�D�O��r':M[D;�q��?��Ն���t�Oĩ�����QkA������z�}pSX��t*���)��x�mK1��˃+�[L�IV������Dqa^5ƏǮ[�h�,�7m�ׅo�Z�Z�aǑ�X�u�>�о��#��+���/�x���S���w,�v�����
����^���P��65%����W*�9@�'�Xdu*�������ʞ\��\��e�]
�Xn4�^�2Ō��^�������.+~sz^��\ ��k
�_ 3eb����3:���N�:�Ri�t8��w)��k��*� ����i:�
dB� ��7[�x�
'�9��N���_�Dlb"|n/\��gO#1.���?v		I���BNv4j��Zu�P��p{8r�_#��1<7�I�ҩj%Ǣ��"f�x	�Q8r�$�л�ۛ���/W�RR���"�Ȋh��z�����@�"G�2�G���!=��V�*]nD�3N�65:R�/�Xi����P~n�>���4�D����`�7��N��^/�L����*@�Q�o�|@���L6QW�9Y�5r8S��~��+��kZ�I�4t��.��n�.Yv�_�+A�i�'{�������J�=�O����'��_�5�r_�Ӊ�d[�9���� �'��1�A?uz1eJ��S��Y܂+0��.��pJ�]���(��_�����	�QI�+�Ye�ץ�%�/^_��=^�H��O:M�#প�Gz� 4�~'	�D�-=d�����v'�z9�U28����t*�vRgkаQ:���k��]�=~޺ǎA��)���^^�f͚����݉���������Y��w�M7wf_�Z#�yI��<�Qx�4����]�h��&�.���ȱ3���Mf@���k|-�T����Acw��p�u�b=��E��^	�Je,Ǣʤ8�*���t�sz���|j@k2���:�!�����t�
�i��xi�襀N����=�K��
���(���!�S� '�F��{S�a�/Y׵�]hsMk�m�	%E>�Ť�o�Đ/���S��]����x�nݺ%W��v��zB��o=��{��;,��$%���O��NY��ᑕU��؃C_d�\�I/Q;+�$	�eL,�^V�.���S��8�]E�*�p��`�Ub�����6G����w��%N�[� He�V��ų�-�a�UXٛ��5�\lp���qI "�V��k{# -V���rZ�j��'O��3�3��v$&&��(a=�4�\��6"Eee�X�a6@�/v[֯[��ݻa֬9�h��O��s#�G�F1t�P���`��8��{�J���G�r�~o��Ѱqz١��R�4a��:�u�����I�
��<��9��8u�d�CgA��'R��|o�j����Ru���i$�p+ha����u�܆�A=Q�uB����Pr �G@�
�^��J �#x���}F	�s�Ч�5	{�mg@���^��l�s���u��V�l?|���E�N�o��aҳ�=���}���W!@�o������2kV�%[�m**-�/x�y�I�Nd�;�����U��	�	(e�X�[��dUK�.����X9�E.dP����.f?�N���( )�j��N@J@K���j�EշZQ��&hw���*�E��r��$5��-����4�JS�V��>�dd���-77��hf/�w�R�B%..�3㋊K��y���[p��I��m'�~��v�G���^JI�)`u�í3#���)u��aZW��M��g�=���$�"a�e��;y�[$����݄��9�%p8����Pk��駟!�܎�u��#��
�����m5<��P��Ti��7@�s����M%*t�*��"�f����?2�������Bu}sd��0"�ݠ�PEɎ���S�(�z���U�WA�� :��$�垟��F��9s�e�z���X��F��b�ӖЅ�#�!c��l�6�!@�?����}��O��ߜ5����G7:�.ÜW����c�V2�=�r��	)`�$���xddd(�� p�B8a�"`�A,��N �]����r�xi���b2�����F�,{�t�8&�C�se�*'l�y������!t!˓hP���0���"̨��ƞq��Y9�-x!!�u�z::Od��ɹ\�111�*U��pyС�(��b����𣙸����|��D�}�����ANN��p�uͿ�=sW��oX��z2S-]�Sv��q�U�N�;������ѽp���D<��SШM��h���д9��Bm�
�Ȕ�N#��=��~�)bU�踨B'Ю�}3U_5���t���̺�ѿ/7�Q����_[��&�#�i�) 9�]\��iiʣ��Ae��E<7�,�;�lۈe���h�E+p�Mw��2Ae���Sg���1��
��q���OMM-�o�[B���:!@�k]����P��hӑɶF=������M�l0z�{�쩜jF�E����X4m�T�Q5�,؞��1�P��%�NB �}Z�fW�ryه'@w;�eN�a�Q�T�[�\(H����PƷ��T=Q�d�D*�wr��`�p_�E!9:������`��]��H��MR�J�����h�w��)�腸Πײ�-!!.Z� �}�6��QVV�����>C�v퐜����$��E�ԉ��v�=HNL��߬FA~<>_���\�g_�F�޽ѻ��X��f"5���_�v��I����l���x=�+-���Y\��D'���+a**ƣMZ!����*��)Ɏ�_!�}�zßt�
&�]�\@W|��L�����C�º����Y�A��⚧G������S��� ��𛊟\�ӸT�X(�c���Z��c@��D��Y��cسOa��Yطw;.���v-Q�v
�ed��[{"`����"�7���ڵ��~nܸq��Fzѿ��_���;8}��s������2��4^�$���a@�|طo���0��$%x˖-�[测���!*WY�J*U*�e6���d5�7d�Y����td�����&K�T�S��1��ɢ��C��"��}2rT�S˶��a��ztЍ�fw�n6$��R�G�,� ��޽{����A Z� ������=��~d�h���:t�}���>cM�����S����׷�*�Eaa>���~M�Ӏ-k�'���F���?l���c�/Ƚx��wb��`�i`Һ���א���{��Bv!z�ꇸ��_�1v�H@K��tv7{��0�E%MC]�W����Wtq�ʠ�� ���j_j �]�+��"�.�� ��s�M(�i� �J��G3�hj�R�S� t�܉~�jT��6 EP����s�"�{�f���[0g���qW�l���w��e�+`��
;�M����r�m�t�kC����~ϼR_!�W���{���f������5�|�i���0�-�S��p�]8z�([�DE,�kd�!z��k^��$�I���;�,Q�r��̂'�$�����{�s����V�A��!:�́)D��j�^Z���BLT{t�uK��Pn-�^�A�ŀبp�*�]^Xm.�Z�px�9S�Z����eC��#L�AJb��C�5�q:�n����4���TQ �·����.{�F��{�qq1H�[��	�˃��� �~؈�˗�[��������-�܂7&N��^��n��0m�س� r�p��i�3�}<;�9N�ۺu+�L�l��]���Of����G�h��qgg|�nΞ�A�^}��Xg�C�ݍ��-_X��r'"Ic@qȊ��v����A,�Q�~��M�p~^@���h�4R�N�Oº�ﹸV���{�6�`O�E����A�"�ưN��Q,/���S�L�+�vZhqBݕ�A�Z���Г���DyY1b�0|4����̟���w7��E�1��o9p�|��%V�h\o��
�?ps��6�UvA/w8�:gݞ5И��>�����p��e�ruj;v�2��o�~"#�дYse>:��E� m!F��6)$����6Υ��T!;]v�ѿ�b���Z�Iij�w��׵��=P±l��ɲ�f >2I)��5�/+Dv~.�j7nm߂G����"))k�ߊu?l���%q��x!PZZ���'�wW�e��Կ4~´?����|�r�h����tj5DE��~R��l1�p��ol/�Y�#P���HLN��d����Bz��[�طw?-Z��n���x���p�M��͉��F���e�Ͽĉӧ��U(�V`��ߠG��ӧ�����`Ѣ��ʺ�VBnqx�x����=8r�.��G��h�� �}��]�5E|��Z����z(���Ao@�H�C΅�>1��ǠzEe�vF�b��8�*��8ZJr�	F�����re�:M���8�2�����(T�}(�9���B�^=���#�M��+ѱ����vEG�T��*m��V�3p9��i�(����!�0�\l޲<�	QhӲrrJ���Yhͱ�E�̧B�K��[����4NQ�5�~�Cz����k�|�o�J

M�'���g������5ɲ���Ç���d��	�jݦ��q�,meģ���	e"�Dzשb�	�x���J���/"''�OU��i�Y��]?"JW�ݻ~�5�݃7&��w�|�&QF3�7o�
�Yy8u�|�b���ܐ����W�{����gp���І!��D�������3Ⱦpz�O|o��
����f�΂7�����F=���h�?�' �L{! -��~;���"^��F-Z5��D�qdAJKKǉS�p��)�Y��w��Q�f��`wT����A�V���Q��G���0`�`�]� y�X��w�ׯ�rrAʸ1�_�ƍ?�ȑ#HJJ���W↶�`�~ &)	��wR��弥ЕXqK��{}I�(p'�瑧����AQ(*�����>?�ڣ��ʿ�BכF�ċ��Q���D7A�k|�^���e��f�[��ՠAr�Fh�.Qw���+�=��m��񹺊nY*?���l����	�
(���3�<���NǮ_��E3��݆��oĖm��sy��EšԧAf���'�0�o���P���/w�Wѷ��^�?qؓ��o��ǃ[���M_�1C�h��Ơ�Z���D7V���AIl"����>���j���t:��s�[ο���8y�d�qz��Cpb��ϑdv�ӿ/�C�=�������?Cdd2zӌf(����S�K    IDAT)���u�`�o�}�X�h6ƍ�>_�Qc&��6�����-�p9��8p��^��e�ߧF?�4��t%Z���2��%��&�&�[dD4��#"-B��dm:t,�����$t���ۃƍ����_�#V,_���0#�&�i�4l�~n���ի�M��`��}��8̘=ޜ�6Ə��/��z�kq�|@��xs����K���_.]�ӁܒR���F�� 11+�/����u��[�Nк=t��:5�[��4�h�/2�iZ�e4m�b�l�l'Ti�q����|��;��/ 5U�n�+�ԈLN�9%q�ç��6��14@��%`��G��s^�����'Q)%�6�4"~W�#G��;�E���Kg�I��HIL@�VעC��a�#@/�p�؊��z�w#>зe(X�O���MB�~u^�K�jڒ�mg��x}�Cꁘ���tT��\�K1�t����h�T��/�\Z��0��.+8ie3^�=�ji���ٳ�DeSeH��Ť������������sx����y�i��KLAZZT�=�s{)�<�w�r�|�>>�|�/�*]4�~Zg^��pΞ=���C;n���{z��v5��5���R�3{>;�Uᑑ�H�O�+�p<C�N�Y�����h^��b�jw �n=X"b�e�6,^���vzrJ<ꤦ@�g����q����cMaزmΜ;����aȐ!������?���~��?o��snC�F�Q�uK>z����
�˯{���G��\K-��������aρ�б�<�*u/����j�X��t�PG+�?��)'�P��JPU�C�i6-m/>C��gC5��ˁ�$=����v+�\�c �ޯ���G� ���2W�u��Q����B����BAN6F�~&N��};�B�9 ��}5jKT**<Zh̑x�ű8�U����6�>|��m�4)����!^�� �|,�Y��y��ܢ����=":n�&����ٿ�S3�5�h� ���*�T��4E�27t�S���mI^u�YYY��Ϊ�I//+�����%3ct�ZQ�FM[a¤��պ_���Q1hԨ|Z-��8���"h�ě/��\��1�	����xq��К��������iŁ;x��m������������B���{Dŧ2xS�N4;�^G�Ah|�]ɘYY����Z���ի�Cn��� 19%e6�>}+��)n��6�z�[����P<Pitp��3��B�鴃����\��Æ��%��~�w����x�١�ر#&My�=���<,��6b#�p�l�o؈G���ZX�`1�j۶m1b�H~M�I��0<[^�h'�\Z���NX�}��*�U!�E���<�$�"@��^23��&ڝ��]��d u����3�i��TЋ��8��g%�~O	���E��M�9iȶ�r�(� �����?�ӕ�p�7#�v
4h���z���}�e��-F���~y��~�[4h�w���!��3�?q���Mޚ;��O6�RRPȀN=t���"&�V��>r�7���(‖��M�3�n�r'�]gL1�̬�e�:�(6/
B��B
�S�N�v�6{�=���PQ^��-3�a�Nl�uN�ɱ����8�>�<sY�9�8�q۵��,���:��M�Pa���k�rka��G�f|�,*�Ǒ�`ҫ���[;_�#�C�U���u�����RSSY�}���S�)d�T,�#ʝ ��L=��5j�ۑ���� �v*�z֮�?lڌ^=�g@/.�ELt�6'�a���'�&���cެ��Z		�3{6��V���Kpzh�GtlΝ;��	f#p�|v���>2Q��X�p1tzڴo�Q/��
���Q�.�޸J��n
y!�Uc$tc�b�����U��x�u�*�R���'m� p��)�x�����aћF͑�_�5*��*��J������眔��4jx�.���ee3�>i�$�:}3>x-�5F�V-p��Y���0ꥵF�݅B�m��w��t�{2C>��J\=�� �깖�{$Ћ�r���,d
�)ѱǎQDobĨZ�g�w㴦��6���&�\�S!2��,A��:P' ���z�ܥ�):�T⥥��x�p{��_;)�&�.ؽ>�V�p�|tZ�"���X��>wٹ�0�԰h�h� ��o�0'�.��h"���״ez��aߞ��j|0�HI�M�2�0����F`�����OOO��t�J��\��&[��G�aʝ�V����"�nj*W�T�RPMR��HN��U��G}w�}��QZ��zuk��v����h����6�]n�j���󚗗��^{���EJB�-a���O��s�qq/<�
�qg[ڿ�f}��~�X���(��Ѿ��3v�i\.�ʩ�&@w��q������z�!5�B�<Y
�yz0�+!?��)r�y��+���.��#��F�\w��_�q����U���&A"�Tp��ύ��\<��3�p�سw�}m �q1�W/�ݫ�@e�@Y�cѸ^�-o�t�F��s:�?wB������Q������<�p�s�b��ʊ*)�E��B���E�޴9��)^��T]S�*��5�t� �*Z^&�1�U+ �/��D�zaR��7��$9h��k�Ώ4[Ă!�AqiW3��N�
��^��������s���0��8����~�l0�TP�I�M3�]p��HLNe�[Y��� H�Z��j�)��ǎ�
]gXX8�IkԘ��6��鋨�D��<���k����FРN-�ujس7v�N�GN�D�N�p��<?r���PpX+�z�w�bc"ѣk���^4n� ����O>BqQ6�e�V���#6&|�ˍ��?�G �SD�kt�ۧ����5\>�ʘZmP,�^��<�-	ңT��4�O�Z�4O��|^/W�Ԃa!�V̲��:o$gpy}�җ�z�4�7�EA^�~�I�]0�lߌU+�a=��hpם���.}p�l���7&�o��
}݄g�?��k�Is�k����x^��kl�()5�z{��w?��P�(/.��b��c��LT�B��(���lkºE�!UsUq�r��Ӎ���T�����>=8-�G}Z-�CGU/E�B�N��)24��s�ˬ�<>N9ӫ=��'0� ���r��r�{���~�W�¨)��A*��8��7�Asu��U�SR�'Mf+..����ܹ��r"@=����u�v9`4����MH����Ɵv����bl޼O���}�&
��Y����jJ�|��[<��s()-��ؿ�\���������U+�����>0t()��?x���p![�lǓOCRb*��#��������"��u�&���Hl�^r�#%y0�r(����w�?����Ѣ18���e%�׫�@��a�������g�q��)�0�y|0�#�%��h:^����[�U��Ѫ*<�X�v:����MF��G<>�i��E5�:�˜��׀���e�Z�Y�mkan���/b��g�7Ep_�|�z��>���覯�`���l�=p��	E�F�(3�	�hik�Q�r"�w@�S�^nǀ�'Ϸ�Ru��j8���PI�!�yUz�=�J�8bj����4�z��aZ��x��N��=�~���XN�=��-ft�y���D8�Ѣ��z�ȑ�(,,�Ł�sp%_/��v�>��h���y�>8=>���}�zu�*�u��P��K����j�_Z�f��G��!+7��zu���Io��U+q[�1��G�ܰg8��Ա}X8w
�5���l޲�{�A�zi�j�;q�=�0p�@q���D��"K�˛�����HPS��⌀Z ��J$�>ZD�e�2�M�ٮ�
��g^�wu+�<�����9�
���~����ѣ0��w�o�N,]<}zuǶ-�1�������V}��;wc����h\w���_��k�=��1�5��O�?��ܵ���\��_���3��U�e�B��0�.��;X�ݮ}6�I�|�^u�޽.997\����=�b��|ue^zp�;����Р�H����F+I5�@��U���$pF�%�XJ�O�Ia0����2B���g�{��:�E��V	�Җ'�+1T��ޤz�=?ː�
z�'��ƍ��s��� :1	�j�D�X�1�?��6��7t��?
��Τwv�g/fa���0~�h��Z���c���P+9	o�6?�q�QHOO�9̈�'�Ι0h�8r��8����Fxx,.\�ۇ��vŀGא WK��}��@	p��@`�����'�p�$]d�Sz�T=�Ǯ�܃��j�V���T�K@��O-\$�^�Y��b�ˣ��;o����X��#4��������ɋ(,�#2�.r�lȳ:؇�:#�ǷFz(D�_���B��ϝ�+�&͟�j���[r/fE|����@W��Q��'�k ����"��VC�L��Ѽ���(�).t��2���栙��Eī��6�y��R���ʓ���"��Nzhb��*�v�jR���x?[	�0�ЋV1�Py��b`�n<�3O��U���T7����i�B�'�8�ݯ��b�����@�LF�k29A����e�К"P�p���1"�ϝ�w�|�'DZ��H�W�M�#�"99w�s/�8�/�Y���������E@qA1�~�-ޙ4	7v�~���GX�`P�pC�FȾp>��]���t���xQr����#��3���P���6"9m�q*�-�� ]}Y�z@� _êGe&�Tk��Զ�����:/��bλ���1~�8L|�<�+�C��0Q�"��K��Uka�J�9>v���D�7���q�{��⮖O�?~!@�����o������l��Ή$@�g�'�����'U�gϞa����j�*ӎ�ߨT�"�U��9ϛ�W�HT�WF��L��_.f���6ѯf�����Ŭs7!+7�����2��Gq�"|�hy'�Q�)�[R}O�)���d����)aᴽ\���Ѿ2S�Q���D�S�;�"��h8��a���M3##�	�e刊�������s�a����xIyV|�O��0#2�7�#}��w_������S�Ga��s7i:�Z��
�~��p¬ע� Z�=�܊���%������棴8��68�t�� 2Zeb��Sa���=w�����6��(���� ��T�UJs����,��~Y��j�`�� -�g*���	�/=+������E�R;J.�|n���0�W0�q��a̞1� &2
u�6A�n�PP���c�0}�|DԪ��������C!��w����p��m���B���Ղo�n,�ɍ�d�X�}v0,�qp�U���~�����d���*>�m�vj=��v41�T(��9VU��e�KG�O'ʝ�6@]t��^�n������$����"�������>/���h�$	�4h�:�=>aâ�2JP� p�����։�dh�*o���>g��G0	���*t�ߑՎz�#"T�@����� �j#�l6��/&��U`��0e�D�ׯ��sg0t�8��n\ߩ#&�7�������左"����԰���>s��?v��F�f��+�Y�	�Ǎ��r��sz�釔�X�tR��M�6x����i�,���I� 2��,x�����\R��Nys�[2���[�7�ʝ_-%��-����z]�
=O熆��{��&U�*���*��ƌ�
}��hެ2[�F F����X��g�ݺv�E�丵�����s��j���_W��a�-|�c���!@>�/���af΍Դ��e�
ٶ�~Vn�����p��vT-!�'�$�#Pg��Z�)�����i��4��/`��������Ʃ*�_�ԫ�r<%�tb������9�A�ۈ���SO4=U�t,��ۥL����X�N�X����������(�?U���Wiu0�l-��6��V�D�åRa��C�z|�d�@�׋�hԊ���/���ۃ�}����F�W��MP���0�lv�6��%���o�:8�J�u�!>Z�/>��O�����]{ѭGv0��n.f�_�Gпo�wyJ�1"�_iO�D���>���/�(@._�ދ��F�
pW��v�|�=�U��T�ә @w��Pܼ��ɺ�q��aʝ��?[�����u��踆0D%���SP����]�ѮM���F����O�շ]Я�k�?��%K��[�{S^vN,Q�/�q�ٝ�)*T��6��"A�MT���9�p�E����a$u�`��3�gU��]9��vHGh��R,��R�B@���8V��9��Do�Ga��nPT�^���&��T�$�Sq
������1�|�	��Z�;���N��+�zAߓ�^��Ĵ0z/��t:x[
�!q=G��r8��� ��"b�WZ��v@�bdI��#\��I�B$MqSD��ɵq�|6\*�p��0D��ꀁBߝX�p�I�<xd�Cօ���bD��)س��8���Fll2/Y���{��ʠN�tb%d�+�.��� ԫ�(dU/)z�liU������xSQ��\���V0�$���.���*r/^��1c0���r_�|��GFZ:r�������'rs�u�XU$�En�2���gd�ր�Z�/sB�^>��q��kݒ���|�XL�"-�L62�J�N��B��J��=rzN���sn��aMձ�!�JVZؤ��	b���ь/�Ԥ��z�^�<E��!�@��ڜ�:��+$�xߪ�|peĕ<U�$��*Y���$D�{<b�L���؅-ͧ���9��~�`7H{�7a	3��t��4z$Ԫ��_~���~z���ԹYO	�>^PoCg0B�7����A���(�2E��v�H�l���vC�*��Q�Ê�p-n����B���tyqw��[/_|�5g�w��}���>�׮��Dh��u�}U������CQ�_򸊫���dv����?s��@m$j}h�
��eCA~.F�z'N�ɓ��`��xY�^c�Y�3�^-̉�� �)j��e��'CY��A�������C�`����?�ZV^��q���0���:UM�B]�I{�d���g�דϱ]�Ke9��)9LI�`(A�~/U�@e?].&�M���J6�H��
�"���W�喂���Uv:�#'_:��\|�~��l6��������S: �th5���C��t�x�B��Ά�8|�y'�j-��>1�/V-��t��ѣa�i���F�ƾ����d|�� v�,@�W��Z���}�"��D���!O<�ʇ����x���9��wz�xѱ	X��L����v�ߧ7���#�~b�E���?�j�j�ߋ�t��}�^��">;�7��P��H����8{���|��pb���@���!<?�;�GNBmN@�ZɿL38������2�m��/����s���a�֊
k�'S_a@�"�CM�`I)�wp�-�q(Յ��%��6�zs	zR�.��I ��:	���'�c��rAQ��.+M�/��� �h�Inv�H���F����m��c��@2��Y���n<�Ä�_�7� �_�����p��۰����~Wg�A��4|��tN�3�Yp���p�B6�-^���g��(v�Y�s��+@�ޏU+f�N�($%D���<�Ϝki�+����u덄�ZX����w������W�T�?�Q������A��[ToU\���������'�5�p�+�'���ñd�Bl��=���d6C�V-q����S4�g�b̤��X�D����S_�33==�^��!��_k�g`���Mg���¢�h��_{�iD�E��
�Ka[��[q�l+�ru�vY�K�La�^���It&�����!+wzMY��}�
	��g�}P��7�j�2D�PSv��b#�������(:��y��H� �*tJ����S��Dxt�#~�q *���?]����	�z    IDATj�G!�V-�6�UL�4	���*�v�bL�`&�}�G������p�����aj,[��-@Rble�x���Ѧu3�۰��o��Ï#6>6l�No�M7ߎ��B��Dl!@�׿���=�?t�~����a@��d��6l>z�}�9{3?���-��[oA�Z�а�58u� ��b����<���2c��^�u� �_��W�+�*�+��c;M���M�~**.�]��X�2tW��Cgz\	��WD����e�|GY�K��F`��k���T8����e����hYM�6�3.A�: �6ȃ�^����N��˛�|=*J9� �o��'!�7:�<n����++�`�B�U��	�$��^�����Dx�Fl�w���ZZ��fa��G`1 ���ѼE3�۷=�0ޘ<�r�f�F�:�#�9W/��I�`�1�[TN�h����<���l�ٹ%�'ѪEdgb��?�O�Gп��[��,���~1HGz���/Z#�H��'��n�{�O>�ϐ��J��c�k�!���)wr\8{#F���?��=ۙro׾%����V�щuq���~���hڨ��w�?ӫujjVͽ"5��C�^�?U���R^Q�t�h�4�1t1��πN�(]���s�ֳ�)[R���+Imj5��I@����TZƂ_��%8˛_p�^����b�n��+g�����Ň y9�[����r��,���-����4��yC&Q/b�8\^LF��0FK8J>8���ki)~X���F��ii2h����ѻo_�Tرh�'xg��,��G? Z���\6��X�Nd�GJB\�"t��	6[1�6/N�:����`�'�"<*=z�Fǎ+Y:�y��H�|����W�_��P(R�|j�;��(b؋�'���}Ό��u�/X�t� ��Q+�.V�����a��DsTa񨝔�����ul�$���+��}���u�ͿmϦ-��1�������Oy�+t��	йbU�\�_��Y��do[
�(�F���W�R'�kmQ z��~��T��-'�)!6r�!�^��$��kH%�t��]�FG�C .� ����K���#��rU=GO*|>g5
Jʘ���V���X������ZT�M?~�����SRРA}L�6cƽ��?����bL~�=,�z=���ч��v"J���B.>+L:+�gԅ��V�Dl�Ǐ�Vƴm�Cl\>�l5ⓒ��^h׮]�����۾V�}�?b<��?c�(*|��֑;ą�ǎ���ձ/W��R�$�g�~��8w��{�N7�ˆ>2����ư��ڷhq�?{��W������U�̿q�ȇ>kͮ�9�9q$����s�2��墡+~uэFV���t	䲚cnA]�>�|yU����~7�'�f�-N.d�\�b�}���5�A6�Ԧ������b��B��kȅ y��MVV���/�S�Ղ�}�</>U湅��f�����C�̓���C�7�VQ�����>�n�Ը�X�.7�
�`������qo"�gF��	�%��|(VV�E��!2B��C��(�,f|��

�q��)t����S���M��x��c��̬e+��V��?n��
:��r�Ο]��D�'�9�)S���W���o{�h��5����D�q��h֬#|3r�v<=��ͳ�q�:{�5ྶ�C�f���׀�>e޼��߳��rŭ�>�����b5g��T���2���FiP��"�s�%�U�kKE:�muRV�r A�^KV�<���(�<����d�x��|&�o�/��W���L���R�L�R^�����}����δ�Qh�_� �^��tk&�0��z3~�{� �����hݸ,JQ	v���0�ˋ�����C���j���`W�֪8�PjE��p\Ӻ>ڷMG�zc��wqp�F�5LEaav�ڃ>�ABb-,�xRS�k��\��c�׃����5�k�_;�`�|S�lH�}ΥДD����a�D:7r�.�X�*�wc��ȼ&��q;�Jm���q��{&9G��vb��)/<խ}�F�
��v��Zo�������ʹE�2�ݽ���4��_���"Lg�y��v%tE�%��M� �+H������7݄<���/�겲��� �@q�\������Nۈ�"���g/�ݤ
]��%8�^���%K�\��J���j|�\T_����
�lm#Cs����' �qq+��氳��-w^��c�;�����W�89rΈ�\1�%
�k�^�"�"�(�� DQQ	J�9���LOO窮���k�8����SԮ�o`��Nթ�^g��Z���e@w��>v�Y�䒥�=����hݬku��+��i>t�]�	s�~�={a��C���#d�� �r7+��I��{��ѧGw�ز�V-B׮q`�1��{ }�=���lܰ�.7y�ɟtV��֎���xӝV_Ċ!����A_��L��骀N,���z��v�ڂş��7��W涵��Zܶ�d��P�z�{�{�G��7���mk�O�>u��y��	K�������P�[����(�Z�X�F�b�E����E4���x���v-"^�"U-��HD�z��z�[D��K��SD��A[d�¢z��{�9r��U�&q��B|^��N���%��,G�J��t:9��ؓ&�A��a�7Z"X�m��݀��N��+�Z����E���S�<������[o�]wu����s�Wlȯ�"�,Ģ/(A�[|�p�����zCQHY��y���[X��X�v#�R�p˭w�}��?ʸ��)���_�EFH,iP���E��4Аy������!C����q����O�����Te֭�{l*���8W�!2�X�{Fx�W�F����������p�~Y_����&-��|��G֗9IK?��_� i���il���UD�J�N�'�r�
F���E�[oP�Y[�c.���xE˔���v0�j+�b�&�o"�->+������U'؉}�
�d��Ы���1k�j*Td�ĢF�SV����	��*%�INI���\^XLj:�/QI��~�~�6H��R�-�=m2��<��?���#�DD�	���+V��1Sq(��n��F*2r`��С��p�f+d_	���>.^<�����bG���b��Ν{`��B��{�]�+t#�S�aU���	��{sK�b�Rݻ��� /Z-����o`İ�q��I̚>	����ذAS��y0Frۚ5����JN�7f��w��e���z��7��5��GH�>}Ł���I˦����^�>D���\NN���}�PtN�N��x� ���!}Y����zU���W���q�"J�ߔ	`,�+"x�rQ� j�W�-+�~�+���bדp�p|��zU?���qȋ�JeeeU�o4 �NQ8B��**�cw6kDN\���|'Hq>:*��"���z���<Я/"�����гgOXLV�\��<�(��`*��g�A��x��e�"ޢC�n�ЯϝhZ�!�K21�Ñ(+˅�̃¢R���{b*6n��Jq�﹏IqT��Q�TX)�7?W��q�� y�!�%#�����r�>�A�1)���fϘ���R��n�+����DN�?��k(�PТQ���<�D�m��/]����a@��^�j�E�,��?�!+7'q���1z�+�<�vE=�T�]RQ��oj阘�Jt��\ >�0�����5�XAQ��5WgW���."��M�#��"�.�����"�)|U�M��Szu������E,PDJ�z/�H�Ӿ	�)B�H�)
�6�N�/Kj?��wP��'3a�F������;�=����Q+=e奰G�'�*kӲ<.z��?JQ(�BPt!=^ؼ~��3�����@'+(�=��~�Ԥ(de��+	�X�QX��$$&�WϾh��
���y|-�	������1��S٥�� ���h��7Bmk�.j��c����8v�,�?W�o�k;^�:��M�άgON�KCG��lR��9�͗�4��C���]����~�3V�ِ����r���}$,�q���6u-Z���ip�Mix�N��
v��dEd+R�"2'*"E0\E:����
���~wQ� L��/�t*�4�E�^�ht���U�₍,X�t޴����kn���M�N7�=�z���h��5:kw�_���vc�׋�H��eճd,1�5#��)w����%�0j�l�q����aAaf�^	Z��t���=	�ع�{|4{n��	��fa��}x��ǡ��g�A��{��h}E�*�~0a@��;��z��^%>
m�G��O"���i��`��]L��� ���l�($%5�>t�9u&����r�7��Gz���.͵�G	��xU~�c3wn�k�m()u$~?w<�y�yx�=0�(
w1�K0�	�(:�n04A�# �/"�.k��EE� ,R��N�%"u�":&�2���S=y��Lm]������Qە��aTb�+S�� �48[���l"��9Ku�����x���c�*�-Eb��cdd$\�
j>��� >:�K����ǁ�9j�p�a�W���?�"P��UW_�-����W`�w�q��cԻ#��X�,�:�v���F��Yb�9E@��c�`�QVZ��[w�o���oW~�ظ���>�n����%@�k.��nOۏJ�{�~���%�B��@�4m-gQE��#��E�>�UL�4	�woe�Ԅ�(�l�!�e�!X��X�T֠B6�^z��<{w�m�w�����Ow�~�O����ԕ�7�'~7g�~�9�"�4t�ʉK�ã���D[���LD�y��ω�Б)��%d�o����^?$Y�DnhT�7@�s���l4r�vQ$�c�F��l2��z�>,6|� s�,�)��'�?,f�O�ޔ� �V�ԅ��G�:��J�VT�ynH��g*U�n/�|rr*��J�b�#��.�SI�#���f\r��� 3*ʋ���Ux�gwn_KM����c�� kD$�?֟U>��s�7	�2ra�GB	a#%;) ]��wH���Nt�zΜ8Ƌ�Ob!��t���3�����>��M	ԕͭX�	�������3PEH��V	*��@���<��������#�0�]��:�$'�Y�6��e�F'ë3A�!-7�5v�K=��M�������s��n��	Ч�ش)�� q�����0��n�	S�C�1"���E5d��	�(2'`usQ�}�>���)��!��)�˩�ʐ7��0[���$�t�(����h�tCSxa ���F�F�#���d�A��1�J�	p��ˌtWE9�f���,���)�$��	��E' ���X��&���j&"�����Ҳ�>u;3���π���]Q��}�G�܃H�>o)�.��lF�>}0a�46T?a:>�49^��C/z"�0BB�v-�L��k��}۰�d_<�����G�� )��]��������ѬY>'�v�r
���ʔȯ���o�=f�T��Bz-䐖���|Ⱥpo��:&M��u�W����e����HM���FP��'Nb��y��i��{�|�g��{\�?�>��n��'���ɬ5;7�%-�p�]�zUJ���sW�N��Ѹ`�U6�f��R����H�E�{Q�Oѹ�OUk����
�#��	|B:d�۫��b�|倪�N�D�����[̰F��O�G�~Y�0��/t!r\3�g�	&�^���CJ2 ��\i)��T��T$@;��q?���%(��h�YPRV���\.KX�Q�M0Z�0G�c�����G~n>�CnkO�f��)�������kq����܋�L��1b�UX�� �F+�����a�Q��<���Z��ρ/?����"�a箽��߃���Ǫ�k��Vw��ŀN��~}­k��Q�}�L�� 5��F� ��L����!;�&M��۠e�&�rK7�$ԃ���V�5���C�Fw�y�>m���Y~����[��<���|�����TXZ��d�����P(>	N'���6.Z�跈�E�-z�#](�����Z5��t��R�5N�u�\�h��:��&"�Z��$!��py��Z�DDEA*ʝp��"**!m&}QF�V#Ar���t)�,HMK���o�AYBI~!|�Rba�k@�sO@B�7 )��6^8Xmv�l,C`��M��T�V�;]U�#@��4
H��<��(h�F8=�y%\ȯ@P�Cyy�o\�޷����3gLF�֭Q�p�G���������s��� ���U�@��F� Ϊ�S���ӏ�I�@iq&Ο���d��c��-x�������_.���}�-Z��F���^����~�~�5DH%C�2-�*#t�~�ee���A���ѽ���i��]+�o����-2�)u�������|4�_o��7�սE�z�����;�S�@�������ؙ��Z�cK~qa��Gb������STL_$��~o�
G�L�.��X$8#Hr�U`E����j�U��z=�����e��0�4HK��AZ$��EG�#����f��B�kѰqSD�#�.w���S�XL��ѧ�-0�%�|D�&`٪���pK:4j�V��]�Ν:��$!�T�g��P$'���#��y�d�88+�����x��[�6>��'q�O�/����>���AEG�L:+,�N�{6�;�ՆPȏk�h�]k�C�8��=���6p�=H�UC�G�Ӈ����tV.�q	�EŢ�����N��v�v�M��/W 7��u�����b��=���v�׭��_.C\|��� Z�l���-ς��C�*��.����^��C^N���|�voƢ�seŭ7߄��Rl�~Q�u`��A�ӏOM���3�_���خi�?�������r�
�1���I�Y�wl-,-J�f�(��`$./G��~)PE:Lo�>��]^^�J�rz�ƀN��t-j�Ec�� Z,�vzoVVV�*��]�׉)��F�FqX��st��65����Ӱ%ă<Ү��jhe��E8{��=��mX��K�_�1�Sbp}�����>8}��lF�+�r?8)�9p �χ�h�lZ����8v�0����?[w���Ebr:"#��"��$��:������/F�b⑗�#3��z�Y�j`�Y�G.�-i���:�&��A����dFBR
J�m-��7��>"[�V+t�*-�͠�A�#�,��.@�@�ۯG����I2��7��u6Ʒ�W#!1}����V���@�A Ls�����{��ՆH�5�:�:T@ '+Ç����o�v,�f!�I)��{�ixa���@�D�MǮ�9n�W���Y�NtYM�Sxܚ��0����_��������5;�;JS(�>��w�,.�Z����Q��0J��`��::�� U����T��p��<�N5�����*�v�-77�����qA���f�ghUǄӨW�v�;�������"���\��?u!EB|j$��Z��3�Q�Hk� �o�sH��e�6�SJ��=0����i�e����Z�=�<�<6n��ي��ڈ���
!>>Ae�+�&G���	����GY�a�Y�W|,�K�^of@?�����.l��4��+)�A�Dz��_����!�~�rt"��..�����F�^A����/��9٧Q^���;�2)��_Ｃ;��>[�b����OV��TE<�E�!�~In��� b�n~ t�������@����yÆ��7���wc���hҰb##P�A�m��ne� f�%��(�MM�>�g��k��ۍu1��_|&�q�i+vn-()J]:et�S��_�F�Ή�N��h#�V�����2��}��!�R$�H� `I�nUɊ��χ��`PQ�����xﭗ�p�k��S���c��P���a�F&ë�h�:9ĩ��NA	��d��Y�n�|�hZ�7����p���>W^s%4z��z>    IDAT��V
"�
L�*�̘3}.^|e0^~k�9�,���$�A��zLl��z��o��k�z����7��&"�^ˀn$�͑��h�N7��;Q�kGyQ!�� B~^z�i��Ƣy��<ǯ����$-d���d�,6(n�r�����O?B����]�ZBX0o:r2Σ�܉��۝=P�qS,�t1�C�<�mk�W��!������_�6��2X�0F�[6	�5:=d��� �b���&�>.��gf�Q�4�k��[��z|���o�����2Q'%i�跞�}m��G^��z�a@��/��sp��}V���۶e䥮�>S�}Ia�T��ÀN�B�E�-ұ}�HN�����uy�؅9�4m��b-$��2��}�����ш��"/��������];݆��J��[���ç����z���#��E@���Ǫo���mlzҸU���i�Z i�����0��Pd�7oB���'˗NFl�ΜG��o��O����\C�G�2�'$&�"�"t5#��өN.���ΨJߺ*`4�]��PH�Hk���tZXb�a�1�C:�4F�=C_�&�j�Q���K�����q�7�Oaa!�����.��\,��\x�<���o9t:\s%�v3�/�oX������}*��٢b��K����>�(G�J�V5q�������{��3�SO�GD���!eh�G������_������#�3s"��p�7k�N��@g����)����G�!�f�9cě��7��C����/���������I��6��M{�:�i�r�6jJ�8�N=ܔ��v����	�	�	�i���6jA��,_��T���gh�� �ޓ��Se��p�"����c}�떶H��� ���ØY_C6F����Mz��
�q�t� �:/�{�h�8^g�*\�2m!J�Q��Ѿ�5�pJ�����9�0j=x��.hX?)��8w� �܀��r���T��%@���j�q�z���;��Lu��@�5�l4��r�+����i_f�0�p�l>�ee�p�8L��"I:ׁ#��W`ʔ)x���q��)�=�2.��}}o|��: �	I�`�hٷ���Y��p:�Q/Վ��hdd�`�����������/��#�=Q�r�0�_=}�j� BZ��e%-�~������˘0u2��)�M�O�8>k7�%6�΂3��(�H���=f���;�i�O�<.�%?�0�_�)��~0��z����ZXZ��Մ������:w��IO�J���Y���(Z��/t� W=2�\���:�&G2A*��Ɏ"xw�H��!.B�����K��Љggr](�*�z\ױ#�=���;E	@k
�i�4�D�x�WT�ܢ
����ƊVTC�[��;�nA�@�HO�":BmH��'�J�)z� 95���z�Qo��#XVTӂ#wz�QH��?x|nx$��b�T��m&9}8��DD\<J����x��c7��)��z��͝�	�зo_Ȓ��C��a�-9��y(�)ĺ�kp��Q��>�}cL4=����p_�gg0)�������Dlڸ��������>��c���z'�S���TG�/_�G�r���	��<����?d@���0h�����5���cD�
�h4�Ww����;�VS�27��E��a��yug�ڽ5�0?�X�K��A��,&yQm�X��5M����Ye���^��p:�7��^�8Z �����.�*���EEŰ�m�i��d��u �q���#�1�"�E�ƍa2!y|(�/ 42�V=l-t: HZ�0��<�%z�V������b���D����#'+fK۞ju&d�ѱ��F��p�	�e����w  s�N�qt>Ծ���P�(�s�������12g�P�zd���o���}��U�����~m۴��bƝwޅ��xu�߰=~�o������9܍д~�Kгǝ�.�Ņ'Тavl�茐� �{�%��b��}pVxЛ7o��2©3��������.�#uLH~d�;π��عk̟���	q�ԩ+m���ؾ����d@O���>��7����K�{W��r���Иٟ֙�z��2Wy���`���Q�WȪh���Z��T� N*����"O`���]����W����)��O0�H��rj^%��a��H
F�	f{r��e��_3E�+�4Ğ�@R|)�)�$mv��i*܀-"Ί
�m5M������\�.hu������hɺ��e�p8UG,
�����o�e��9�F����(s����	:�{�π�3@��0}�<����Bh޼>�>'Jʊ�V���
�����f��'���_z#����/b��X�h!�N��u+�E�:�К(/�×��Y\ �ۇ�k���G|r*��>�3g/��$,��Z���������#tJ�O�9�����!�4���xԭ��x:[$�O���:�zi��f����m6,��/|�~�O����K>���k�Z��X�>o�8
K��R���@�Nx���\��	;UA���>���wѯN���VU|N�xU�u-�0��ϋ6T1YT��VZ�r=�$2e	V�f���!҉�K��f����n�9f8�:ؾ4�h� J�J���^7�����	�
��Z�|���t�����R�����h6���,��#�VzhZ������
�LV@�bŒ�1m�8��D[p���m؀翸ȁ&M������9���Y�L�.	�$#!6�O���M�`��	z`1q��n�f���3g�f���Տ���
K0�ͷXX���8�^ٺv�o����c�+!����!�b�q�'�R���ѹ�5�Mп��D�2�{CZ;�Iq�q1��?��]:�*O��s�7��S�~Vkښm�2r�j}9n�}2�*�.�⸷���T�НN'G�������~�"���	�q:2^�~t�~��oA�#��A�֫��R�z���$pYS^����J����g��T����!Lo���(��� ���j��kz�No}�R��B�}�
i�]��O%�O�g�X*���-��)����xVX\����(f���
;���ь���ѣ�m8�g;Z4����
�b�`�F����_�5�v!`�#&!�N��.X�zvik���7^	��\�e"��a�J�綵%K�e-w"�}���,&���/WS��A~���Yj��� =��*�����{#p��n̙=	7tꀮ7݈]�!"�6��@�_��Ukp"��	G�|�֎�څ��j����a@����$��?kV������;k:�-|��|;p�S�D�S]ш�f�Y���?&&F�&���W�|g�2��C���"UD��9��� ݉8��đ.��(:&Os�Q%$��j���v�� �$^pP�L�˖����*'f:��T�W��IT���D=�"�
��u۵$�A�ٴE���/#2*�[e�+�Nz�t��)�Z"�;Y��v���}���%��X�QvlQX�a�=K���m��e+DYM��<�̈́��h�8�a��@�:s$V��kZmh��;=�N������Ipg�f7��q��a��m�w��	���>�,v|��:�}2^}�ut�B�`O�V�A'e2:��V33 X$�]����k^V&�y����G�q�=)1j�B�-���l�;��#dO����{�ΰ�Z�\��a�0�_W�>�S�֚�q�ֲ���+gLƒ��bߎ휾&��Py��Ȣ�ˑ'1�	�9M��dj�M�k�BDC��E$N���u��w��FѮQG=ު�*����,գ=� �����v�f�r���������s{�G%��}ު�;�Gm+��A��Y��2l�*��7��HF��+���"�����+��)·X�88��$R3iU��(���%�;g\��pA�񂣴��7E�׋R���#'���c`�G��,���:EF�F��S��(�&=�B���9�.p!���z'5n��|�Éw��,wġ��@�p��-y���|�w��3@j�� 1%H$5���B���@>�wl¢����v !2m[����(��� 0F#%!z���_�um۰����~����s�}æmY����?�V���͛$�5���B��@[ 7TYY���Cit"�	���@O�c�2�~�H^��п���@���hL�V�U��AqIby\J�GXmPB�j�j2� �)�NNh:�J�#���J��h�����%�������8Z��3������` ��),$�`��A�T�'�w���h)�O /#�nCv�g�=@Oa�_��?� �
��v��KZ�!�/�6 K�m��Bb�k��(�F%�(����܉�����4�:qK�/���ǡ(!�;���=� !>��Z��AC���f͚U:/��笆X������v�DI�Z!R�g~HQn���1���_��(n�tn����d���7��B��k�m�����xu����ey����
�?�5>¤Yҧ�Y�=�����qc�m�R���i���ZW% %Pus��E��Hn��\0�YN �`��>��x�_WJ���:פI^�T�t:O���Ft���.����Nrt����Ո�"��z<��d�қ��(/wTF�Z�D�^x*'���b�G�)&,&kUƂ�EoвY��@Y��-V	�k�JG���
/�Ng�F�$(�!_(��l�� ���z����B����+�@RT4RRR0��7q��Q�1tVl܆CY�0E��窀��M�1������ְXM(/��'󧰶=-2�l݉;�u�5"k�mD^~!�5M�5��>��
���׋:­�5����(�%Z��F��Qav6�~C�z'OŜ��ѶMt�r+Z5o����(q�0'$��3�d�v������=�mk5v9k|�0���%��`ܴ�is���^ꬨ�d�,�d.vo�3���p'P&���iv�?h��isU��j�ԓ�Q�.Τ:��:�
��_A��}�S�b2s���,��n��X� V�Q�v�V��,����S�ܪ�����왧ł��F�R]����nR�}�&����Tӧ4�ڲ��sTk��-dbc���^�qqq�i5�z�י b�ktL�#�/CD6� �M���/��GBBLײ�c�����ګ(s�c��͘8e*6�9�o6�CdB���p��Ѕd�!�A�cG�ň���̉#qk��زu9���܎��TtZ����+hڼg(�A�v��(6��{x��i�PC4$� �/
��0x������ν��G�^w )*'��F�>�¯��\�-^�Y%����;i��=�)���5>p�k���0���Rg�ܴ3����cFs�N��#�:E�������ggg��z��q�Z�	l�f;�i���*�]�DU�E�p" b��)�P���r��yj#?q���r�lF-=���|D��n��	��c�=2.��A���@�dZ|~��l�(-�٨��jf`B�J%�Փ�f�<WS��{��̆*=¡yr8ʑ������iC������4_�مe�,A�t�`�ү8�i5����ے���s����/�ơ�G����X�u?],ETb-������2�r��*�ݰ�l(*����BN�9DFD��oW���BrR��f9�~CA�&͙�_}�8�0������ ]G�N�I��%EB^F�O��C�ٷ�fMB��uqC���*�`���H���Ɇ�R`OD\����a��ݹU���;���59a@��ٿDc���r��bGy�GÇ���رi#����Q� �"eJ1Ʒ`xWW�c��S�+���.�sJ�ӾH�R�QQ^έf���#l{d,���2�L���)j�=(�`҇Դ�^g���U(=O M�p:~"ӑMkH������Jw9R�sy|0��(-u@�'g5U����hLe9��U���$4��N:n2�	jX܆#t����q"�!�e��f�2��³�p�~<��;�FBr�L���m�K���m{��hV��H��$�;��lF�(�������uq�q��~8�.�#�qW��hP�1�._����{�7��Ss/�*#�0�_��g�	�d.3}A�� �	�Fa@��0{�,:�̓pB')�pյ��4 "���!���L���a-����5=r�k�
\��'��,u�����>:E�k��k�0������`�S
� ��M�����j�]��B)mՉL�ګ��ɍ�C�+�~2.�GE��G��ud�Q���֠��+�`�"MV4o���̭qy9Y���hҨ1�L������֓fk���+"��8����y�����㢱a�w(.�c�'�6ۣ���.p�<l3JlcZЂ�T�h��dd�t=��DǢ����YV$DE�Bb�9U�f2"*!���KD4��x����3�*кy3ȒEE�� �FD�^�ǟ,�K�`�LX����^RT )�y���hݢ!4z�?~?��{��b@w�}���;�V�.�o؂�F����7m�}��3(a2�%x���!�E�.��V���{�"��2f̘����3&0)�_����z��k� �nS8{�M��|������<���7_�6�:������/xQzJ�g|������/de���h.ϙ��{� ���P�l�2U�=��W�(�T����X����Y���eg2�����ϝ�N���"(�v�JX-�R�� ))	3f���)Sٟ��N�X��aŦ�P$=-˾��Y�a�r��$co���� :\{+�p9tNG��N��U�p��Q^<hu:�'�B�N7����n�������js-]�)wJ���]PR8�N$8����<z����H�j�[H
 ��g
<(شtJ ���A�z�k�۝�s���k?�1A%�cT"\�XDŧ�2XyI!,=��m��#}0y�H|��صs=Nކ�H+�^�_���1D�%�o�#2*��V��t8*�</�:U�>���hCL���Y'���"��x�Uv⻐q�&��bD���M�@�F���k ��=u�D[��f�x�G8B���Y�����~3>�*e܊U��k�|s0
N÷_�D0B%ӛ�q�Q�]��'''37�S�NUi�S�n�[�z̅����W�[d:��'�_����lټQ�&�H�y7aͺx󭡰ڣq��1�Z�_��#�Maт�(-Ƞ2;���m�k��̀~�wB��?�o/
��P�N:6�����AO-f
4j���q��]��Jց�sW�����(�N�:?j��l��CAP��/Sﰖ�ZRH%B�=V�<�)w��2g�:�Vj
�>�?]�Vm�`ʴ�о�T�D�i���}^�fì� ڤE�h=4�Ǝ�pb�GSѮus?y
�6lēO<I��?
�������4��s��r�E&F��2��f����C�$��H�ɀSG�`�ȑ=r�ރgM�-];�VR
⒑��щ�a�O��／GΡ~���^~�{��5���5<p�i��p)����%k���<u��}�[֭�v%���ALU���X�*�~�%��R��v��I~��)B����f��U?+LLպ��D'Z���}�V���U��;�AC2���-�����ɧ�FL\n���eL&|��b~_��M���yp�@	XS�n�&�~9�����B/t�Ǐ�����W,�
�Ng@'Q���zܻ}��y���u��g����y"�Q-��uh��em��"� �(�Nj_:�Yu�SHJ������`��J��"���''!&.=z��_���зa��C���t�̉ḧ0�q���t@�-G�]����iצ)��M0�d��c��x��g�L���\S'�����a�[�TJ�Z����c�����h��W�F@��F����q�`|0�}d�^����ЪeC�����7Kףn��p�@����6t`ƈ�m8��w���7��ݟ2�    IDAT\C_�v��������q��P� �SUN ��.�_�Ujm�ni�v���`�>��*FW�RU�5B� ]�00V��W�X9����WU�#
EAQ���܃��D�r�,�b4����/y�ѲE3̛5�Y��F���7�U:B��q�]wW�՝={�A�E�F�f�"d_<�&��q�-
O������7ue�T�A��,&�՚?��+���S	�5J�	{�0���-jt|Vr[�Fbϙ|��!9V��c�֍�km7����o0�<\��z��������P2�X�!�f2��(��D�UMy.�J�]�]����8}������{�j�ĩ��PV�°!����e>~E����	a�{�}�S���2{
��t�?yo|�&M¶]�1}�$��a�Ьi+|�dK�Z��%���4�JI�9��z]߾}�>��.k�����K38��u����x�pdُ/|#��p�X� *��X>է��&@��N�8&��t��;1��@��6�S�)�#f�uz?m�V,�����ka4�E�z�����nꂴZ����mӂcْo��xe�v�9c*J�	)�i^�n]t��3����X��;���ً+۵��?F���@H��ߠ	���sX�n=:u�����j���Sp��� ��
z�͊@P���L�ɪ�<zHoƎ�����a��U�������Cs�Έ���������l}g6�:�=�
У-&��!P^�Y��:��KO=΋��<zb��39C�����2`�ν��<�M$&���3��
_;*T��.�M�̀ t�@p���+{@��'Or�}�ȑؽ~�1��V�}z��)���Ł��h��ȫ�vr�ι�Ѫ~������~����??m���W� =��,�hLt�2�nB&Ux�S$N1�����H�](��MVDDG��Q�����2� ]��Eݖ ���b�7�zʱe�z�F��\�� ��;u�������.^��n�Rt��cǌ����{�5:���G�>(*)�m�w�z���38t� ���̘6/��Ť��'��a�!X�v���:�c7�̐d����bFe�1����	i!�u;�7�����M��zP�a|�� �_&�,Ŵɣ1����./�3O=�V͛q��nÖ;1m�t2��ea��,�bS�ҋ��0-3�C��D�=�߁�� �W�_���[Ы�}hw�՘>{��_|�5^Q�>1�%Y%�_�9!:���Cp�":�
r'H�|tR�;�ofM�����������L�h�m�4G�+�F���P��q�>y�,�n3j''�>�a����b_�C
�%��� }�-�.w��?xǶobR���E�L)r}S�"!	+�]	tE*����&52'�ur��P�"3?h���2�[��א$7��
�ˍzr)}M�`O>�����ՓA��vlGaa>�v�'�%Ejk]�GE�wG���w��~��N���=�йs'����8z�0�3oTT4�.Y��[����7�J&'�2�F)Q�\P����P����lM�n��&��-/�#�^C,�t��⃮2|8a��*ʊ@�CB��:`��}x���L��(�ݹ_�������[a6���CJ|�ʤ���7�G��X��v�jt��f���^̞;����y��@o�@�F4A5�N�t����z8	�)�NϚF��5��-[0o�2�k��{7u��6����nŅ�RD$�a΢����YD�{g��r�vM���Sk����a@��+p	Ɵ6���	+���p��,xo.܃�_~����W˼�<fh�yWAjf-BA��sZ�#�p�2��z!TC�gkS6P�A>vْ��x�3{:6�[�R��Y�Y��O�����.�܂��2>��;w 77}���e�E�L�3�������G��}�$fO�8�����W���SG�<y�!���n��,]���މ����%�dU�\�{�|>���5"4�\N��WAg��3/n�r�h���Y�GD������.�c������SкeS:{����Y����Ͼ��N`���u64�9q���Ï�(=n��	�YYȾx��7@�fPTX���v���7�;�c��i0[�x���HM��z���\�N���_/���PT�^&_ ��A�qw���Y�1꽑(sa��ב^;���͛�##�	��Vt�s�, h@����7mPo�;�=�#�r��kZ�#�����%�X�S�n؞[XXg��W�s�aδa�X�lF�؇�ku�&�7��N�I ä8�ۍ���RT����:M�����X��#��/�#::�%`�R ���?q2̖t��3��X��;dd\��?�F��(e7R���m;v���㸻{OU��b���ؾO?�͛5Av�E>�~u�<HI��ѣ�ছoA|BA���U�?���/R��|/ ^)�z*����6����rs�M�~�قF-Zc�����������YR �<�ЃHIM@qq!Gc��x��*v㛍��
�F5�,���A/b,2��2�'��.E��Q�w��i���qM�Nx������G믶�i�[O b�S������K���!�f��{I!�B~���;ƀN��{��0� �N��u㫥k������`�L�d�BRL��٣_�����%���À^��i������+�ߞSPPg��7ql�&l۴f�����S�{�nDGG1��"���V�����mC5����Q�&m�wo�Ͽ�s��{+S���6��FEEa��i�k�X��2̞9Q��A?�S�&L��`H����zxѰe�f��f�чB����r: �0Y�l�Bl��{�������gegb��%0�4�_Ξa�P"��Ux��1���pw�ް�#95M��ܜ>J�	�� d?��5ݓ������hݖ������j-}�	�����
�^���)q�(*-FI�I	q�*�ko茷��Ć�9��"��������@jGkpU�FhҨ)�%��=���N���	�hղ={�|0v�ԯ���!%�64Z@�^A�\H,}&ʑ%G@\�_sW���;q&����(��M[�������Ou#���Y��W}~�O����s�Ӛ��"�U`�j��.,�d������%
�����N]��ި%�����7z|L�у�ug端k��҅�����腭~Z�r_�z{��Y��1c���j�2fJ�v:��Į]����Dfz�&9Y��lGJ_B�f�h�f��F*l�j���
E��wѲ���ɸ%�F�Zܞ
��⯾������_���!>!�Ǡ�7i܌AIo��G�ޜ.��z��u(*.���?�v�ڢ����g��[�;���O������kZ��:q���F��=��~��qzG�e�^�=���oѪU+�����$�:�\p��,����o�6(�%�?����V�Y���<&,}�y'����i���{��Yú��E<�����ð��0}(*�G\r
Vlއ-ǊP��3$��fRl��wu�խ㚫:`�Uسs=��28�޵�u�|���3=�܃��Z�j,�A��u�PPmd繟 zu��E@�v��7�����~]j@��������- ����CAJ��bXG�C )X�N�#;�b��Y3~֬_����A�d��W͛�F����H���w�L���a5i�=�g���3~�8ï�5g�>O�Y����
�kv���:b<y����T��I���_B
��ك��xv��E%��b1f��&P�٦�Ѩ�͠��3N	r4O��S��]ڟ��SI#݊3'O��u�>���a�T���H���#,YZ�~}x�>x�>���z�Ma�1E�_�գ���|�����[RR���MZ�����H�MK`�pV�J�jדf�_e��Ε�	�zph=C֯����u;s?��+$���7��]P�iɋ1����飸��~x��GѨe+�uZ\ۺ9��֮�'_x�rdH�X(d�*�`�}��`���µW��RA�]�%��Dq�9�����[z!)�V~�
�o�v
��Cse�����΀BER�̲"#��m���H�r�# ���I�ߴ���z�M��Oq�?�� tr����t�S$Dz�ļ��{�a��q7y"�o\�%�~�����-�"11��4��0G����r�6D��f�?⮰}�o�#�������w?i�W��V��[PR���С(>wϝ���H�s��2��=55E^��=���j�yRdM���h��C6�*K�l��� ���$�Ϡ+ QBmU*_K�ݕLrY
p$�ѳÉ��h�%	T����j�{����U���鋞#y�PK��	y,���臅_�d<##�h��K=<9���B�9��U;����dY��������4t�ԣ�5�0n�B�-�����-+��7^�7�?èw��k��I�ֈ����E�v���/£����"h�C���>xOa.�?��
��II�8�gt��nR���X�j5���+0mؼm+n��V�n��I����:� t������_�,g
��������[#t2��-�/e0~n.���B���@��_a��_�C�Upr�!����;zr��1s�$%�`�s/`���U�C��m��e�AdU Ƣ?2y��ulf���k�g��o����g�7:���}Vk�Wkv��ޔ%��c��eX�rG�D��h:2:
[�nE��yf��F$5YQ�ZHj���e��f����� I�9��meݙ�WE�9�;�UҲL0�eURV��$�ٷ���5E
��<��ͩ����%D]`Vի+{�	��>�I��t�t�9���F6v��KKKa�?@��YR���8) ��΋�>��_7���������3gpE�kx��6#�ݕ�#�nc��YA�� ���}�tC���0'�W]��W�C~�9���K(p80~��X�/^�^��W�Pʝ�{�a�J��=���\�N�6C�Z������C���C� *&�6mD��;��uF\b
B��
q����������F����P�Տ ��&�߂:�|��� �'�7l���=柜�OFW��������V������q:�C+� ���c�3*:v�����`�"��t("* "*'8�k���}���׹�y��\���Q{�����}�����vN�y�k{�H@��m6㩑#1�՗��j&��\.}z�BKDÊ;�]p�Ϙ�>�?��ܽCN�۷�8%m�7>m��o|�~뮏�8�lԧ��jhii���/�y�n��]��	x9A|��W�ҭ�OA$��e;��רMM����|��#��G,�`����g6;�膁H8����mP'����n�;x{�L��^h�A��N��T����(���հ#_���ɞ׬�w: �Ty�Q���y;�y������nz��*�`�: �D����`��������**����1l޴g�ٓ�MőW�_}�#I��r�.t�TE̢����2,TWQ�����B�2��j5���deX�7"��mG�Àjf�I$QT��_��1c�G4f��s��=�w�/�i���>}�!7���p�f� @�����B����k7ܯ �����{�����~��I��~�X��c��=������[�qkz!-�haEeze�$$���u�1���ĳOcc��h�jQ,��g]���@�汿�)9 :ЕݓF�?�-m���5�w�����^۟�l��S;�8��ʚ��F��n�ˣ^`��Vorr+[�z5r�m-�%�޽;�9�8�DY�E,�{��$U��cb2g�4�Ku!� �x:���3��5�*?�,���)�ԩ��fR��4S��9���4$
d8�1�S���TuR��t�4�l�I�cܺo����*��i�@�Nb���dbc/RH���0H�vKKK� h�ۋ�@,�~�-�/_�G��s�nt�݊7t޶��p�Q�����×[�P}=ƍy[�Y����� �H"��g���⮺�ZL��_��	�D:�.7�pF2
!�	Y��[��C�`Ѣi���E*���}�GYY,X� \t1��w4rra�t�l�;�L;5�P���uh�&�W�"���_��#��o�_��M��;�NķVP線l�m��ϱ̿l),d����U�1v��x��g�����⹼��(>t?b >�x	do>$⸨.��9��ؽ'�<�g���!�\��Cl�C�¿9yv���,�vX��{X4�#�X���A�,����&�U�ٱ$�w��z�:�4�����:lذ����E�0}! T�*�B,��А�=�������M M�z�
�Z& Z�&�YśL��V$U0�N���Dr#���p!k�?e�[ݴ��;�D�x�@/2y��UL{q�Nqg�����y�M�{�?���HfYp(��g͚eW�Z�'�|*�.��J�4D���{̉���W�h������F�����
�p�#�����v֣?��sغ�����@�¦&x9i�m�!B��=^�?|-f�z�9��X���X�=A,��k�{�yx�q��-�����se�	rF�&����7U���}p������������ڷ�8�׀�o��~��b�/�G��ph��~��Vr1܉�B�$�da��x�	>�ql��f6�y�$\{���' WDU\����jU���C�O��c�?~F�>��|� ������}5������Z�&;Ž=�M8ԟ]�HN@U]Sǀ�H�p�עW�^̭�g�-��5�Q% *(�C��q.�m!kZ�NlxjM��0-&�Ѭ��h��ry�L��5�6���*�t�g��ļ��:m�l\sssA@-+�"�씪�v T�j�5��Cu�l�B�I�B�"�ыg�T��:����y1CU:-4HOߥK���-�F�2��:�V��cΚ:o���G�б�]D���~���@&�'3����/C,܄�n��p��wvlۆiS�bѢE��?cgy|�	I��N>��d)IH@7R�>����sf�ǖ�^�=��G��ݰp�B\�(��>_��؀h4�5dsz��o��;�V�`�o~�)�\�ߴ(�����η�=�ϋ��>�����x�T�
��`d��~�&��}�1l/߅y_͇%�hj��ҡ���'��_ԑ=�%E�a�(p���=��O��&[��y����U��ϟ��7����.�X�|OEE�i�=D����#?/�[�,Cs��c���I1��O<�D����'@�9�i޾C)��$=̩�&}-�-�� Ϧ�n�S�m/������mrA`�-2�rL%3���f&��΋�@��e��.@V�t���s�-�����f�ی}�o"�i����j(�é�<��������,����hq�a���m"�N&�ѹr����tVC~^�m��J0�^U��3 S/��:�E��=}n�y�-��\�\�]x>v��Ì������K/�֝��c5L�I]�%��@0��efy��RҸq���f�b�^�p�[�^(�-Ŋ+��?\�3tt����GV,PC0	���/���; L��W��|�Y<���~u~;����m@�tJ�S�g-{<dd`e�ؾ�[n����U��9���0�g�;�ޒn�_���0�P��w�|��>{�w������>m��?}��l����v��ҕU���>�,ʷl��I����9������K������������/�%R�����՟��2۬��x�ގ�"6;�";i�utpj�Ӭ�@�@�gϦα�.b-��oZְ���bڱ�n��A8����u،v��әb�ڼ�U��G4��|>d�o���:�Z 45���g�-2���ق�8D�ˣP"��[�"	��vچ:��0�/����M��t
ޞ3������h�x�z
9>�r��{do����5h��q�E��1��WA�`�"dU
|IB�RM���!��^���e����z�w��9s���u�]�n�S�    IDAT�	Щ�$:�:����A��3߿�ҦE����o������߲�����ؠ�n��S�+8~�f=^y�E��vV�Ŕ��0��Jqí��s��W�"��|�8Q=���N2���m��:��@��|�;�;��d�ʖh��e��]�S&C���cSe����r�gN֪]�ve����^�r߽c'K�|� T���8���~E����453�2N�5�����^d.�Tl?x=K^��ӨZ����V��#�LrZmTj�S�:�C��oj��NkYTP��4�L�er�!әH4�3|	��(��ʻC�ܭ �!E 1�]��2�ݻv�1H���Ʉ�ew�z�?3�XQqC��1��	���?"�KY&���;���� I㖻��_F<���/ߌ4hF"��B'� R�L�e�%�q�%�i���pѓz�J�`ٲe8묳0p�q��r`����2�ߥ���:�*��_���ҹ�#fm.�='�$:�!���_�b�b���ݤ�V[֬���g@ߵf̛�? ��ǉ�^�?���ȦXupǫ�a֎q��C�ﵻ��g�������O:���puc(����KK�����1=�	ԉ`Fd7�?hϴ5�����Ќ� ��TWW���n�����U�y�L9�d�B��Xj��yA@��Ɩf�&I���2��ND"!���҂�dp��\��:Wܙ���f��/u�Śl@C��T�g�,J��H��,�#�u~nD�b`�����^uA�i�or%��$��Mr��?G��n�o޴�G=x$PX�����5�x8�G�G�@��0��]��Hǚ1��Q��`f"�;�������/AEu�ʛK��2-]�@�)�g�<�,���4l޴N�&q�Q��{ >�l��|�aH�pmC��1h>�ǳ֪�������
�������r���=����/[�6��ω��Ǌ�FM
����ͫ�`��W0|䣨j�Ƭ�3!�i��ǵ7݇�މ@QWXa�ڶ�����'�8������<�m{�Ϟ�6@�g�����͘��噟��onn��#� �P��y.��>��t
{��AN^?ZZ��m���oW��� GGlpbd��L���1"���h��f�suz�*�Td�Inó<���N��m����Fv�I��I�KD�t��c2�q(2W��X�� MmGͤD7�x�u��bG�i"�Q����Q[_y�����O�i�n���c��U�D�����A"���gr��3-r�t=n��L~�&2)G�Ϝ���d�X�Ȇ�#�v��/>���}��uM	\����B%����რ�$}�nJ�Q�$e`d�PD>o7�x֬�>��[*��uG��ݰ`�\������!�σaR���47�A�B�Z*�'@��g������_T��lU��'��?i��/���m�NL��^��y'���Z �_�L��·kV�Ï�ǽ߇��嘳p&��fF���������#'#Hr��z܈[N��I�f�����_�m���9��_���ٳۿ2��5�r�9j6-]�%�?窘f�Ty9gÆ�JzH����l��AEn=�������Cgdu��]���I�:�%u���������Y6��g]#KR���;y�9-����j�����-�H�s�v�gm���v�+�!��*|쎲���<R�;>$"!8�DRYT�����癴���K���|Ĩoe�/�tn���z�&���Rw�[���!cfl�}<���;�L��/jV��IB�����8�gO<5�$"5��Z��N�x�%�� ,g ������蜕 �)�c�,�iO*x<��mx��бC�"i��9�z��k���������R���%Hmp����~0���7~���.�(��!����?���g�7�ϕ�C���~	���v���٩i?����]����v��Z$�X�A�eJ��Nݠ��Vr���߈��*��t*�9Z��m�j2r�+��e����f��;��O9�o�l����֟l�����v��_���zMum]��c^��m���)"77A7A>�iJ��{xn�L2���:
���M@+��o˴��v��	C�`�N�@��K�w#�"Ǳ�e`�[�1j�(l۱��<D�	�T��+�D4����IgT�Μ=[�~HNH7�^?�2���Mr4+��EI��5�-���1����n��' M�xnn��H��p�5W㼳����61C���{0u�9H��p��d��]�>�tV�tPT�CǼy���X�����^���L��W �P�%Ņ�47�{����d5$�)�C�S�����4N>v �����r�b���x��H�2�:�����b�;y�ӌ�x
Ґ-��p�1\u������p�"���#���,��+x,�;�8th�	W z�g[��ׁ,d@?k��%��q���7���-)���.�}�~����̭l��+�V�{ �:��{(�k� [���B�qL���G��{~��_������/#��p?�
�Ց���v�^4�2<&`����(JģX��K̜5�]s95�is>��raOy��#��;L�ÀN�<G�V���]'���������� ��ε��G2~ƌ��3�il�����d<7�x��,�����솟6������ÝK g�drkKe��Ѐ�߬C�@F$���GR*��O�Ul~ ����x^�uע��	JQ	W�Ł\�"a$�t(��ݷ]���C$����y5u-��k���GV�ÒT��!��,��^�����|\�`a��}x�T�oj���C�� ���RУ���Å���O�Pųc�.���������!�18��*��?�yPANw18$�֮D]}���	�ˏX�D��Btz�Y:�N\�����������&�{���8�UxEg7W\|�F�Á���/��˯����5{��}6xRD-=��$iJA�,(䏟mƝם��?����<����w?�?�
��t`e���P�H%�:��2)�)����ߞ�t6"��Bq�����h_Z�j r�� �ܑ��R���]*wk�o@c��:��~�/>��;D��D?2ҍ,�浒�n���(m�d��C��`g?�ݭ�mJDX0H�g�wDI�{�#HI���Dv�^t�o����%du���O�'B����.-.9XH�g�8���?dck��1�aP�
).�p��Yg���G^NY�h�
ꖆ���!�J�&L�Īe+1g�L�p���f�.�������q���p�_FÛ[�����E6���kV��Н��l������b��~���_��ٚPK�d���X�r)�L�ɡB�-D[�aXD3��J��% ���{�[D<����F<�����}(��EC$���`��D2(zH�:2Z�L+�	�0Ϗ9Ӧ���/B](-��x.S��킠��RV�?]�p$ꫫЩ�=�8�<��(�_�5�ʁ��B��n'R-5�xp?��Ͻ��w|x�1X��lٱ��Bh�Y)�+��������b�7k�j����3�%K���[o��HF��W��םr�	����
<�����p���Pֱ��q+���~��_�D:�d��>x[��c>X �D"�����#�C�Sı����K/���}�R.��ձo��n@TW���������'�M�"A�d:�p��x莋���w�v˜5߫���Ю3|����	7��N����5Ȓ��be���� �w�Ѹ��wH���E�w�.6�!��hn!M���3�0����u�l$D#� &�����Y�@�d�K]���<�cI�w�yX�dK���p���Éw���J�@�>C2Hb�Ӌ�O���Y�II~HUj�V��&k���������uAE%�H^�a���2h���w&���<&cR\o�>}x�4�!wE�WRo�^�{��Q�"������pyx!&(����5<nv[�cb��zhV����q�-;a�u,�b9>�7��B�>�Nò�HDǣO�Ņ���WSU�+�%2(t����o=�������_;�6@?.��3>������[�%��~�5��g�cL�!�&�2z`	z�:v�H����>�'��3�e���uH���o����U7݂�."k��L�=?�t�3q�V
ss���a��Y�q�UX�a���ږ�t�
��4��0q���밎p�v�#������;��TH�bxr��P#тsO��������2�>{6�۲{���S����-�+�h��9Ca˪���[o�2�~۶m������-@��=ك��v^'r(�2`fR�,���a���1��x�I#Q_~)����`?�S�&|��<?�e�����F]���t:�|��P2iӽ��u8D�d��������ո��Q�żo�!#���H  ��=1��Cc[ڧz<x���|�$��N8d:w�N���bB��-s[���S���fhH��H'ȥ�O�ْ7�L�9�-�#7'Ǯ�@U���E\�fCt"�eY�GF@D,�ʘ:v������{_��0O���rNj	���?�ҹ�����Ug;�ٳ�H�����$����������'���������+@&C�Ĺ�cw(���`�!/j��Z��ڗ����x��me��L�ڷg�O�3vڠf?���Eu!�A�~FEB���Q����fB�=�-�`;$�c	(��v�z0��������҅��ı���ӣ&qG���y��z���o<��!��t��s��ы���wz��kC�o��Sŵ����)\�^&�Y"܄�{��I�3=�.]�`����6�X$��@eU5�KK���_#��C3E�p2���H�c��U�_��<Lz�m\z��'���J2�]>d"ax��U↫��c��� F���ߛ�P$���*͘H
^XT��R5ѫC }{t����dA3u4�B�:e&��"�WQO����0����{2�F>6j�Jb����:��C(�!�1�p�Q\\����@ia�����u��vXw<��s��b((*B4�cky-<yܪ�J~��I���t�[�$��U;���9��W �\��������F]K6~��w���ކ�HsW����V2�X&W�
�"p�6�؏;o8˾���� 􌎒�2?h0���=�L*���`�s&Mmh���6�Gt�el}M-���d��y�l�K�L�OcuQ��=`�K�r�0�H��ʗ��~���Ӷ�ȒtM	dmU��
z/�)�g��'âVo��E;�e��=�'i�A�:��P�����&)#6i{�` �h����F1�ċ �ے�"�E�a:�!	#''��-Ѥ��{��0WޡP3G��y��9'��<v��e�-Lh\D�Kc�g Ny$Pׁ��D����� �t�΅H#�MBϤ9�H4$^0��;�e�&�Y��)Crp�u�����������X
y�lØ�7�p֐��t�賾�B?.�;�gw5e����p��>��=;0�ѐ����h<͕����؞�q��	th_�)3��3QxV^����~��B̤�X�B�YQ�!��JD�]^X����|:g2�?�\T��!������Izv)�����ASCrA����ٛ+�]���g_Bu(��H_ ���sNF�#�1�xou9:u�#��B�)�'G<�m�*��I�%C�����ki�e�յ�ؽ{7���c��/X�[~��m;�[�n���U��ODca���`����ѫ'W���|4���jIA� )"�k�1�z�:���|(� �ZLx�E<����TW`���q�����sG�47�#���mxf�S�no5���xd��!+Y.Ju1t�����
���oD�i7� ~����ر������z]\%�C� s�v 7IJn���y��n#k�,��$�)�t���Ģ��d��ٻ �\�T'i^_���T�����|U��Y��O��}dD�wrhFm��lt �r�[e��T�3��"�,�Pe�E,�d�`�T�d8�������ar+� ���*d�G�4���<g'K�H4�����@�D$$�>�8�H��U>��5j�x�IN�ڊS�LZ`PG��x��,h��I�@�8Ŷ8VtZ6�����CU(C�t���ǽ���Mp{�M:���q'\�[�x
�� �p�<6�+٦��m�YC�n�C��V���Hqo}�|mm}Kɔѣ�o�6�x�i��d��h�$\���"�JF�:����[e�UN-M!��77���!a	�C���řA)�x"A�PTP���<̝=w\wV��%=z�1E��f�/���^x���a�7�WP��6�����'���������P,���>S�y	�mX�����c��u8��SqΙ��%�X�ŗ��OJ⚆��aʴ��u=��I,��0�D��|�O �L��t��MCN9��&ܾ���e˖@u;�qV�Ct!(A}Șn�����_��ɓ1w�F@r!��b�p��D��
s�p�J:���%�]U50O<6�*0m�;���J�ީ�m�cf�L&�����1��[�ł)���0�^��C`B&}�:u_TdM���x,���D*��=m��-
�Q��s�п�1�>c6b)��¢|���7k�Fu�n��PPPA�������8�sر���n[�lF�.��#�y�����о}w@H��x<X��2a�<�7U��w�BUU{�Su��'y�?�����XU���ZTV���F~~�Ĳ�~܎��v��.C}c��#�CU7u^h�@ �i����E���!���N�:����裏�a��if����H�N`^��k/���9�?�+FSS#�W���j?�֕�%��T�ՠ�S��p*���I
r�H"e۾f5x�>��Ux��M�1@Q~lZ�=4�_�g�w8�S�J���$�fӸ�n>��9Du��a�U��-���e�X�������'F�)X��;��s!8�H�uh�0�� #a@�-G����n�r��"��h�w�BKBCJ	 m)Pe'(��2��=�PTT��g���=�p$gq)�Z�p�.т���G�"���{L�6��|�]�~7�\ݵ�(
B�(���U�m�!�H�����1Gv�$ƍ���%X�q-.�������K`%3���k�uG=D���G��ŗ��?��/�0
�h
-�M�N�9dzC�+׮������0d�)l��t���Ω���
�SFCS#W������@CDd�h�|�ɻ�hʇ�d�&d�D2����]�ߟ{2�j�E�c!dST�y�e�Gr��_�5{È���sV�id*C�@[�e�"q����(<^���mEy�n$S1f2]S���n�۝\�%LU�J��D��~�����T��aL�6� ��sσ�t¡X��+�U���^���w�þ��ش�[�q�8�w�5R;���ѵkg�~��X�~-w7V�^���ϻ ��0$�_.[�x4���?������M�x�u�g2`�g�E��%2d�I��vcɗ����^:�
Ϊ'@޲edE�_��zC}3�D�c��>o���.Z�}�8��;������w�bݺuL,$�"-h��wB�������A� ��p�W`��7�uӷ8�S�����WUagE|E�H����v(���DD�(�ă���(!���~��&��})�m������?��+��d�*�XE4�y�Ɓ��4��x��⯜�6@?n��~Z6���É���r$C�#�=Kv��C(៕�ѭ�~��q�}�R6�0G���t��d��={��E��h�YvB��=�d<�3����vm�y�7m"����UԲ(�X4w"J��>� :tꊊ�J�u����{0����q���ݕ�����3qX�B�����/Aq;є
���(7�����أ�b��H�Y̙?�� �Ǭ� ]�������s����DnE�ܕ�G�b<��3mKU�J��Р@�G[ԋl�v�7���y�a��������h�TL]��B�^��x�    IDATXi�I��CH�C���G?�Kν�\|~�5,q�����d��'b�JZ+��e�bK]2�!;]"�)0�E��S�����<�]"��Q�j"��ڿ��FG��N�hh�
�p��T.�D�����S<�?�=,]�OB~A�k���u�Ep��nE��=�v㷘9g.{�s��8���P'NĞ=�pd�޸��K�j��ٵk������g�E"�Ƨ�-ƒe_�y6l�8+W��pb��}���ܹ3����4�?��ù�&���/�D�v����w1�~��)زe+�����:�0 S�L��)�Owޅ��������ɂO��p���a�3�~��bT�W�C��r�)%��Mع{7W�=�$�zޞ��۲�xw�{7J���g׬Z	=��I���i'Ayy%>�� -��`	A@���`!����^(�x��qA�r�M4l5�ۃU���ʨ��G��3�db�9S� ��/5�1��cNkc�O�_?�6@?.=�����b]C(^4}�8lۼO>�<����&ƴ�N��r`�1j�c=�C��FT��̂�WI�2��\�56ǡ�}l|bZY8��&h	�gڂہ��Z(Z�u��[�#��3G~���g�푹���o�	ULO<�(F�x����8�~��ڛ��]��5n{�����:i
?�u��nGtGײN��I�0` F<�4�/^�X:�EK�"��@������|��7�N�;���沤�_��F�%���;�\�䦨ȦӬ��6I���#��U^���L���vu}%&}�6|�-����;zp)N��%w�;n���r,� �}�x�<��q���@i�	8!��O��d�"�<�XW�������@"��:{���� C�y,��Y
ʣ�v�[��03M�����~�ݼ�+V����ǟz���7�⋐�s�ә�ODQ֭�=�x�>���ӭkwn�WT������i�a |��W1o�|*Ǝ��U��[Q�n���h!E�v����'_k�޽z�c�a��믿�������íwލ�+V���c#�#�҂��ӧOG�.]��o /� S�NŘ1o��}��U,�#	��'� �ۍY�f��0���f��7߄��]��aW��];y��ʫ�s��GG`��y��7w�\clܸw�uK2�|�t(i��!�;��bD,��B�ia	r�ֱk����� ��6D�a��M"���A�E���%{�S�����s�$
����ǝ��cw���Cl���{`��/�<?iΚ���ƍE*äI2�*���(�!���c�z!���@%�/�e2:��e�C�z����I9�Pe �Gn���3��A�r�hڷ�Ё����ܳ5��1�C(�-a��؅�{ʑ�_�m�u+��������n��o߇� ��Q��;t�����lS�jA�~=9֕��C)|�q|�d3"�$�/�	M�iy� �,_���*9}^�:�J;u����X�z5:u�Ν���f�d�=���D�P%���M��_�A�,Byuk�_z�I���X|�b#��<���a�i¡���΋��oׯ�;��d�r�u��m�@*�f�D�S�}),�|[�9 �=xnN,p-E�4�W%�&'>Rp�&2��i �6�BM�0�IH��Hἳ3��Hc�ƍ�펻0������PQU�L2�+.�=��s�u�z�[�G��������Wp��]�vx���t�R��޻l�K�/��#F<�;＋A����HW^5���Tկ_�����t�=3��=W�d�s�Wb�M�:'�{aI	x�q|��<��?3�1�Jb��s�i���cQSS�Hj���`��x�B@ݳ_�r��5k��Ӊ��<���g�y��AZ��#���E��/���=˜��3�cܘ�||�W�����PZZ�3�<�� >��	\7<� �:�b�a�s�;Ud�EOr�a�|�4���`Et�!�Qr Kא=",��A�?
��)�`�$��%COd�2�W����~w܏�擮��*�C��0m�a��.\�
y��r=���T2���<&�8�H���`�'�sdo�ݽ�I;Z"���D2���"xyp8\�֥��)��'PI"kDn��t���	E];r`K��}()(Dư��^�v��+�^���mdӏ��T�4��o�A]m5N8v ֮�3g��eW]��5�&�X���Zj�R(�!���u�f��atl��}�G�w'c��M&�z헨��7�TV��-?�����9g6w�;�D44��8��去
ǡ���z���&�%��Rk:��2˞4��L����$B)���!�X�ݍ�CFIng��u=� P@������&�S��8���m=}�B|4k>�5��r'�"]��;��T�qI�@B�lI��	���S�q�����IHj4������T�u��Rat(��������
w�y��x*�S���N��b��oYP�o/F?�4N?�t�]������s�q�J߱c��P�>~�[L�������k���ODQQ�|�	�\���<� W�D&�>u��]�{��7o����Y6F��#F �`��O���^�o�{yA�z�M�����ޚ��}���^��{2���'!?/+W��Kc�"Ob�С���+��i�@��ԟ�yޏ.����%��kY�G�O��d:�)ӧ�g�^x���x�n��8��3��Ïb�GS����"����C�t@��G�N4ɮ�H-
��A�^�Y ;��8`)'�I�y�y��?:�A���Z�!�U��=�挹��;o���T6i�a��m+Y]RYB6�?j�H�9d<��N��.�[b1-K�X����ťAm�t�&c�c:��y��v�^Bq��,D"%�ܹKÌ�#�����3g�BAI)���r��G�S�nx�ٗ�v���_8�S�8LlٰnՃH2��X#6}����~��[�+�l�ĩ���3�(ؿ{'�,Z���^8}^477"��zx䗴�Kc���/`9�������� �֐��v���A$�8��%xr\h	7C7$�"�Bp��uz�V7Ӳ�<�$�5ըؽ�h3�:�CSs�hوg,&�=|��X�t5ޞ��+"ɯȥ,IndN�2�466"�Aai��D6�S���y��*�G"p��#Y����Nsd�+{`�d���ePm�T��&��ʪr(2��8�]�{��[M�\��c,�j��k�x�~������ѣv���2��z�=V�l[�u�Vmբ���f�4������ۦ�|*�����Ȥ}I1v���#	�62�����uNN.��r���#�|�����.��Pp��*���ү���e[�4�e{Ա K��ȣ�ѩS�x���]�x�wtln��6�<}D�qvE�!�֡�p�����N�B����\ȝ^-�hI0��,��:� 0�h����ZiE.�^����۬_��</��C?t���is�x��O�Ꞡ��2�MR+ς7@s}R��J��C�,/�5���DŊ�A� ���s�h$�9��c�$�Z��F���v;!�"+�2��pI
tjZ��1��7+���u��k�6l޼�SȠеc'|��f�z��xu���n�TTVc͊��ض	{w��J]S#��a
&:�k�bqi	�	Sf}���yO�S�k��:i��ѹC)�L�������Ź�Ͽ����,�>h���%�=*Y�f�4���	�dooÊ��s�3�O�GqA�T���3�BS�̙8��v+Zj����m|J&�� ��}�AX����%����)]32T9~B�..��L�r��=���yk4��&�}�m(+�Q/����>��%�W��W�BT�$'t�;UD���<o/.�G,b6��)2P���L��7�S|>��$�iQI�Y�>�Q{�[�q)��A�����k#�t�;����[����i�iy��_�Mea��|}�)d���!7�յu�� �;��r�455q��Lg�q9��֊�E$�,J�ߧ}�{��MS��R��c6�!G:Y��M4�;*n7���jF���u cXv:ai4�Dx;�S�I�t�� �6�"��$��GRU^�q������Ŋ
�ERfZG��
���u��ԯ�)��y��Ց��!p�}����>^Tw�Lq��M��V]
��)�#��LRId�:��ө�t$v�"͌���tB�lKά`!ih�ȳ���aĚ��^خt�M��pkh��ux�l�%B�*�,��;�Ǟ�۰b���UV։�рϏ��:\~�0<��s�[U��P˿\�D�>��tKƎ];QS_K7�TT��RJ\�T0q�|�75cٗ��u_������]:wFm�>쯨Ď�{a�*.�G���4Ų��x�JXGNc�H��u �N�o��V���FڄBd62Gq8�NG�p%Κ�o�;��+~�^=��G�>�1o�W<���͊��v;"��A�Tu��sΦ&4K��J��D=�d�
c_}Lx#�[o���<
{�U��ݻ�Ų�vݭ� B	�.7���D�#8[���3i�����m�t�9�븺T$��q~d2���FQ�B�m�ʤJ����CUm�-c"��rWH�����
�'vk�*+, �&���������]���l*ɠl�B�Hd�̱����������,� ��Bc}��O�`;yhaT_[c�gт�ey���/)0%�y�a��\��t������A��9yy<n!6��pC�X_�6��Һ�K��M��/
@���
���r,C�ȼ�Z�;�	n�Ӗ"J�z�̢@͆_�ˍ�����c�W���+�����<7i����p���$CA*�CX�-$u$�q���d��+H�_�?Բ���8��I;aJ�U�)��Hߤi4���t�vꄌ��kz}� {g��j^�=ь9S?����Вh��ACsg��1�M��~���p�c�aOU-�ugN��_/@qa.|���
��l��p����ӏ?���3?^����0��o�S�B�5l�~���p4=��������%q�g��)�5�GƐ��E&/�oI�LP�����U9�$�p��L6�tڀ���9�u�
Y�6���9�0��G�\[��:A�cx�ч0}�,쫨�֭[q�M7"���x)"��lk"&��v�LxN�"��#O���A�t�*�ɬ�x����D<p�p��ivh��_-��g������ $7����ʐG;������YzE�D�#;_�����E��c��x\n$	���Nj��FU-$����)�kGill�5�B�GLA42��s�V�	��J'�$ ��?k���v)P�������ΕI]�I�����!+N��f������"o)�����M|hVo���G)��%_�T*�ҲN�3\(̿fVc%����Waw���h0��)xŋā�Gn ��iډI��:W�:D#M�dMǋ4��E�d9 X�ݡ�0�ţʐ�.)��}�G_��w<��� ���oN���YKVEe�7�'y��	-��"HE��
$q:�֥**���-8	
��I?D"�Q����l�SU�J�8@"�hC=,C@a���<
��Dj3�L��d�XD+��{ N!�`��%+Pz�Z�p�$X*�v��y��3�$.<�Tto��� �`a������Bx��x`��0� �@Yi��s;�̜�2PҩG�����:��r�^�G�T�3o1����HY�����yO�r���"�e�[��T>��Gɴ'��)�T\0�4�L�{�?�
�N�+��0߇�G�`��܅_�����YٍQ�Ά��犗S>��N���| BT�$�ǻN�W���T���ň���7Ǝ��x1s��8�ԓQؾ���p��C!���S˟4x��D6M I�.biQ{�"A�0M�����"R�tRLH���8t�h.O��T"�"I9�Ԅe�p{\�h���\���f�H�d��1@�̜�kj����R���$�`�^��������XR�(K(��e.��eX�ɏ�.2��X2�:���
���q�y[��F&-�9Je#9)h���fy�����������syJ�#���&�Ñً//���qu��h�D��h�����bX�3�J�Z�t��i���nȬ�$)�M�x�nI"��N֯�Wｩ��g��:�6@?.��Y�z=7u᪈��|�|�]���ܪ��H46@��F*D$d���" m}����F� 7��(>7���������� �<��p4���m	��+#�EQtb���m�jlٴG�p,��c�o�GFb�+�Т;��A��tI8��T(	LBii1�++���K$q�eC1≧
'�Ԝ�`=�ĵW_���}�ޭ#��0p�Qhi��9u�'ࣙ���-���+Eʒ�6d!3��,��A�HƎ��p��o;g��K��0�gj�+l�C���4bδ�x���I���}�%l\�y9�hIix𱑸��PMc��k ys`P������%��]��|�:�C�?���Z��Z׹�\�54q��q#��"@��v#�Q5K�]�I�G�Į/H"GU+���1�g�t����4i�	�,@"na[������4��I�bp����)��3�h�Z�d!,#� ^�	w�˄I��ߩ@6�O���%MTֶ�]Yd���(r�d��r�
`*N�9�[.��T��0�VU�`� ��h�@5^Wϭp���}Zڡ���yr��΅fZ(n��,�����a`v�p�Z����*��W��TڄC��{�g��(<�t!�^�_�@�Y�SE4�`�_���KH����E�s���;��� :e"�E_���/lg9��m�!{�'������Z�R}AJ#pH��\�s�RO�M3S��)jV�#[,��$*� ��\6��CVv:�L��zV�𓔨��+��v�^v*+;�3"J�xΆ(,��$B�voszUXze�A���+�Y�o�C4�k��Fi�vpy���JT�'Y*�L�������i�OČi�p���X�|�Yga�g�PY݀P8	����ѲiN+�z��8n`��a|�n5���8��m�&�9���#�W�� "3dG�H�]��C�T-���yܲI�s��fƲ.:�M�E�n@�t亹3�@W�*��"��x4������f@�@��>�~�~��	�) ���f��i�A A�+z1�+,X��\�Udf��� ������2m����rX&�9��<;&�{��ˆ�-mÒ��ʐ�x�w�,�ꔸǻI�b�Ds'-<��E�;�ch�_{�%E���U��=y��	U@0����zԃrT1a@E8b΂%(AE�zP1G2{:w�w�.<［�]}������XLUwծ��������g����q��cዔ�rEfJPB�|A�ٻ��F"����!�i|����3�?�W�t��8$�`�5�I`'��!�"ܪ�{p߃s��b�e�l
�$B��T�Tk+|4f���e���-t��J�Lw�gRI%�a�nh����/+c׳DC��A)/C^P�[�2'�W�&BȲ�&;F�d�wZ�Q�^"# �����IV6y!nz>�3f�
�5��Z6����9I��M$���'�U���O�B���������ޅ�}Ԥ�N�y�y���!�hA@$)Q��:�03�6#*�lO������L:Ӧ9A$Z�f�� �F�3���ߵ�[���1ä��
gg#"2����RK2@��H��YC~��CЧ{O�<�;���K��|�u7>��#+�l"��0%7�j�K���٭+ҙ{L����h��&�Ӡ0U�� ��d3IX�$j۔b`�^�jS��T
o���mߍhQ�hl�ꮂ�c�*9�y݋�f�5���� 1��N�`Ôu��%ƻ�B�$�)�i�nf.�N���@M�
�qF�o��k���E^�U���2dͣ���2�υ�Z�%�k:���E�yڇT娢����*�JLB��z�P��(Q;'a[�y	���ͣ���'��Ht9�SK��sԹ��N-~�ݩz�L�k+�������    IDAT�ű�:ֿ���%%_ D}��$ٚ�?�%���3���}H4lg��#G��t�F�p=�6s�ɥ,��:~jG2_ͺg�=�������B�e6�OhlB�9Q��dO�o|���6|�=��'�*�Y5���N�r�B�%Ο]Z��%\Q'��BHvı�JdH|�z_�
�T�w󀑄�g�����ȥ=Z"-�5���ϥ��)ȶ�Y����Sb�
\��6Ĥ�@�V+�
��}h�%�G�o�~�X+\��%���|,�z�׭O,�0�Bz*� I��-�I�A�f�s=�b��F�>h��gҳ����N4.�hӃ��cG�ݴ:9�]"���_�  �G�+����BC+����UuP(�dVG8�!��ٶQ|��Yt�} ���f�A�tXrd[�E���p�%:oF6Ê\�M�4����g�Q���]��Xy����[&���02��H$�$Й� )�d�K�=��%(Jp�j���>���%t��=�W���PL�pl��$vV.�������!wC2�����b��W���aJ1�R����n��R�D�+3�E�Z��?O�E��*�9+��]���.��iq�:%t��v���Q���6S�f�CSb�G.4/wJJ&wsh�@	��T ��T�8pB�b%]�ЉS�+͌@_�D;J��ĚU�p���%�]Y�k&Q�[�.<�����߃_��~�6����8󜋐ə(��ѫW����X�zsc=:�V��Tk
���V��ڍ?BԂ��g[�.'��G�SC$�"��2��n�.� _����h�+x�[�5% �6���~+��� Q�V6�#��S��pT$�EZ`�]f�;��`@U���f�ڰz�@A6��"QW�@@��wē98�ZI)�45�~��>+k<4�#N�����V��BB�??�,[�g��U���/;��Y�YE!?2��9�W�B�X[É��妠��%��u��W7a?XAwE�@Q}��2h۱�bVM��z�m��W#	�N�T�`[��
QS��D��{���儕MPU�BS]�Aհ�0��J��s����S���1�J:���f�2T�œ(.+��"�Ȧ[��M�jja�,a�0"a8>�+@j�Ӣ�t�)��fr%Nml�R��-υIy����Ʀ�ц%�</v\�Q��w-�4�ϠK�6����(�ػ=zu�f]w-ďۛ1���H�� v6�aI!�	��ʁH�@-s�O�V�A�q)�{�4��]��w�؎m�ƻ�Q�g�*[n��k�ӵ�kB�
�ꂪ¥���\�3?�1�6��]9�G�z�Խ��;�/�@���km���wu���%<�����;#Pq�Q#X+���������_�I7⋯?Cm�C!�
l[��_A}CNu/0~��;|����IX�t���<���|��ؔ���3�WE�$�; �w��/M���Ǒj�s���QTY)����M��{7�#�^�j�W���a��L�,��D^"��!*�Z��#�&�$�:-@\R۵�n��I�B2��T �Qe�i+��P e8x��uH.|%5h��Њ�̜3���=��ao�O��U*���30���o}t����h���������	矱�mYtU&�-
�ZJb��/����;�Ti�HGG�;l�b�[Z!Q��*H.����!�t�Bqm5���͐�y��$���JCH�P�:�\�A<�E&Q�浄\�uT��9!�Si�B~��;'�(j�	G��Ց۳��BqQ����`�t0T
�_�_�ֱ^�*m3�HXE4���a��h�0��S0-J�5m #L��j��۔��AK|g��󃜄KdJ�.	�P_��Dj���-C��.�p�'tB��_��@m��;0�;p�m7"���ѡ���@O41�o[}o��9N;����oA	�~>����	1NI�Z�4���FP،ސ���9%_��h#�6)��.��q�i��k���Ŀ斻@�a�{3t���/����KD{�7��I��S@#�����K��0��焾��%��F
'��<��	ӒX2��qcQ�/����d��Z�6U�x��y�Ǜ��g_`�1g0��kU*p��X5���P��?���۰	[w�ă3g�ť�`kJ@^Ta�yh��cc��m�3��#F���d
��Cah�0ϬEBKS3�%4�	1��$�꾼���&t�)�j�����+�K��3ivʙ"���e
���� �
�Ц�l�ke>�ӣ˺�=���xS�τP�����?�j]��>������D�e�N����G^�<�
�X�������/�pϳ/��?r�J"GH��]�f⻶�>�k�J��}���>//{���v���e[`�+��UT�u)�d2�'�.)=��w�D �c�+�P�l@Iq�����K� }����������㞻�DǪr�(mn�gpS�OE,��%+pϜ�Q�� �u#ф~];a�7aώ�h׶���gvq���),���Ԅ���o��9ФYO���J�޽����O�Hm����9��ոMO`#�,)�̦�dF�fa/،�*R��p2%ГJ�e0ʜ��-wZ𨂍����҂�q˵W�$(����߭R>��;wC����8d��Ǟ_�PQ��"+ҞEF�j��/�E?S����%d���x����m^�� n��_RK�{-J�&ϟ�,A�@q6�������i8���|�C0I��oB�{(�_��r�ZWʹР�H�ނղ���[6�y$29m�+0j�ܧ;2���M����;����i3om�G�l��Ƴ�m"���@�>������b>P��O?���|�<�k&N�{�l�[Z`)D������OÞ];1��aÇ0{�l��14v�%U�� �t��&u!�^_I�%w[w����JX�>S�=E�>E��Ȳ#
=Y�T����f��+23)pM �D���vEihmM��3�޹�?zb-\�����_9v��QwL�U#��]3��8v��!��']��~�x��Uf�{�=S��R>�Ğ�x��9i����������85�7�olM�ƺ�h��/��Iv�
�D�P\U�T"��ĭIlxg6�h�u��Z�x奊�
�RM����ٔײe�SB��{�X��7W�t'B�!����1�o/t�,�3f0G�+GA�B��$QJ���gJ��"��N�JH�<��s�>����_y-R��D0R9b]wj3��<����`tM��]���D��i�*C`�/j){�h��k�Bv��K���3�Č�o��'qh�0j�H�CMU�z��|�m�:�|�nI��ϿF���H�:!{�U=F��`.�{ �IB0l�AT&�+g:�6P[ݶ�>�R�l��)V��F�7���8�Nx���a����򬜖.I�R��VDo�	�'�BR�T�(���˝�:ԥf'8�� �V<�F=�y�t���!�ѳKG�Q,-bXh6���mQS���x#����܇aC�C�!��p'�g�.����>��i{��~+-]�O��닰���(��XO>��صeb�"���./�R&�B�1����ʊx�a:���ܖ��PD^�{��'�WYA��iZ�h^W�%j\S���OzG�=Y�<zwl�/�+�����_�����ߟ~����_2�ɷ�R��6f�z�G<W �fa��"PH���-n�k�f��d����-�����^);������ׯ][��w�
���g-��D`z�8y8>��UE��v}=�{}5N:���P6��VN��`���d
:y����N�7�Xdi�đ#G���3�?�8"�x���9,,S
`��w�����XT���^�!���_~?��En��bd��K�/��\ ��-2q�-����R(ARD#yU���	AN�r�"�8���Q��r��R
�E��Խr���[�i;�z�5����׻�C~�d�L��i�nڄcO:Z$���^w�ÿ�6��������̜��.�6濲�l؀@0��<	�M�����#�Z�I���&;ڞ��#�\���y" f�g��P4��=� 	ٸ2y�p�T�`��id^��O0�<��m��]XQб��A�(�0�&��#���}lt2���3�4�7!�\lٶ�|��~k-�-��᧟��pn�w�)A"ш�f�d4<�.I��C�U,mv�Ǭ����O`K�BʦI�Ur!�S�X��"�?/�`�ct�H��	�pI��8$c\G&��E2�~���~U�� O?"����.���x��4��;��"�]q=ږ.:}��KO<���~/i�SƜ=���:n��jw�t�C=z��TH�%��s�-$��9��?�����;���56jS����k=���O�[/���o��+kVo�ak��_|��kE?�� -d.��NChj��+�����;oB$�b���`�U��أO`���L�fyY	�v����u��Q'a�������=��z�ZƢ~�ƘSO�a}����㢿���>Z��=��MM�}�i_�kS�[�q2<��S�Je�t�R<0g6�r�����E�z�_Pվ�:oI ��CP4���%�T=�����?Z�{���HF�d�A��Dc��R�&T<���&��٧p��W!���Cz��K.�ꕯa��ñ��Uxe�J\>�*�?֮]�V�WL��C��C�]�iwMg��|VGiu[�?�2�v�t�.i0,2	r��M)�9O#��ѻ{G<��,��q�om�s��i8��1(�l������Sg��t�G��}���:w\5̟�F#��9�d.��%�|�5�ڭ\͏e�_���s�����0�Bl&by_�b���>\��@P#��,��O��hۦ-��4l�e%�W���ɮ-?ᓏ����M@�z�mSEv��?✳�b���[��ڷp��ix������͘>�v,[���r,هP��
�<&pm����r2WCa��;[��S��|>Ċ���YF��-	n�[>Z,�xb}P%�2��|���I��/h9ȷ���֧yx�5v.���}P�㮼�~��򫯾j{�=w�uک�t��.{��Æ�X����o($����/^�j�ԧ�sDIxt���-g1��˿���9k�����%����C�� ,�¤��XeT2�7�%�1����vұGaҕ��Ԃk���K&L�w_�}z#���[o��9s��Ư�WT��|	��ꃃ�˯���Z��t�N9���ƲE�a�a}Q�gν�Bl�ǧ��h�L�+����O9N6�����T�����5o�G�~��A\s�](n�����
%}��ڽd1���{�ĹV�R���ل�&�9J�4c�(��p�m̕���e��Ԇ��{k^�M����_~�e&��ڀP��T��R^H�?�"�t����7�������Ȓ�o���w�A8B�1���m�t�B8��x�@��E�`�Y[f�j��~;�x�U��qXFÏ���Mw܉X(��Ӧ!RR���7^w-F�s�}��b4�����Ÿ/��7^�����@�=p�%1宩�}�@y܉P#%�f	]��O�*�iٞ;Ѵ� ��]x1d��F+O�F��mצ=W�9Gg�[+g2=�\��>�#F��TIiG;�w�b���9�ջV��.��q����/������V�<b��){��$��A,�rǉ\��l�,���ˣeO���)-f~:�Z��a�f!i��E@(��O�M���5�Թ3BT7�Xf+�W�*��%���{��t�7]���;�ޡC���6X:��Ba��"PH�����x�������J���5=�pAȒ�7oo����������w�Z2rY@����ycQM9|"km�+/>���z��,��Ɯ�}zq����W2��ǥ\�t2�����'^�L�B��	��z=z������-3fC(n���X�{p���8���x����s�e���Ba|��wxe�j����5��'ӈ�S�ҥڵ��O[���L���'݀�N��u}H%�H�[�E��C��
�̐,*!ۙ&�I���Kr���HF����N0���E0��y�v,_�+�o܃l>�p4�`3B��x�/F(�܇Ɗ+���f��m�*+��c��c�A���q�M���o�f>�V�Y�+����Ȋ�����" ���2xx�t�{kҩf�}:.�p"���z��"�o�����C�ݰ���dR������&���8��ӱh�t��	�;�]z)�=��x3�9i42$L�|v\K�,��6dգ��0KH���^}GC�s%��yvqs�^(+�51��'Op����?��:�?o4��V>��Y�� ͫ�OpY>�$e�;����1k�#����d�qD��H�5���A�n��R�,�d�;-$sL�ѭN�c�WJԁH����њ�#�$Q�� SI����mZ*	3���J�1E���N�h�pP�n'?p��~�r�_lXw�'�ظ����֫��X��7������cE����X���l^^�b��O�0{�����է�f�r㉿��B3���o}tt���%�$K`�V������hƲyO����0h@\1�BTU� ��n�)g�����c�s/b�ĉ�r�\p�x�K*V�xj�}��2`f=��h)���p�)'�o�n���k����oi@��v�񗟱e�Vl޼�}>��c=|(+�QB'���}���O�#�=�K��NEW�� �y������l�ҧ�{�	�xI�8�W�,�J7#/�f�ϓ%�P'�4��b"$�*6J�1D�L'�1Ou��B29n�S���5��f�P ��&G�����,�H]�2�� [[�L�&�xf[���c�P��{�,�·�م�>�{�~I�%����^�s��W;l&����(<c?㴓9y���A��d+^���o��~C�A�^�+'!�ᬱ硺s��m�M?mf�>��u|!^p��mPI<�`�<+Մ%���SND��-�#au�v�. �ӓ%� ���*�&���e7�Jo� ����2���n��I_��a|~X���=�߀�V���4K�ʲ�����H������'ݚ`!�|� ¥Eܭ!�����I'�G��
Y��m$�^�K��P���!�� AW4R�ki��Iz��t�$��P�F��X�����8n�������-�}�~ç�v��!ѹ[ב�HM��}��q������󙿴l��iO̟~�i���ךּl��ߝ��M��ztыK�S�2�#.����i.o!ڮ
�`×Mb���0d�A,�zH�Y�=��󯿃����4jʪ���ʍ�G���~�ݛ���k��G�De�q����:ɓ6����CѶ4�Gg�D�>ݘ�^\Z�H��?��+&��d0�����۲�TVU�_6�i�q�WC�9&=�IW�=�R�7	�ҧ���5���#uO��@$�&QB �⇾�Ȱ	3�z�aM���!*G(����C�d��N�CR5��%?zj�S���$dR)C~�?��ap2!:-
�}��Ln^$��W=3�G@�1PLvl�Wz�@�9��L=����op��#q���`���J��@R�M8��c����CR�\��w�������qPo����*8X��eth�]��@I۶���l|�e+�Ί��]@f��4�܅|�l�D3^|�1�9��e**+��(���T--T6�ڊ��r^�I��֦:;�H|��hnjEuU%;���Y�R�[q��֦������:�me���;��y��eI���cH0�D����'	�4s�IŐ� .y���@��8x��RYD���Y���(��?
ˑ`�
w���'S��=��ɭ���H�&N+ڗE���+�u��-����w;Ʒl�-Y���^}�9���BB����sWH����Og���o����N=c�un�b�С�����`�9�����V�eks+�d��:L�AQ�j8���U/=�^�:�$ !���%�,��R褚�h��L=�6�U����0���Ɖǝ���շ߃��}x�H��J����NAPs���O���K ��4'�̥`�IF3~g%�  UIDAT�ri��#������]�x��U��p&����Ma�s�ٜ��,��E�w��r�N�kh��TE����6� ����(hI�>�@5e�ihA��i�����M�Fz�^�O	�	�}�e��g$���ӆ�!4�����c�-j�࿩�6�<$�+z����x6����|lUJ����$Z���;2�C~�T�eQ�B%=w3'C�������k�k�Ke�ڵU��	ybP?Õ�ͥY������%Q��*a��@|4@w�p�̬�`$���BIiR�,R-�(�kAB2K`D���F �����P[�D����,K-�E�ؾ�	Z�,�J����!�[,��*@sE��H D>�
��V�W�t����J���0����u��u�4(� b�$$�B$�u�D�^Mup�i�,��V���$:W�6_s���ǜ|���{�e˖�;�֮�x`�l�^�GW�*��k���F������n��|������3��n2�#�O:��s�������U7�������lț�HL�E��ðl�նc+K1�ǫ��DkC#��E~��"�06}�5&�1��3Ix��oB��ʉ�����p��greuǔ{�x�
���P8��=?�4������CrLO�(�%Ռ~޶cWMG�'O�� �L�g��M�uɼ�Q���3k�_S�&�RAT��E�.D�"�ɩ��|�)a�+�J֕pP� ��"eIU����O1�;
c{S��Y$JcA����r���3����њ�@��^�`DO��2�,8�(+�V4�4~��? k��EYFK:	Q�`�*���hH�&�Ee,P#)��REKjw
� d�\��W��'��A(������"�l
>Mb _��� �vo�� 4�A7�Ƒ�&!�ʛ ����^sNu<�y�q<���3z"��W��W	��C�i�c���|��ⲿ���q��w��]5ο�4�7��/���Ϳ����0��z��i3���_��_�9܇��jp��q��I8�����q�M7A��<C�$��c�Z�<�w<�����"D~��,��jE��sN� O@O�
*�	Q�MRXS�S�gCK���&!�XW�AR��\���+�n5��^v�����ݦ*7n�iӦŽ�u�޾s�S˂e��w�pܟ7����w�|�K_[u������ǡcU�{Ǟ|���n�����X���u�Ei�@��S�H%���ԅ�>0I�łF/�4JB�V�+�P@c	OYSoMB�m��Q��U��m����ߜ��O�i���D��-��e���75�q��1�⊶�2j�i�	$SiFKS�rlv�"K̼nrH���Y,�!s��\&�~�?���6� 6v@���9��$t��²������;�#"��Z<;�>N�?�o��)�8j8&]yn��*L�r+��q���/�g�s�8�B�;�R4gnU���M�9�N����9��6��t3���>I���`Μq�y��+'�s�>����<� R�yWA��|����G4-a��8!��.hqC] �G����N�/��N�j�ﹷ�IE$
=�E�߸�ݺtF��}��g����W"���k�v��=�T�rұ�����s�̝������O7~������;/-^���#G��Ï<�c��cǲ����-[�A�T�m����A�~��x�gx<p���;�A�����CM��hߩ#N;��K�@�JS6�!�;B�SW�: �y1�?sF.�d]e	�p�1�~������5|�(�(�0��ȄG/2�o�Fށ�M#�N�����0��8��*��^������K��v\���)u{v�ֽ{��C��7,#�¶�E����������|j��v���k���+/ׯ�_��{.���/_�ї�=��?�bE3_0��j4/&���v��If I2����q��a�r����z���s�Ű��t�0�������[UQѦ=���syz�76֣��E!Q���©'����
��[n����~{�Y�0�����9�N*f�'tV��hNmp�Enj�
G��R�k+J�l��)��5Ѣ"L�\K�b~4��	�\=����\�7�E]PU[�ję'һ�ɆOp�q�e7����S�GD�@���g���'����=�l��,�:���q��`S�����k�'Zx���c�-���f��'��ϡ�]{<���X0o>����}�F��a��v]{�Ǟ�.�)u�i�{f*�G�m�ǻ'KJ�a��|ީ���r���%�������~��hmA,������m��w߰�}8�`�3p����Wa����C6��$I�3>�K�,��g��iӦᤓN�q��m۶a��i8p ����q<���[���	=��KJp�\�;P�.U����b'(�T�=b1jS[J�X�)5��ڤ(��{�VI���jQ3�����������9������}��\7����f��>��(���b0�V�ϜGl��u��������+w�u�(s��m8t��s��A�ٟ}U�β;����ci�U��*4gì T��kp S�-�5�ϋ@��ɧ����(˓G�A���-63���y�p�B��X��Ug�����`{�~�$���+��_c�=o�I�Y�HZ�����]����C��K�^�������j˽���m-ErU����6��E2��O�͚T!�!�7_R��$�(�흗z��bkZ����*v�ԲRW�P.��H��E�c�VJ7��
�k&�U�D՝�\B�g`K�o����F�;����B9�m�wYFrǰ�ӏ~Jw�ӐV�%�û��;G=��)�*m�����eZ��L�Q����A�T��eN��d��p,��LUK��2����#p$&�]BH����73݅��#�{���h�a[�`�
u��d��	/jpه��%A�:�S5���q?0C[(<~�򥠋���=��;fcl�*a	ȟ�$e�B�ۨ.���c��ã�p �}���+ &��.��z:���������i����ŋ.��/C�8v��q�N�EX���ˤ�gƌF�o9�g��8�?3����Wo {��������SM��u�|���Q�Wq�71�b�@���h�aDb�S�h�h���V�~01�l�p����f�����s�ݞ��S伶����}���{��2���%J�!�����xQ�ӯ��&�Ei�256Ł6���Y�Zӛ����;��m�)d�����7,�y�n����F�+؀>�1��<�F=��*m>�kU�hr8i�Jd��T>!Ӧ?�a�������e|Jx�8w�_a�{I9��ف�l��dQG���Yz5���:��9#�x�Q�Tɺ�H�frp�͛m���|��ވ
^�&�?:�ӄ�}
^ff���
�Ig��V��T@dlh8�����e�z�=��^F�m�{/ǚ��^77k�nGm����\^�픸��a�[�D�:��+�$b���dx���J����*��HŖ+���s������¯�������Зw�ȁM�I�\�,4�)�S ��f�3�g^�p�� ��f�r�V����_�|��5blb�ЭB#X���k��qH�ݹ���I�ZC��D��,oR�M�����?�S��f�\]�v,@�+n�^z�[H}�=J���^/�S6�?�I��猽jTw�X�r�:�@v�������E�&��t�ʵt�ra"L�V�"�T&�݌`6��	�@���F��Au��y���g����3�u�\F�ܫHP�0A*ZEi�Nӏ1�4j}��A�F����|(�J,`��Z"d���R/����e�����̧2�Xq�a���1��zk��ͧ~[�n}�����K�����u\��� ��O�V�>���2;=��j�7�`y��|N�Q:IB.��E�12f��ӷ�ID[[P�ihd[!��5��d�Jz�p�y��q�5R�(<"݁S�&���8�]{k�qu��ھ�ra��z�~��I��umT�7L�Z��"�j����Dl{ӕ���>BY�
����O p��_M7�a���!ёiqf̴�����&�y�^��bLywDB��� �����5�.��ktx=;�z�@���h����.(�Tu<���Z�9)�Ԇ��	X¶J^��잲xt L,�?����H��nA%5�&�ʘ�œ)��N���A-����ڲ^�i��ե����gOr��k<Җ�	�G�IW���%Y�_f�C>� �xBU��g�a��i����٩lܗ�	��������X�����d��[��+�T�25]���I�B���	��k'�����}�2��b��C/O�}���؄\��J��~
y4U�n͞&�z1P+4����a��Fޢ�4s�[��s� �B#r�M�r-u���S��/G�<��R���V���A����*��p��ް����KW�|����h� 99u����49��_�Dkc�_I���;P�R��~zG�����eO�.�Sx�n>��Y�N*�+}�+Aޝ��=��A�˧l�2����|�Grjh��w&�����w�g	�����zd����Bɺ��!bf��fP���v!�O$�@�Fƚ'���o��I�R���d]�Ck���g`�t�D[�I�6���@=�sT�c�jk���&=�:mlh�������o�j�I�8f?�������HُV��]���KP��i�h&��� �@��T�F�����Զ4h���Ң�����.��b�����hg���n`7�h���/�/�v�)�*������F]�g��c�K|��G��|���>^B�A�mf�C�ϋ�,��0^r1����;3Ԯ'�K��O�0]�#��7!]S�~�p �>U,�uu�4����1�Wv�";H�K'�!��{FK��C�vG�E�G�;U��\�]���`�~����ù'�"�w�1J��U�	l��h!��D�ĄB�"��p���'{ �f�ũ�EokqD���
Xs.`�"���P�hl��.��F�g��"��[��t/8��ߟr;�%p�θ~>�<�5߮y�oug|q&����Rk8>;��چ�ϛ^�$�V=���w��- Ǫ"����.�ؖʌ�p�>����]0v��D���ĥ��D/����{�S�w����!���1�@N���ף��9f�b�>5q�
ǂ}%r��a��U�:�h`�8Bf{�k���f �z�+ygI�J!v[͗��t�lL�Tc�>�U�o��7�W$�;��?��>\��5�&t�^��z��k�qW@��ѡ���"���O�)܀E:ѓ��1�V���8,N��`�6{�X�[�O��7;�p��Z���^�U�@��j�6s���e�Ȇ�!�_8==�������Z�oW��|���m����rI����� f�fE ~��>ڍ�&�w���4�,��������4I�o;������J�W�ds������%$�����8BTΏ�ha? ��*��Z��S�,�[�լ^.��Q�&A|�����@�0+��FbY��m���<^鬇E��S���` �=���r�I�
TLt��7�tX�6#)@�J��H���^#_��rl=P�*_���E�{��r�x����>a*Ty ����y=��O�O\������*�T��J�L<p:�^&���4���(y:��LmM3�J(�{j�bm�2�T���A�-\K%,8"y1���ITGM�	��v�[��v�ːK���W :�|Sr5��'����e��[�h(b@�5@�q�iLPm]����D$�U�'���*�Lw��^�d�RK�'�Jv��dD����j�*>���G��h@0�[73�-��0~�T�)Y�h��$��up�۩S)��R:���%Iu�wq�G_-�@�K��d��pH+% $�
����h׹?��?�eJA�����0���bYs�\�l��M�{k*����ߍb6L �{��wd�=l�*7C����漱��/O3�E,����(ɯ-��ŕ&�-V��6��!h4���7V�����<�
?���JF��*T(M���1 '}�>Б�����0�0ᔑH�PZ��I�	��106�Q�`>L��83�B�˛�,1���N%�3�[��H���@��M�Ԥ��Z_�qPD�ۅ?�X�@*�]�\9��y(JO�t"��L��k�d�L�<���/��4�\덿�	~3.ٺ�g���AdM�3I�&�.J�p:VG�F����(0N�0>@��lU�H�ƽ�b�}��vJ�&O��~]]��G|\�`���;4� ��|ƤjZ���"�JB�Ty�VA���ޜ�)�Jg��%Vn���o+\����u\-4�`�pgȋ�퓏�,1�
�Ĭ���!_��4�%g�����V�N�y~bP�ç�����+�GF}{��&)��b�����ns��p pΛ�7������#�]�T�x��;/�e����|�KH��U��9����R�a�)t���s��O�7��B�y���(>g ']W������ɫ��w��a��5B{���cQ�E�nx(d �9��9W�5k�h���57���y� �SR�m�3��X�E���t�sV�j��r�(:�*`z�_Vw��a$mb5�]������W )���?Ԕg�wj0�ܯy���Zi���O��6���S�/ίp�W&�w��<h��֯<��Y;+����ۍ�+���]�S`�䱵�����e�b.E����,:i�Ub�J�_|m�Z1,ۓ��p�qm�tn*Apb�o8����0�7�Zb.[#T��<A�����aû1t]�E���l'�"X{AA�
=�lx�G�j��c�	�{vA<ζ�Yoj`��Po����+rsR.����%�bSjs�M��.u��q���۴�����+#���a&.�W�(��ץ]!Wb�c�T��b�V�;���dND+��h��V@�=M�2	��M���n�R��/������/����P���pOW������y�{q7؇���q��]��;Gb//�����%s�\Ht+��ō�	�U�R~�PK   Ŧ�X�i�R�I �I /   images/5472dc22-a170-4182-a291-403007edeea8.png 5@ʿ�PNG

   IHDR  �  ^   sQ�   sRGB ���    IDATx^��]�u%��?Wկ�P�D"�3$J�ܒ,�d�e�n��vK�����Kv�r[NK����%y[�$�J�2sI�ȁ�(T�U?������`�g��v�����"?������ܳ��'\��^���k3���6���k3��~�?�'�y�$I � nb I����D)�����{m^��3�$TI*���[���p5���8���S�*�3����g�����\}��zJ)�����/��ٽ9Qr�$I̫���\�YPM �Y���ɞ�?�^��y^Y��o`���?�����Z�W-�'Ib=�����Kkm#W�"�DYFdY
!�a%�z^�C�Q0�C��1cS�A)�"�A,�$I'*H��]�+���.-����ڢ�f�+��r�l�4{C)���K� v�
�"k��]�);�'�et;}K��
� 1��5�(_��U� ��7b�M��U���<��+ާT.�����k�P�W���qv���v���;�O �i���T���Jlۆ�����[�ִ�$�-�x�Q�w3I�H����G)#�f�ϘV�Dqdr�q"3�u�P)��9bK���u��c�ʵ��PP����}+nV !�{~.I��q�K��Jg���2\�l7v�-31�wVjK�a�*���Q��M$����{�̕m��e�R�}ˈle�Fd���ŃcF�%c�Z�s�����99�H�����$񽁲3�(h���a(U)�=e�q�j�T���O�Q�b�2���������\�� �`&HL�N�84ݜ�m����r��xx��C� Il�zs<�g�Ʀ�$ʵ�0�c�qel,q�$�} �:����ǆ��R>�>+�� ^$*6c�1#Ӷ�$
�~���Pŉ��0c7��9f^#�|V�|E���]ʴ�����r��ʱ�/@dF��Ï��a�~W�7o�2/�e'ʌbγe9��{�l�08�IĹ��xs_�s�P�C���F��>���5�9�@��4��6,ʹ��ʽ�߷��g���q�$g��f� �l��+���<�C �s}�E�A�I�8.��*xQ�Dv���<�R*ŽA߰m3)�*�l��R����`����D�3�(��2�$N�$6��B���x��`�F��5��3I��gq����be*+v�2e�MeĥJ)�9�P!{�A��$ʰl$�L�4�DI#��A�3B����p�$�8�|&I#��B�^�e�b�4��9lK�V�6���Z�b���wz�\9�3e��T�q=��r�ML�D^`�*V��K"?��f�H��B�2)ӊ�
��%H">'Ts�q�M�(V��\�T&��¢��zA�q��J9,��,�e��k:��(H~�q���\T(���nmi<7t��ؾ����W%�S������G�����sB�#*�� �Tg�*6,q�z�kY��V�^�s̤�lƑ׍L�Xr�R�鈃~F���4��4�p�-ǽn�,��{N�g�g�v��֖jP�;��T+hk8��Z���f�lvz�aRQGV�����X�hԓ��P�T$�a;I��)ߏ�Pu�7Le�Ib�\�
�)e�|>G�z�N#1�8%��ȗ�Fo��T*���n��P�j���T0�C�"_�l�J���PɄ���(�m)�F����/l�H"��W�J�Ȁ�$	�ǆ	SEql�q$� 
�$g�	7����m�����2`h\3ް�?�T��n�o$�Q�T�y^���h������v۲m+	�Q%��(�1�<W�q�(���#��0l�U�c$��q�QS���KhB�1��X��5��v�8��{Q>_�<�C����B�hz�Qä7�(�`�P�����B���m�r�R������M��X��e3���)Ħiҽ3�8E��4D����0*_([�8"$$Q�R����
����˪8�	��LLZV4
�Ģ�(
)(\�$�υ��@U��S���� �冖e
��h�A�5Olۡ�&�B�۶��a#�$��qNT$����wΪ�/�0�4�{~�\�8D�EN�DGA%�J��P"Eȉ���B\/B�xi���n�+j �M�˖UF�����$�^��Ee��Q���J�����ȵ�(�7��k��f��A?H�=�vs.(L��C�RyQ�KŸ�j�q]b����Te��N���I���c�d��b�ʥ$�T����'!�+>'S��Ib��Ǹ?�4��\A%���	uRG����0ʊ�gN6��$��DV�q��0��(4�D���������7���8�L�4��v[ٮ���`���q3�W�</���r����m�=&''U�\�;ݮ��u�n�k��Eʕ2���$��8r,��Ca�}��}_Y�ͧ0FGG~���"��Sl�0�a�f���P��D ]+?���/Z@F���AE��$�m'�^'1L3�L�;D�<	��B���&��Z���H!TTUq��Dsn��܏��;��{65���\v�����}�o������?v��һ�~8��x�v��yt���Pt��N��2z�:r���k��t�R�{mLO��"�R.Ppم~2P�&��ǡŭ��aF��t����(�"
B�nvL
f�P�mێ)�	b�zӥ��91>�9w�v�9h�
/� �T�:w:#�X!7Jj,Ϗ�-Vnm���
�����(Qp��۬��#��;��(0B���2�t��HLz1�laj�4�.����'�ҳ�7,77,��A�c��Ub�U�
���þJ4�m�� 3Fd D^�T��0��'q���*��������$�/��&  1U�aXP�������)�K��a9vL��v��Y��LӔ�E��A��[P�0��f%J�ĴĲ89;1�*Ra�1�^�y/�8�����X@3�'�2o�� *�b�(*���)�2�Ģ'nt[���Y����08^�4m�`Gyi�Z�����h8�\1��*�|6E0OJ��!�#s�L����P1א/ޣ���u�8�cE����1e�k�g�.�f0��-#�I#�n�m�du?��l�b�p���ٶ���|4L��U.���ͦ1R��U��4]�I���:M����	�� �0y-�8��x��X��tU�;H�8�M�]U9SY|�9I[�;��A�H>�g��S�@޴�A��6��Bz�9'�C�ވ��B�-���@��:�*�[7���9����Q(T�f�e
���i��J1�U/��&���sM��v��\�b���@��6]7OyQ��^��]��pn)�_�H�Y��L�a�9������wYLˆ��"o�&e��4��T63�̬ꎑr9�E�^�Q�)�R�����*	����<1���Β���^��m�QKKK��b�~������!��L�x���u�L�e^h{sׯ_/c[^��3r����?�������ʪ��$��|ޥxƦI�!L��.~:�F�R	-S��j�|.j��vy�����e��2�LXF�u�C�I�������{����5p�U臓�y���|�B��r���v�pLy� ����u�p� �k�N�����-\�5�c�u�n�;+0������T#`[����5X\\§>��e}zT�7)=~V6L��9
���D���7b��Xi�!B�ޠ��c�2$^@���pu�·{��	KC0M�nA��i.���\.S�#LBq?N�
0~���Dh	�T��D��`���(���?K���@M� q샌�eF�n��Y�"`RA\$�"�� �c��;L0�/ g�t���Q[�k���ăֈ) � �qe�x��+�P*V0�z��H�c��䳥�=�OUJ~',���u�2>*ΓI&��g"�]HVd
O�0	a8HyT��]��J������#��4T��Ғ<���T2��9�\���h`ݺu�t�J��\S��(��c ^U��afыKr���I�+���h51;;�f�����t�%��V���@&$_��@Qp �����7��g�t���/�����q��1v�YyI�5�s���@�K��s]�=%l��y��^��x�y�H��O����*e[2�NyXu�5��'iؓ���9��؋�B����g�yv+�K�t�WJ����rn�,���z�c��jX�v-����a||ǎC�Z��z�9���G0#�qD��E���ز�E��H0p�=�@4��p���\aJ,1�d���6��D�x�!��|9[�(�C�c�T*��z��1����4�(�����.�}�ޓ����:��df,Ӕq���Q$�U��@�Pޗz��(���H=o z�P�c>�Ȣf'������enŰ� J �C���
Z'Ҩ�m4�1V�5G���̗�+��!$Q%'J�h��]7o����Ի?�G)���S�^u��r#��G��'V�G~x�i�&:+����ț
q�IC^֒�mІ�oa����܉���r�x8"t�NW�M�� �SSS��g?�5k�`rrJ����5���!$��
7�"��S6���f֭=����T$a�ju�v�M���z0�f֬�Ï|_�֓p��0��<l'�7�(�X&��l,w���3,�Vo�^�� ��]4mG �6Q4eQ��I��0 -R�!8+�xmro(�
����F��(3>�j�h�<�{"���(�����X7>	R�Ξ��P�.bl��n��������B,�������`ڴ��䨸,� >n|�,���熊�J��v�Q���%Q0�\�"��=�n�+ �mА��A�/G��L=��9�Tf\�^�#F���(kn�N���Q��5��U66�Pm7?K��|R��P��+W)`*N�'�)�2g᪲��y]�(ށ��-W���MNN��b���C{~�2�*C�@�r�U�34@�{T�a���|Q�|.�|/��Q���ƴ��j�3e�����\�3�[�6	bR���c]�d�;4�Oꁃ�J1\ȴ�i��2�N��Z�ky�z���=a�\Y4��y<p�\<ss�c�]���&���y'�"�}F���&�ͺ�7י�������=�F����w
��������r�;�+�IB���|&ej4�ǫl��^��v����yO�,�.�(��62ഇ�3�m���́�S�ȴ5�l\g�Y�c>_\5Zā���|����)����ؠNku�L���ع���İ�M��"4&�S2ݐL�9�e��ԛ�����s��H�^'�	F��]���8������z�a!T
�<,�cr��|ҩ��7������߾��-J�M�O�z������g}�O7�Zjy�ё���8w�0Z����[��ڍ����i�1=��%^�n��2&Ǉp��1w�<�A�D�P[���L�R���X ���`p��(�N��k��F0P ]���EI��TJ6��y��-TF���
y���Ba��Ǥ������3<��ؼ�f4=�7l؀��)ahM�
�`r��;����E�Ac���r���O�F��:�>s�?��S}��M�{]%Da;���%f�p�έؽm#�N����I�^��B����S������a���SSh�,��'�@%o�6	�6nB���>O扔�� J@%Aϖ�ึ�9 �.�����r�
��{B��J�ʘ������D���J@���U@�:� �Ա�� u�M+"qT|T���rΞ=+��,�� -���*:**o�w>W���xm���Ξ='�@OwaaA��{Q�SΨ(y]��b��zn��O-c�x]*l&�6�-����X���{Fd���[�Q�S�N�(���1�p�8f˲�@ �Ԗ��/��Q�T(��,ǻ��ё1*4�8^�=c\������ɮKy!`� �jP�zj�K�.A�U�z�ɸ�hh�V��,���8��!���1�{0#�4�ȫ o�w+��?A��X����z���X�705=�f�	�g�1`���2�y(�*�3�O�c��賹�#����'3����F�X4�.����a �ɜ��6���^Ȼ�:�@��+C��{��p=��vl�L&�Z&��C�X�CC���y	����<��.
���/��flT�G133#{/��3�teeE��Gc����"?t����8u���3q8Rv��A֧T*���O�8�7�]~V؄4���gr%a�Y5��kfF&��t��i8n�R�	7�OM�z��C���1�|,7�����P`F��L�M�U��S��|�Co|��O�LL��Sy�:@�_Kf�ϯ}総���0ܲ�s�g�����_�nۉ\t�mnݾ������+��=�ܱ��"��+�H���@D��Mμ/ҢJӁ��Kڨ�a�g ����q���:��M��mM�������V>��" �a|b
�KLL��G~����/>��^���)�:y=��P�_��p������sX\\Ď�������7����Yl�ua��<�|�E/���J�0���C(x���
�j�����eL�U��:@�Z-�޻ož�oÚ�2J6��!��D�@I&��(tB����x�E8r��@�Bl�f�/�#W�<ZD� Ցx� �@�Ey�VC�n��طo�=*	7-�xiiy�[��2Kc�(K�5�C�Q���k�}�6?~��(�v�)k�y¼�� �M��|Q�b�u���+���m���l�Ļ�΂md�e��	O�9w�(�;w�8����3�񊗬=t��z����܇�[;�FL^#�%�@�5�G��0�wQĮ���	�4�<��)�����M�B�� xX���3��y/Xd�8�4P����'�ŋѬ7`�#��>׉ʚ�q��)	�8��@�g�����82>h4����w���	h\2%���CehF�Z����ή� Fl��sS�F��Hwz}1��|�����1�=t��p�ޝ8q�i�9�"Ɔ�0��sb�ƣ�7��e�n��?��={d�(G�e��4
	��Iݕih�-ejD��33k��Oh��|O�H�b�* ̂�iP����U�ݰ����[����|������$����8�|1��@��#�aff�>�8�c#:�g�أ<1�������K"�H��M�"�Ө�gVJ��=�9HW��2V�c�䄟#��z|q.*����H�_���Y�;~�����1�I2�����gN��2��2�A&��<�B�E��ը��Y(򝽷�x��9���{���y�QD�c�W��&�|���~��R�m��p.B\>yEx��>�7ݵ���`a�����Cl6B����XZ�������Ҹ��_J�R@��N����+�)eI+��(� R֤�$��83��x
���>IDP�b�ݒ�>R��_#�O�џb�ف��clj
##��w�=�z=l\?�r���?�u;y
c��hu�����������c�(�Q�T�/��H@'�F���ۘ����,3![ׯ�;��Fl�<��3�($��L����ʲ�F����g_<�ǟ|Z<��R��<�ߏJ���n�w�m5e.�0@�����X�����'Fq���q��>C��@���f��Y���d������b��׉Q ��m�4[uy��S(w��5�2�N�A�_�~=v�ލ'N��BE�<��b+��K!<}v�#@D�ea�2֭[�]�v�ĉS2f~�ʃT#�ޛ
Ŷɳ�ʅBN���ebrg7��B�v:4t��>�W�N�c�F{��F=��!9;�[�máC�@���~���A�y��s	�ĉ0��,�j�u��ĥ�s릧�%&������>@�$S�d�(��K�/��ޏ�N4��wm�sy��`B_B�A4�FǪ2_�fC�a�;-�<׃ J���1[�uyxD����Ÿe����(��c�4��b��陵X$�d�Z+�Ӄ�DX3Z����p���8q�y��Fb�Ҽ�B:a~���Dp���T4�p��7�39rD�����J@'�+�wz��gM���P'ݼ�a��y���v8,-_��ҫN9%�E��˺
P&�0~�7o�`jfVVj���%n~�K�������    IDAT��$%,����v����5x��'P���&�7����"����3hS�,��{��l��֬ŉS'eOQ6���iA�Ua�����/!�(<������Oabr.ΡX�a~��֪^H��t���rM����ܗ\�8R"#�VO��H�,��&jK��l��U�����KsX�q�FG�f�L~�ֽ��������QJ[���׫���������W���	�<F�8q�������x����[7��Fހ�	*�<ry�<��..\8+�7i�+�n"
�}H��N� θe� '�u�d
�d�	��IQ�C<�4�a��N�*�{�I��Wo`^+��Ή���'���֬_���*|�MZ1RQG1����T��������8w�"n��n�t�Xn��W_�^�˽X�o*xteI���(K,
<�~�8&FKPa���T���/߉�ދ�|Z�-���Pt�<���a1ʂDl��	��<�/}�a��u�X'�D)��7��jb�� 
O6h�n:e�IqJbXPFǫ���}8r�P�d9z��x#�|T�Y\=ۼ��,�ZYnڴ7޸[ ,��.�� ��w����\���H�͖-[p��7��CW���nW�T����H��x�!����I��X����
�=�=t��@�Q�����4%�2���(��[6bv�,��Q=z��4뢈)�un(�"'80����7�q��s���x��$.\�$�9b
c�\g��`�刲�<�n'��t-^:�_�[���T����I^�N�(u>3���߶m�$�E����=-��������d�t���$IK1�6mڀ��*�W���9&�Q�4I���%����b��߸e&�f���C��`�֭��h�6��+5���p�m�A<X���/`��Y0�c��|��ljΡ0{�`�0{�� y����� �_+&M,%bB?/��B���( ����`�/���D�₀, ��ߌi�e-6n�(2M������9Yw�C(R
'N�ևYH�L�$��v�7o��=�\���� ˋ+b_��+m���g�I<^ظy�lڌ�/[��/2`�Isl�}%ɥ�6��z �u�����أO�::�N�'@��+/���P�]W������e>$I3��=R�OO��ɓ'Q�۸q�N��P[�ƥ��a�wa�7�s_y��p��ض�\z�����_�����b��/��/���ݣ�d��~�r���@:���!�����������o�F����-͋'Ie595*� �w�:���%���
IQeJ�ԭ��K2� _���LL.A�B�Y����D���J+��Z���P��9�u����n_gs
{�?`���(<��o�@��}����ַ�5�n�p����&����훸���{�#ܵ�xϏ��u�ۏ���=�mĥq�XkE�4+0���С Z�����J��/�h�x��>���w��.���bv;�8ƒ�Q'`]j�zT�$��A�J�Ծ�n�ǳ�=����8s�x�:�&:��;�,-J�����t�ĵ�r^�axt��s/�9�~�y	�e� �=�U@�D��ɽ�(��n�	��S9�����Щ0d#��S�wk��
p�Νؿ���$1*�̻�R��ێJɐd.=Om�q�رC�3�;�s�G����c���Z� �K�iʳУ!3��"yʟd�&�ȵ1����NMO��FƂ���Q�Ϝ9���O�F}Qܦ��t�=F��7� ��O=�533��z� K��JNA$����G(�|^��w_��7๧��1z�Y�6�/͡�1W@'=e��H�!R��}}y�����x��ؼ��ʾ#�1}MkK2����R�r��0[�n�cS3x��02:��5���B��b*L���43��;7���
����`��˗.#fވ�d���! ���µf>��}Lϒ θr�#��uX1|%�F�럅]�dA^~�e�����ZmE�[t�l�CĽO����5�w������SO�:6���y�.�K1*�`�X���/�v��~�Nlݺ�?��j&:u
C-�C�H|*�(�:�t���^��^zi5�ι��=��դY)m��2�]����Lcѳ'{F�W+x��Uc2M��[���$��wWw�qy�4�4�P�(r��P)�K'�4bT�9	v�	{t=w�� ��A|��Ϣ�`��-شe#�.]<�{������_�c�^u��R=Y��?���½^�`j�>�������� ^�(�J����cya��fӄ�gϼ����jy�v6�z���g(�,��ă3-�|]�aIl�+V�M&qIbkGi�2A�Yĺ��J�XS�h��=M1R)�$�D�?Ų~�#����a\��1H���Y#Id^����r+Ν9�/�̮߄���/��?������3�7p���K"�n}Ø�4Z�,7��������~Ղ�T��o}��f����]J��E�#�4(I>v~��
��X�DA��h�s�y|�k_��Y^\�J���"��֪ř�)d�lʡ
q��pw�u�=,^_a*�v��
�w3�D���ꘔ��o��FQ���No���s4v��>��c��$0�z��؎C���.�l��P�<J]�s1
i�"��c��W��T�����]˞������K��%�.��������3h���4p$VK@j]9�۬� B�v�V�/� 6����	2\W~�Ư�������`���خ��z�{�	lX7+�<=y��W�jrO��+=�8VR��[�\���n��>&`+U��K.��cY!�،�1[�NQlH{��0�c8��)]3�l 
B�z}1 ���%�r�N[���&4Nn�ša|�����b�$\�� rJ��^3����ؾik��x扇�oՠ��X��6Z�a-}d��Z�^$����1q�w�\�HBc����Pu��~q����`�r-��Cn���Й�@�)�8'KT��;ti����x�f����7��'�Â����	�=Ӻ���кT�RP��o�.��qH�i�39O��Ԡ����}f�=9Fz��]w����"��x��T]M��c]|�%��y2�����RF�/������?���98���Q���]����O�1r��#F#�f��pm���ߕ�[2G̛���n�}�>|��_Eb������q�f\�x�U)��}?��߻w�V�6�A�W�\l�����&���@�TD�oc�ch�.�G��6�a�Mp� ^{΀�R���$�D����KB1�;�J��rUk�ԛ͔���c��E�M*Y�a�A�vb��%��Ip��&�ō)�/�M\�u�R�Y�N�0�%#��9���>&�)zA��7܄`�G!W��.�èז�ҁè-7�凿�V?�{~�������b]8hIf��&���N��J2TI����7|Xa?����}?�/�kv0Q*�ҽ���I=n�,\,%!��S6��t� �� B~��~��Fd	�G��C���^��=<LJ�(A��fI/��i���ܬ%���0Pb��`��������i��TF�J_ZvH ������Q���q�?&ʎ���c��;X����S�g�i���Q��Y�;�;��s�gs�º"wO^�	gT`dx�,@���;�e`�3�
ntt�n�w݀mۯų�<�N`2�9��
�k9XƤs
4D%B��*e1��W��l�(��Y�v<k��d���֕��j���X aӦM���9P��8^�S��_�!�4fhԑ&�x��ge>�g�pᢀv&�N�8�p��JJ�������`�r8t�f֮Em��3�0�n3�b@��c��6�N�ǿ��o"fހJ�4���5��C��2,ybn����w�]���f0403���*׏���ꉎ�RN^��׉�O��d6<_�qiRe�DX��f/�/K#S�n�z0� e����5�!���9�������%�`�1fu�4
$4#�L,��0_�jg��1?Cy&�S��L���ٷ�!����ϐ��kPv9���ۇ�������$A�Av�L�u��!���C1ԋ�SSر};9"��kX�ư���,*y��~�F��,��0]R�1�l����7�+_{Ny�����ci�bob����'�W߸g�ߍ�����O4���_���=�@�5@�5�aO���S����i�m��u�<u\�pQ��$*Q��y�ݒ�����d�+���<�������4�ݜ��%���t�J��(��(,c���`��n� V"��2>o��Y��'��P*��+g�~T( 
���ff� ��a�M���&'�s�.\�8��J�新c�^O���>��u�\�mU;�g�w)y������ӈb�
0T �p������CH��s�4?R�|I���8`��4�a�	6�!=C[��.^���â�9���d^`�ʆg"a���4����ʔz��р���|g^	�Q�R��0!)�d4*0ifPQ�e`��.�<K�mm��)�gFF������ܹG�*�G K4Z-*�\bZ�Ҁ8MF�czB��8zY�.�F���9�$��,��̌�M[6���# �"�g͎�V��R����G'��i�flܸD��%?���JC�$�W�Xi#"%�`�'-*4ҭtR�R�D�>N�X[�&M�4�r	2��z�6\�s���w���Ռ~~��"5��V+K��~�S�S��@p�8�fF+@i�	k��<:P`��t^��{�B��?��;�åK�q�Ai=�y��r�I�
;�m@�v�v�NQ�c�Ҽ��U�ِ&�i�\;������=@DB6���q�yܜ3� p��\�\��o�m���#ݸ��#{,d,h�E�2����]�D��߿_�sΗd�Ǳ\�L�6�4sI�j@�1F���g��+2�
�ϟ%R_�Z�묌��L#������Ҭ~��)��W��o�8�����޳�&|�+_#�L$s-��+:�����8K%�aL�ܶu+>�ߥ���4.�Ma��-��98v�ȼ��ȳM����f���Y��*f���jya�*>�����~��]�/�#����Џԓ���K��ӎ1����$U,�gN`��Q����߱㴽6��/����&�NlD�[�`ia.k-�j�@"}������ߐ�	�������&�l���9�ӋLN����B�c��8%����+]�lvLC�:m�lT0N�����_�����@ J��)����f-n��N��Ma�م��`���/>�%,�t�O�晈TN(w]�IK�
��8qHL��p��a������_� ��&�������pB�|6�禲M�=]J��M�I�-���ӧ��#��(,fms�,/�$KY����G,ㆤmݰD�ɋE�u��R擁w��P�LX��5�Z�/�f5��	��SW�Y<���m�)�o5��1d��}lF�	P�Y�Vbuc�2�dv�*�*?�veM3@'U�m�U��j@'�S�2/DӷJ䉠�9�P	S�>��s���aʜ��c�R��i��͍ziG,�\2Ɋr�y�&�R��k����z(&�?%H�����;zUd�z��h�k0�H#JwK;������y�ק�"��a�Y��\���a�?��%u��3ڗ�#0$��b���N[��AMS���� )�{��*q��f���%�<{I���Jd��/a�Z���[Q[8�'b|�5�=�]�KkřDH������G`&�P^3��.�,�j@��bP1���LKw�q���/�R޹�8gY2eff47���gF"!vb;v��#cX\���h��{���a���l�I<�$����a� �{����r�?Y�~��s^��GE>����؇A*9鹬լ�+�R�Q*av�:)��|d�Ю7E�	�s?1%��hh�P�)��5�g�,j椏by�N�"��$�P����8����-n�iu:����>�M���>�i�F'��؄��8�T�$���O���;�Ig?�^�:@?�Kf��Ï�B���R��iD}���p��q�����u�:��t�0�����P�MF
@��M�vb��C��D�5�t)	�i�c
�O��c�UY�`��&0�s��S�Kf�͛��R��X��BM����EX,�X����f�Z��5�׋� �ϔ���0S�x~��{�c�NH�Y�q���w�G>z��)�������k��Ad��ݗ�`~���� u����/5Vx�iw��x�&�9^so�~�C?�
����Kc���aU���f t�1�}�Q�����/1C�}PA//-�;�vh��ɼS�� -ԠJ���o��q�� +uQ�4̉���jR��z�a���7o��1�`����w�<d�t0�r��1�G�fz͌��	`T*����N�mi�7�yD�*&`�RE�$B�ONL������H�QQ��J�gߗD�1c�rBeŲR��n��R7��y�N��H�Q\*/6��2�	x!��5�شq��)��Y�_��=���f2�N��h|���1����$2cժ����2�y_	Q������G��
�^L�"0s]�,�w�ќd���rV��{g�]�J	o}�[�0�!��K^G!���ںDf$e��1SƦ�yֆ�9�w_x�\�F���������@���=w݉#���,~	�4ure���媄A����-Xy/�1��Ac�c��,��zs����D�P�7�f��0����B?l��,u��e+���96�1_4l�$Z��� ��G��� �Q������v��h������/-c��B?s�,%���~	�p�+�u�YӞ�9+�2c�����
SA��P���FْpS�ѐ��OͲE���]�961����k+5��a�<s
8���~X���0HHM3�Rj�F3���Я�^C!�Ò��������� �N�U3���8|��Zmں7�ً�ni�]D��a�A{��>����=��X._y����d���g�y�ǃT~s���y�ks�-[6�ÎM;��+'1_�G���h����ų���������m�l#��+J{g�m0�8F�Ѱ��׎Vќ��/�����c��m��_���d�\� ۰�k<{�斖0�e3�7m0_jv�cDʔR!fr�ޤA��8�h�|�w~F9��fL�(�+���x�|��k��\��c�N�,A9؅
F��b��C��~^�� އ��x]T�6:�sx����/��{P2x֔�q���)��6��X��.�w
�e�ιI2���?����7�-���|����u���|����,W6���Ȱ�\T�Tr���P���VBY�f�W��-�rY,nz�'NO3�W�J��,7>�q*�@�d���#[�V�B��Y��7�Ki{C�=��X���#�kd5�ҡ�J!������W�$.z�W�)e�q�D&ޤNjJ���&�oT"uf�3�R7���Y2�^"��Y%@�)����̮Y+^��#GV�� ��ԭHӞ�i�3cȆ��a(��TF��V��m�IBhʼPZ8V�7�@��a>���]1A��Ȍ$>_YH��D����paH&3 x���F���%3���|(f�s�ȼ�ϝ� l?���o�/����ݖ��?��}�c��dޚ+u#�n�~�ӑ�67�,�~JyK�X�랻%$#�u�֗9	d���+��]I��66�*��K�x��}?�N��b�,s\o���roJ�g[d����$L ,�0,�s�7������NΑZs�J�I�:$���y�M����?��5�y�OmiE���E&���2ԹV�RI�L9�4�i���F.�%k���Ȍ<����̌[�kB\?�S�Wv���x�,5���փ�%�l�ҰdN �Gؔ&c�h(�<c1�	�̐�+ł��/-��!�l�7�O>�|(M�E��9��0������o���k�����F�'�����(ɡ�B���Rf<@}�\#�Pn�Nv�4pK���;����f�����G1^�H�W�}g�M�$������6��GŐ�����S1�?���ai���2; 3@̿B4�Ę���
��:��    IDAT���$���w�������PU6��������g����~/8
��H�b��a���W�$��.�4�v�Vx�CcӰJC0�xA�5����d��0q��I�Q�ͅ���x��ϼy����G��Z�<�S(/������I��>m>!�t!ݗ~�.���RQ��% Iu�C]_[[B�IM2ș��^zaT
C��'�r�n��W�zL�LEA����r�����z3�]�=�#��-L���q��6b��f�-�|�1e�����g�5���8� �c9�ز�Z���r\�!.��DI,�4��e�.s�I�zbjR��4u?CC�m:3��f�l[g�gYɬ����J��Ⳉ�v��r�3�*�B��f7Y��@J0暌UG�y��2���5ݒ7K�˼Dޛ�ͨ�,S��Y�,����V��CBY"��ga[Z݆�t���xV	�$��u=��W���Q�ie���nX]��ŋs�<��O@;r������K/\e��<%a��?�dkJ���^'� ��$��a���x�f�E$����R�ɜ��R�;��}��<�RE{�4Ĺ�Yr@ M"�3���X���yo����*&�..�D�);�	�I�aeFOXIR�7�t�Ŀ?���霟D���@�,��$?&�)1uۖ{҈`
N��o�>��R�L���R����de|��:Y�:�+L����u��UB�uhq��2�E�av�Z��{�PY*)s��:�W�\�K�����:�߼/<
+_Fuf=jd�r�g;�������� �*s��F����>u��Sk�L�G�Y\�����c(�
e���R�9LOOp�?}����o�ȃ�<��uɂ�FnY��W�\`jbG@AEx����[YB���-��

��M�\Y��$�I�]�.,7��g�Ŧ�q�}�ǩ�94>O��ĄX����@���d��o��������\3��ɩO��\J��
3;���O��#�`�P�N��#�9]��&�]�̼?q�$�D���[��7߿����D��{�:[C7���P9	�*@ϒh�t9��ItД�?���h�F?,e#]��3#U��SV�|	��G��0�arj7ߴW���1�,\n���R�dY�VTv����]��aǶ��?��s�֓
�ʙ�&�.?�Lw6ߡ��i���!���ӧOiO!�{�)N+t��J&�%��&�Y�?������_��#��M����l��(jB���}w�u��'��K�K��$��K������`����J�/}��-�6�gE�c�<��Y� ;�I���`��v�����C��LkvJLGa�8v #C�-��s%�w�4l����W��r�r	/�? ��DŐ�tE�3"IT�f\��M�ds̸'���t�c�Ҭ��Be��4������6�3J�6i/��|��@�铟�$>�ψ!B@������$\��@c$K���ה;�=N�\e�#���~p�Y?�Ò��Ga������NqL���=B���M���M��:���}.Y��s��?Ęݺc�<?�"�&24�wR��XE� _��r�$�^w�-���c�yT�{]�ac�Ҽܟ�{iP�Y\���9.�'���)ϬN�����J�@;IYÙ�0�<s�{4,XSO��w���$U; �w���LQ�fa� ���o[�J�d���z�D��a�"������19�C#�xq�AT�'����p��'8��+��������U�~��l���y�?\�����!�o`˚x��G ���q���I*��J���n�7���w�¹S8u���-g9W�C��e�HPjS�in-��n�_6\<y�<�*E����%���m,_�����	�
�-��W_~������kw����u�G�ulGw�S�蹱%���o��
���ش��R� ���dV����a�TC�g��%�<�u�XK�X��W<�D��2{Y��+g��V�xPõ�F������4�Czȱ�.=���'������
��]@|�r�ֶT*�l�O|⏰0��˗�P_i�Z~�ՙ���i�L�b�nY)M%�X6<7)7$�6��5��y�F��J�	c�c�qi�9��P��|�I�����+�ݮ *�J憧\�0���:++5Z����<��.=n����oX�^���8���F��_ ��&=
�ns=d	�T��I0==)-M��e9`%���Y��>Z��' �H �ʑ�睴2�8��Ǒ���y��Y��Y��~��e5��P����N?�;Q�<Y�XJ�$�/�K�{R���W �¹��.��X���Go�c�<���� �� ��s�]�9J|&���1u�#��*�kp�y�!�����0[)	���c��>s3��HX��{�B�ݖ�������k��x8w<+��GØIT�NG �?gc�����&�>E� ;24,)���С)]�%�I"\���r.�'A�G�f%�4B���2�TI�A�2bP[����?i	�K8P��uk�<���<I�c/	ʢ�C�Kr��O7L��i�DF�$Z4X�9��1�(�˦0b���0���y-�#�C��?S�d^:׋7Y��A"͔U�d�-��˟�i_�gV>ǰ�ypt��.}#s�}��rf��y�n*#��v���i��g���+cv�u8�� ����~����_xﭻ�\i�������?��l��_}�W��}�* bkӕ&�zcy�������G����H9גX1����Q�8��E���2��6�E�w�����^���סv�fG�M��2ʅ�4���$ **iP���l'/\���;�o}�����t�e��8s�<f֮����e<�9���Wpi~�]B�4
ǥ��{gg�ryH�k9�V��������`+��pO`���pu8�R��q�v;O���W�nՑwx:R�������}���� �v���{0��T.^O�WOO�"��֡�s�8�v�_��W���R�Vw�b)���0�R�,l��6f&'d�Kr���K��4��S�4�J+����l���
�%9|���M&�^3#L �ᱝ�ã�+!���-̾�M�,[֣���L,���V�XXX��PYփ/*���Y*}�D[�+����⭉��	��"�D%�z��	��C3�iZh���1�Vb��Y̚m`ƾ�+�`���P�3��
���$ ��I*w>{֠E{�,U�DL.b2e�Aw���1��W+4L�#��ug#����Y�7��������5��ݱ܊��\��E18�3��	����^��Y	��[���{��9��!���?3p�5��4'=��	<��7�[dm��s��ܜ;wF�l����Z�������)zu�����L��,E֓_��:�nd��|�z���tV�BY'��3������w�`� :BJ�v�,&&�$�e�̑`�2������B��i�'����ц�>@��LYɚ]�m ��^�L��x�i�)Ku����`\5k���[��`�љl����\#���8����J�����bVӈl�t�"��e�Z9?!y��ٹ��F��a\d) �b�N��.�dB9t��R	������y3�/�,�����z�Ov`%�`�q�3�6I�Ӆ�PN#��0�hB��P���W~��?��� ����r��/|�|�-]2��BgiU׆4���7ྻ�c�Hy��g{X�>�	^ǏB��:R©G`�ޔ�|�~'�#n��|��!����ќ����F�.���>�g��C�ﶣ�=?D�݆�0�<��<��C_�"~�~��C���t�E��H���4��~�Ku(�E�8"��
q�h��x�[߁w����'���?�	�n#� n����5�(V��h$c�%^�󡓘^�Nl�p�4*a���_�����bv��<�d���=���m��\��ݥn>"t��- �z�|�+_������J1KΨ(���y}�}�W.V�����j41Qeh[��NZ֕y��q��eYa����铞�咀���P�+���L�bk5�bq��
�I+x���:���j:�T���$��������_/�y��I���Ln*pR��s�1�6z~|6Z�R��Ö�� L�t�e��Ԁ☲#��� Tx��e�ٳH�Q��gh����(U�x�f�&����N��:Q~��:�;��ڽ.�~�˖�����sҹ���J{Sf�K*gZ�ϳ�,CV:'DDC��s|���hu8M�S�I��s�ߥ�f��kĥs�3xf(so���b��jc��5���/��;J��j��yr�4� r6�&l��`��F���&�$�069�A� (�������:���~�[��ޟ�b��i4}���瞽w��U�����͚ж%N�]��jy<GFj��;_Cԡ��W�r��5ȇ�cPɴ WV�=�=Jt<>>�&��ȌԦ���Q�/�c���'�b�%i�0}w�WB%�N�	"4B����z%�D�����11�!~ҭ��W���(i$����J2,/¢/�t&��4G���r��<8�P�`�]wAG�X��i6�$G
�� r��5JG2�
�p]�W��B��1mc�����1��]O�_��6I��.B}c�V�D����nɈ����i�p�D%�L7M.h�G�A�l��%	y|F����w��;}�p8��1	�3���l��tD5�La*�5������^W>v?�%���[���T�����u��j��ٗ�����	k����� ��
Y��1?�[LoB.�G�D
��V�UX[E�D[� ��q�i.]Ҕ�)�JfD�ٺ�%��I�2{zV�����\�̌�@e* f|�\Mqmd"Q5̅$-Y}<�ƛ�<{[l��.�f�:x�!d
y�(/u�����q���� ��a�X����>9�Wq�o/�n{l#G�cv��֚�ǣ?Ҭ�[�	O[UX����9�j�f>�_�M�q�D[SW]~��95^�/p3��V�sȹ�WN?*9�ŀ^v�/\��>���q�\�K}�ƺzi��z���ȌF�j�W���;�� �G`�Q��(�%����MV��s�D:��f�(�\G�	x?�ԃ#�� XJ
7
:iq�:���/��� �x�q�1>�i�2f���8��N&uNDr�aE���x"!$RҒlܢ�2P�٤���^g��;�/V\���?W`����Xd�
҅!�YqV�d��#A�Ӛi����M���ȳ��:�eU����>�M�l�afg����mɉv\��iY�&8�
�H=j�lh�;��B����x��z���vu�(�m
�b�ܼ���b7
�ݽ��6ySZV��~����U:��<'��);n�ͬ�ypƆ���Y���ꔒ�|�TPx ����;��|"V�_��ۨ?VK,l
����WǙ8`��Z��A$R�6(a�ϋ$�dj~��RB{�R��`\�\s���"�_�v�8I��z�w&A��I��{�Ă|A���\�:oGS��k�Fl�>'����n�j����.��A�,q�j�5������Ug����č$X�I&@j�V�"�9��g��p��l���
��ID�Ї����Ux�ߝ;ﻀ>*C����v��oܵ1[>8����*���Ơ�l?��c��k[p���~]Hql����|� M�d��f�
)?���I#�Lal�e�����w�����0��C]�*d��f`wk�3�
���|Mt3}x�_��7>�r8�+V�;�Ǳ���]�ʤ��fe%/v͛�J���j,�j���j���ԆL�"���G�3�:D�o��I<M�`�H=RL���c�"�U�p;�E�uV��3v�%X��ӉukW��!�H��������T\z�9�jR�lS����z�Y٪���O�KЃ��} kA�������X�b��.z�w�߈�Z��ͤP�XH��j���:�3Uu*�M���K�egcw�n�
lN��d
^���E�w�;�yA���Y�S~�7�IS'�g�̟�swo�H�($�q�y������S���?<�`����[o��u�QGc������@�@�U��:�]ׯY�p("�԰����a�����+��[������͜Ƿ����5nPDc�9HX���
����ʲ�	3��7�-8�fT�&����M�a��r._D'�����j�H���z��������߱��s5	n���W�b!'fMX�m�ؠ��Ii��Z��V��ɒc�b��c4ю׎A`��U҆��4��y�#f���Q��a���eH3p��l����'�S�$���`��`Y��""@�2V��.�n� �k�����4XAɰ��%�\'��F|fI<����&���hD�6?�QϏ3ݢ���㘱��uת����w܁�T� 9�V���e)��X�Z��/ϋ���g�v"�� ���h���]OB�F�}�=�{��	B�T�p��,��?U�\;T�db&�,"�����u��/��'JK��B�x�1�L�g�����z����+.>뻀>�b/�W'���W��ɹ��$c]���>���>������;mM��l�TV}�@���|��3466�TΡs�ZUhdbV	�J�Il{K>}�]l;uZk��ő昙�#_d��-��`�l�.&B="��H�3(���ە,Up��?��x%�c�)m#W({�b�_q�^�\���k��R�͇D:�1�:��λ�Y����#R�,ȽP�i����15-v�!%q��lY��L:�x<�"j"^��7\�m���3O�fu:;|r���iVC:aU�D�TD*_@���+���n���X�z�4	�n�ڳ/��مtrH��A� ��UH�3�:BЦ"s��y=�T�V�D�����y8M"ez ��s��m `E� Ξ�*�G�O|�^t��C�M؎J�Xd�3H��ƫ
��\�r������ YJI�ޛ~��H8���'���/�xB�-���KV�ֳ��O���& ̌�b���\*%BY��hؼ4bK�a6si�ԩ�>Dbc��d��	y�2���y#�_�]��1a���qF�
F˚���@�<���I�!ӓ��v&����U�2��`�Q�x���zu�>`�Φ��ĕVs�W����鏣��h؊�V�����SX�)�e7kr�!?昼o4M�H��*O�?�3*e��?|_�CS�+���MgS�9cK��Ձ?�C>[�oH�rGBg�M�0�����S���Dq]m�H���$~��BQߝ����6!?�����U2�~1�`ߚ��V#�N�թ8��a}�\|�Ŏ51���"��P�JQ��lo���Uy(����������[`�4����-bUGZ�\�L�G�\CZ�{n��?�
��}�*�m�`[�@ȯn�Ȫ�~����(�x�e{�֪:��lS@�����r}�?�N�練�({�Ε<�f��X��w�����o�����.�Y���%F��7�~��	&41�%	�В�&R��wKc���Cl=��Ѡ���{{t��S�+��/�q�H���d�f1��!��bњ��˗��aG�3�>1)��Y&n.�2.��J,]��P[P����<��Igs���X��9so������Y(�HM\��1��L�������^��&��F4�G�D��;�m���~|��z�5Iu�����j�T��՝�>v�,g����E�d�7��=����V,!�#9Ї�`<ܰK9�a`��:Mp�:�T�b��i�i*�w>�{���٘�o�w?�>B�%tVcƬ��`�����ѣ|�]w2�����A�o�����ˤ�3�|����/���� �gܙN9������ ��K�=3vu���'�T��AX���A��IA6�FCm�>+|n�V��"��'�Pr��䁉	+�#?R�u<67�X4�$����#��>����
��A��B-�o�����|,Ú�	h/���}�y��l�ȶ��0)�w
~ؠ��h�0��3�B���b���|�#&��s�	W�g���6���p���$6`�n���}4 �’l�\�+�VG    IDAT���֥�`@ <]�b�=��a�jd���C������������z��B>�i�5�!O���'�n>�LA��K���r�?�G6��{��g�}^�C�{�XSR6�C�!�l���z�u�)������e��g f��k��a�r� Q����M��^c���L���K(r3�s���;A�3���gm�mfo�� ��K��33N����_�F@U� �ʶ����4��H3۪����܎�s�	��y�17��5":��ٲMˑ_�-�i��B�{6�b{��0տ��p!�!$'A/R�pc���(�P]/\}��~2g����<����u=��r�|��+�=Y�n6i*�{���Y�p���c��D!���!� H9-8[ۚ��[C�-��$����
n�_}� ��0��	Y�.�S�r�2TP��0#�a������i�sEd=,Y�k��ã�E�?��i��TW���Q������
,Z�5|���t(��üP�CT�2����M��@2WF��A��5�ml�
�V5j�[�*���l�lc�1�)0�ߋtfH��UBJ9�6Ű�6�������Sڴ����朸��U�
$R���E�j�Jt����A"�CooJL[����������K��4���΁������CB�2��7UM��@�/�QY�;��M���"!�v�S>��p��S[o\�XI�vc�f�aC����;$�z2��'�<9"_z�g�4�l�[o�]Jv�6���1 0��� �pȑ�����TnG�RiB���O�Qm��	mr�r�^�B,�t���-��"Z[��g��\ �?7!Ul��DBA���ly-�;�v�K�D�ؒ�6��F^O,&I� �J��D(��5����c���&������dՓ�ϭ�����|}]C���7�#�_n��m�O���lT�7*���g-D?���dB������:2�;�����fT�wL?^{	׹��I��p�6�a[�S����'�A�5��n]�L�j�Y��hZ�a�z�6I��`K���ʦ�deg}J�����n%�\�dċt��k�h�s�
�1U��
��c$���|�|�룎<�r>[��W_{Ӧ�Ę�"�1c������8\/V��V���i��+0Cԃ�юn�5������7_o�m<��]g�,�C���F���+Z��ir�e4Y��>�,0��6�G����U�.75WQ����"A�p�����dδ���X>ސ�~�so�9���Ud��+�)A9Gvx#~��6�w��($�����ۥ��J)�����0~�8V�Z�P�T�d�����26���˿A ��N[�D׺��sd*OU��9ʅ8K�+�fD�d�d�^��Y��n���>�yo���0P�\��>�|��Lb��~���sl���U0a�4�L��|�>�A�|A�(�ɹZxPr��
� \�_�V�m�b��|�o� �M�?;�biӹq���C{}UDbn��l@��Ŗ�'cڔ�h���������C*�A���39t�'�He��x5(W��T������&��N ��P7\��4��]L@�jv<��d�P�&l��moL��G	����\�h�bzg���0׭ݠ~8�eYI�#��`,A�G�@��(�����6�on��>�,ZZ��|��*�y�R�I��}G�K��)x_�\�/�9�<�1��P���0֠v��p+8V���6���
`���W�G.��^�c1dhAj��N��=Y̸��hp���-$���v�LoX��W������#�,�U�hvKJ��YiV��t{$��m���#�����Gv����r��
8|�qlP1S]�f�k�V��)�6ꏎO������G�k���`oߙ�߄�p�7P���zcbö[JTV���^'�l�X�4Lb�u�Zf��@�s�ƹM2�r��,i��?9-<�J6��{�ѹ���#��i�CĀ�ɱ/��[��޿�}�O�P��BQ!����ͬ���3�|�L6���z
�]qJe�JZ���uA{&����<�Z%N!�`m�r�X���?g�z�ʜEUl@���v���L�f�-{���:����kI!;{:��r���h��s>Z���8���!�)F�S-�B���ͯ}��ӿc�ۀ�Aon�ߞx����)�C��h�H�� �C]��޳q�>["� �d�K���1�N�U.a��-�ª�%#� UT����/��� �}�!��cW�3)�	+��Q�L#��QeR��QΉn��ٯ�4�W����/a�.{`��["M7�0���u�s��ƥ�]�ϿX�hi�ں&.���n��1`x�c�^x�Qj����j�>$�}ʌ�z	En7U6�(��p�Ňe�*5$?����2u<\�R�^��D|��+�{Ɇ�"��`(��'E \K���)d�U�#�Jd�i���VD�,�]jh�� �Uq��I�ˡT,�^�R�kl�����l�2�a�1�q�_䩚�:1�����_.Z����+���� 8��/�=�P�{�Z�RŁ�)�C�2��πN�>V�d���:�����\s������4���2�����T҆j��E0sLI�����u����6�2P1�sl��U�2�O��ц�m�v��I���e�1�=P�q��2_)�TE���0I��+n�1^w*�Q	������)�6�'i���*�Y�A� p���O�VF�^�gl7qڄ�jF!���l�����|��	��P�Q��,��q���sr�����T���*�k�$(�&��y]y}��Go�v��&�����;�,g����xXb�%X���k�,�Ό�G�sM%8��7����QI i�;G%��1��e�k����w&�b�(Pm1��D
��`��7�4&�\��M����z��.��=^{�M$��#1�g#�����;>`,`�@mu�-��̈́�׍�)t��A�6��q?�|<�D�J}�9����e���o�w�v����f����w�">#K�8�q���<�Ī�ʡ^\$��h���A1��x�o���w��� ��Nz���p��+V�(�JV��sQ�f�X��d�(�R�Puh�lV�$am=k&2��6�G���D(�I���5~/�|�.��i���V䆇�*{B�M���d}�W2������L��������,� �1�"���^vz8n�T���ҕW�˾])��/F ���'���B\cS�t+�Q����ԩ:f0�]�F��|����x�KZqڸ4{����EM�2
�xJ�D�(璈��h� �@&�����^ZVP�x�!,]ۂ|�T���C:_��i��^.7�D| �La?�:�:�8�ݩk_4�F�@X�H����2�|^b,R��jMY����2����e��D�y���1e�4445ᕗ_ø���kہ_�������ۅƦt"Bg_���TY��?7w�\m������{O_?��hhn��=��:�8�`�z�(��zc;�8�0nX��͂��hR7���q]�!TIV>�s��e�꫒�hF�(f��-��w�+�ꉚX�6�^�'+'
�2#����\;�y,~�Þ��^��
qN �wI�j���+sC�d�C���
��~���n�#n@���M���X���WB3�nZ��n�kzx>�l�0`A)"Z��9��QX"eS��wU7jKQe3��aB[�
�n��m��?#J�s���klP���#e6�Sit�D�q£ Q-Nި��t��+7CL ���]B"Fd�sƔ#j�Q[K�y���9P��7:� �p�qz��|��JHe�/���i���J�,bb�x��k�uk֔�0������� oӜ?�S�kh��LP�>Hh\�Xs<!=L8�@��ߙ �J^DBGSj���웒͇�2��n�Z�ᚚ������aWu�}ϼt�@%07�
"7�r�6̧U��-t{�TQ�$�b�l��,�a���H��йa��լ�sٔnt����q��W*���.�Vӧ���^[�^kM0$/vn�.G���l̓:������o �|� {�� 4����]}h7^z�P02�P�W��]����X��.�Ʉi=L
ՐG��Z$/K)j�{|[�G���R�c�7�"�.F8䃻B� �z���h��,Ԋ5!T�L�,xC��9�}U���PJ`���(��Ӛ3�C�nN�FFB��d��/��Z̚5�ب��cՊo�n��mmB:E��<*�#���GE���2�b|�Wn��(�bfY�V������A����k��<a�$s�	"'=��c�4q�!�}�O���
ֻ�<����ڰ�FC��x\s��䌚XZ?N���sDv#bC#��R2cP��Mb�S}�RtDaL�¯"�kG$����o�w7�lL:L�'�l�T���7a%@ܨ��/d�:���� i
p�EL���$��r�:o�,�7��ܜP��0�л}f��u�X�:U�ZKNϖ0n���`ʏJ��&��r;Om�Ò�F�[L6�&���e>���Aǎӹ��>z�NLr��>��y�θ?%x�}�`GX�&e�k���p�R�;�f9��ꙥ�N�P􇗆��DR	;c�O�5�}qĲ�~�/�v�@T��0V^�gd�[	�S��Ϧ�❫�h,fP4Ώ��Z(�-h�Kn5I��n"=Ӝ�%��p@x��=�� �ᵆ6���kIϺ�v&f�����O�!-�p��i��eǍ�S\����G%���ً�d1�s�b��8�� ��� &D�S)�՗����s���G=Mve'>��w�WBs3U?�E �L�C��|F�� a"WY�0�#�u�_�͖�p�qG��gr�!�B@��1f�dT�rfZ�L3V������j�d ���TF��'oz�ЊU����J�TF��GwrO��*v�e7��>��3 I�Xc�3Y��E��$n��H������R,�f�Z��4��A��x�-U��[�8x�HgJ��4�ɍ}�X}k������4�Ķz�|����˒|U+��G�����NeKX��+V첯����S&�ú��b���.@��[z�����&��r���T=H�����Sa��g�=�Z�\�?�q8D(��2yU�����6�L++�P0��5+V�{'�9��{�L&�/M���7D�yœ�����΅��+������)��#8蠃��s��믾�I?��f�/��%�ѡjj���h�<U��mm6C��ѯ��+��=�Ｍ�m1cKL�6�>�<��C"{�jee��kZ���0�+UrA��;��ԲpH8�xa�hbSj�s�$)J!-Hh�#_�ha����Ȟ�<R$����#��L�ژisƁ,���Մ�����F(2g:	o��<ܰM�l���|h�/W{�n���޻.���g��ʙ�;U����37oa�͗	��7Di8�XS��D(����`* n�j)d�:�
&��H�"ڌ�@�\q��A0�*r���f*@^OB��E�{����X��W.���:�~~&o�y3CI�67 ��"�븙l
�u�� �59.c%��Z�=Gcj3��Qb��kI1�2+b�v%�4�ŖmB�F��򴆨VA(lf��E�#~��Y���z���TrK����"w���E��
[���X�:�1I��M�O!���GI��m�~p��� 9B��8�3�:jf��(��8�3���	���|�x�� �.�������MR�`��e '�J7�5����є�X�j������8�;a�Q}��섻�y�ξrd�l��=d��np���R�*2��K��B�J5Q2���6�i�L�t""��DH���0��2~^{�d���sP��k�
�54!�H:paU08�0Hv�n���N|�pf��{�3}�a�����ߞ���R�]�,��d�ӄ��K/�K/Ek�d�e�Ň0a�d�C����P>��ĵ��}��@�PUPoj�@ C��twnD]Ћ�-Q\rީh��RΠ��\*��A���eu��W�8v<������U�~�ͧNE6����?���&�l\����M'���7��n/�u�
$�PT�Π��ЀH(��˗Jk���E=nhʸe�\�b�@6=�H��-s#��*�2gǶ�K[[��!jOW%���47% ���\�ZkǸ	Hf��s�}��koi��0+V���)������п���m��3�k���
{�|�m�ɍ�Ǖ L��Q�����ѿ?,V2�{\��v���'��c�z'*���V=V�jT�6�t*�����9�1Š�HE*�?�1QԆ	M��I�bl!yŵ S�"6Lv(
"'@�5��A�U��*8c�U����m����[7��Q#T%"W�踰�q�ot"Y�x���ճ/��$W*5�9�l�ッ#������)�t����P؆V�2��ufp��e@03�&�6D5�n$�{����PR3*@()p�+m����Tb�=�m�Ur:�낏�����Ֆ��\��� *r��}�34dl�h�C�d�&��A��U�-5A���(��I/(u����ؙo�s�t���ֳ �@�����)%GGJ8�J8�M#xc�mF&98�XS��~��u��s�Tv#i��1{��HF�*�vv�~�?=0����u?��R�_��v��cZ˜R`��U�̈́�$SL�xx�ę�9�i;0xrP.0���pWb HU���X�rUd1�	�ף�v!�*`����xمg�������N��o��[ퟫ���#N��U����څJ.#R\9��[Tm1tu��>����Z�)jk��l6iE;չ��
��X��l=kW��:�oi��� �L¯ L�"�y*�������D��:6��;�@�Y��t���ǸͰ�5LW�/�M�ˮ���_!�A$Z�b��3>.V�Qy,�!W(+x����E�5����P�׬G[CB�$�:�8Lۈ��fg�ks#ap��E��@�H�7�u���ٍ�K�bζ���O>@����I�Nı�C,,��X��%P,�>��I5��v��M�����M�Ɩ3675����Ԉ+�t&��jgsbE�J%�W@�̑.
�p��}$��o��6x}��]�8��5#m"����;c���˅�E���s��_����$�>s뭴2xs���P�jK�.�?R�E�7ɵ��Y�2���{�_饗b���rb�����?���x�T��t��(�s�om	�r�Y0�if�
O�ܳ\k~�H��H���0�*�5Lb�6$�*�"E����T���*rڸ�F���;��wn^�l Rm��(�&���;mp����x$"b��g�#RR1�kU��紆_	R��B�&�1H0uG29�^1�3Ʌ:�h�mQ�ݨ�5�S����B�T�ؒplo�T�V�T�R�Z����M[����GɘZ�_�Œ�~	�3�!�K=�Io�[$Q��M'3hӊޞ�w4;�eϑ�CD��	Q���:i��Ւ�r��,"�I+ôrz9FJ$ŧ�9�%soxlJ9�BZ�Nl2�3���Q�ڪ��&>L��HsDN�Gި�1�`E#y��[[�u��y>�|�y|Fm����mmB9��S���M��������I�CChjm���N4��4�&)T����kZE&����<9Ob�P��E%a�.�]d�LK����~���Udp��mGu�ӅS�ps�ເ>*���_	�������&�Z)Pf��u#��ZF�M�w�tN��b>�B6�R!�#~t fL��T�^�#	 �IGD�������ӵ,B]0���X�t)ܬ"�Y�h�!���r��Hf3hnmAǔI�|�������%сb�8�<a�h�X�>��au��^e�_~%��f%B�Dcu7��=�(2��{�Jg��
>��B��'��+�"x�!4��A6S�ؖ�)�vީ�bj���k�r�r��Λ
$�b
F��2v��ZI���鏏��=�@�q����������Ť��������H�<��a�["RS���^m�+��¸�c�L�2Y��|�|�_��ޗ3GÔ�k\�>�du{��78�Ǿ�[�;��Cp��)X�"    IDAT
� M@��_�f��6,_��(�Q�R��;Oi���ݍ����L��E�kj��8��� �����oV,���{0��@GF;=�Ǐ��wݣM�ni��Ѓ�0�-]��N<Q6�W_}��
�3_O8�Wg��Xm-��{�طl��q�a�sC�+&7����747֒4F��4�\I:
D4)AF6Mn�����_��l�dF�X�RŁ�9W˪D��N��@�f�RU*v�)Om���T��J.8w-�;��"��~�"�J�� *܅�&@:	{����咪B��: �h5�'a�7�y�-��*8���c�	����$��$)��?{�����{m���3�%�?��9������Emȅ��\�v�ZU�s]-W���B�ҷ��=98���F�Le��I�ܧ����2g��VK��r��¢��U}���!l��>y<�<�M�� !w��Yl�fb�H�*1d��k��3ْ��c5�Q�V�4�i���DM����ƶ�;�۹.m����;��c#�=�?��1�|GҺu���Rm��p8$L⍜���B�
n\�U^?J�d¢��ϼ&��R���`���|9Rޖs�uHЎ� �i%����0	 $����G��U@G5Wl�^��B����qwv�=Ͽ5?^���9�r>�(�\�b��=s:22CC�|��E�R
�PΧ��R���.��9|������J����	3�b��\�T]��W�\-���hlmAS{3b55p���ú�]���!��L��RU�a�kA���ͩ��{�.GOw?|� �.���ނ��'�ù� 	lƺ���]=�����!��Z�ח�G�}	�?�hЇ�7�?��<�k㛯a�ڕ�d��>�PV�H��'�x��7�Œo�6f�t�/��y��?Œ�_���y�`����٧�`��5x��bٷ+�٤]�*;�q��˵�	
!w���6�l~s��H	~{�����o
��&@!tU�nZ��VX���_}�5hh��5����p���%	��(KJ��dN�w0�PU_u��qc�~��'M#5�B]mN��i��]z/V���'�����G�o�^~�6�h��8n��h����>���W������FÒ�_�K�k���U��?c�L�Њ%YG)�����|+L2��~����KhmoC&�����ʥ�Î(G4�2Uu��rf8�`�1j!/@�b1t�~�CV����f��#�C��cFa�A�T�E�̨���&tuv"H����2P	��X�Ѐ��.�,������\*U��-`�ƥ�:���͠	�<o��)GXѣ�	+0�� aN���0���qc�M+ϑ�z�̝18+�c��,���Љ.��1c���e˾�$v��LvlDƎ��H���{L_���oa�so`�wi����������J��!o�x�Lb�{�T�î/r�)gb�E/��o���|������r��usC������
-�M��V}#L����s8M��M��T�.C|8�L�b���*��]�֡}�x�Gk������ئڰ�SI��uk�4�ɑ��w��vx������'� '?�9���>:��7�S�q	�e�S�[- ������Q�]�Ǖ���=3�5HSY0����` �DKG��E�j����Þ����ٿ>r��4i�����O)��:�_��D�RH�.D�d��0��/���l�}6��E�_�,ii�AA���N�	~'JS.u2m
	2s��Wh��pЌxQƕ�-i����QC�^��8օ�QA:��&;Lӄh_@pt"�B��y���Ud���4�ι�?��3��@1G��c�v�A�iם��ڈ�dB�}���hikC0X������ c�MA"��-��C��iȦ�����0��ݝ�@�&Foƍ��Ȩ�r��w>�����{q�����%���Q�$q�Eb�mfc��/��k����Gwo�a���UҚZD*���7�<��,�Z�q��c��w���&�y�'�z�H=r��騳R�bρ�*S7h��ꪫ$���������7v���AJT���۟L���j�� ���Ki�󼆆S�a���78���܋/h�>}*�O�/��`�}��v�yW���S�F1v�xͤSz�r�ܔv�e'\|�E�͈+Be����!��λ�ۃ��1����$lD��4��Fe�� ɂ����'2n�D��$����yn��l��E����_1�����Y���+�m��àJ�a�ZA'a���ղ�	�g�+n����u�Z�.jjb�Z�͍2��3g��+^W��u��A����D���b�;I5�/�c�E�}&O�e�H%�q�J�N���b}�m?�Θ�P���K���a̟;��~{������[�l�2�5��I�*5+=� 
���tV�|��iӦᣏ>�믿�Q.���y�d���n�1x�L��o�EE���ˍ��n��>]�{܄�X��k�pT����A�����V��j��p��n��<�hXE U��^�Ԑ
y�jkGFC��#�NB��&�p˹��'o6��sN9��X��r�4�a8G�1�w�
!���5
��X]�]Y��?/[g��8�V���p^�����}��5�������V��R���O<Q�̃>������i��)���5שIR�J]��K�@�Vq�I,��4����i�SO=��X�z���x
���?x���
T�Lg%�M^�T�`��*:^��7��]@�˼�S�����Gt.���a\�8�������<�:���#�f��Xk׬p�7�j��8VR)�˰��M�2�z��\n~DCU/�DJ��p	���W��l�"�9_{��(�p|��GWO��m�}��C�c �~��*P�3%�)U��ѥ�p�U����6}�^�h�WH�r��4!i@o_
��m���f��g_Cm�8�h-{��W��ރ\2�H�o��>����L!C}�r��)n��N��E��O=�x��gѵq&t��fӦa|�X��.x�g��Ob�FƊ
4���5�Ɠ��NINt h"B��쮻�/��>5+O'H���z=�K�53+�J��Y�fa�	X�x�����z��U-�:����W� .]qf�/>�<fo��$+fڢN�:;�#�|�imz�hoiiÃ�]=�=��x0~=�|m�mc0y�d�]�]]�:/&MM:���^mT��'bAh�S�@XY�B�x���RQ��D&M��j��iS��a�]w�����x��tބ�1qM�<I�d��K%1c���|�i�֊��zNm	Μ�|�)X�d	>���	~$�יM���$�#"�k!h�/��d�$TI��O$�P߀drX�{��gk��a8N�VUu��t��� �h����$��u�$��#u�e�갤9���a��EN�=��ǵ�k�Ɗ�� ����CԵ��{p/��"�{���k�E$Vk����ᦩ��]o�t]R���Ar�f���k�ꫯ�z���?V�H���֩�cPa��9I#�a���Ԛ�T�붝=�7{��9�%0��M�L���&�H#=g
R���nL�8�'N��）��~�a�g�\��ч�~��?8�+���==;~�,���9�u��}�]1}�4�����t��rk�Tȇ������E#0<�a��-岪v��2#����n{�g��Ɋ�ͷ���5F^�_l�0��q� 2�/_�� N��/�o9���ѷa#���&,�v9��vD�[M;�i%� �Č(*]ݒi�Lh���IZ��J�$�	���J�(���0e
��n<�����X�f�>#�mgo�c�9g��WZ�[l��x2��^��hMC�o��!TC�*�o�^�⢳���O{���~��;�!� ���Cy��N���v����n�o���UA_��nxk[�6��� Z[���G�	���-���g*FE�r���<`����U�K%�J�8���e�0W1��"���Y�r1slL��^*���/Z���t�[�1m��z����_/]���v��B�Mx�ŗ1,BL=�u�#�c��h3	���]1e�AW�;��"/��-�b�T�����`ђ/��'#�9w�|�C�}!l��v
��<�j0�����H'ND�رx㭷�"ŖC2�Ѧ����˅��V���E�nB�x]np4� q�W^��"�0Z�vv���kd�KL��18���I��۽�K�ǌ\�d��J��2�P����>V�.MK≔>ϳ��f^���iӱϾ����^զ��>�h���VҶ�~����s睯�7g��L:���u�0{�Y����M���>{�LT��L�2O=�,n��VL�2=}�#�`J��3�p��8����g�R�:�������G���O��Љ+��C���0B!F���ub�8�z�M�z�Bm�3gn�x ���
���T��^��ͿS�M1���K!�],����~���LH�;SЦOM{~)H8?�����~�>n��I��W��/<���[��g�c�m�!\O%?�E�q7
�x<�~�98��3��_��'��8=�0�p�	���+0c�L�������4���fYI\��v�LK��=��sx衇������a�}�A8餓q��?E��a$�$A�R#��i��ӏ���u�B���><��c�46�����ե���%	�]9ҭ�벷�2v�M����}���3���e����W+랻���̝wމ��+��74!O�1	bU=<4��v�'��x���pؑG*�:�����߯�Ы�t���k�t-�13�k�yw1�����p޹�b�]wÆ���'	�'ʲp�b�e� ~��Q�Ԩ�E5F>�z���C��矏���/X�r%���r|�٧��;��o��W���mY���o��y��XI�\�B �ߏ���约?���8�C������7�3��.��:���/ttLP�͖"�n�$�V�ǟxF{5�Aԡ��A�:�\?>�P��g�~:b5&���᪢������L�'L�˯���>��~��� �A�j��b@�KW\tּ�*�Q�ӡ��{�y��x5���A�]En��8�Gs��GK?�y�r9����s�����|�l��C;�C)�-�*�@�:��25�-�>3ko<7�p�ƌp�WUUEȗ�)����de!e"
J8��A�?!e�ԇ'�;_B&�Ess�=�<A�<�j�������'�|@�l��t��6���=�����Rه�T�`��Y$�e<�سՎC���j������#x��'��X�X8�x| .O._�7`�=�F*�CW!��$^��{ӦLl��J�x����ꚙ;{�C��~�H7T2�yM�X۝��0�5�` �
h�Z�I�\+�U��gDv97�χ,[��6�^CC����@L8�~��7v�)a�����Ѝ���]��aG���&��Xe��֋,�de츉����㮻�[�Ǡ��M����~o����a��Z��8���a�a�m��G��w�� �ׯGsS+r�������E����I���c�³Ͻ��ϛO�$7?��~�i�{�-h�0	���xM�6�ñ����7N8�0D���& ��ч�-�]���_	˵�^��,�>yl	׸��v�	��|%�z�3L�a�ӽ>��-�c�0]~��ذ���ӄ3=P��l�cZq�e���SNRF�:o����w�y��<�l�e<c��V�"�䢋d.��7Z3é�&���z��p�}���/���?��7x�Oi�;��������⨣�Bb0����.�/��R.�u$9�G8��
G����<�9'"F�Q����-w�w�D���B�4��3����8Lnl��/�����Z�u��̥��;�+�;�h�u��hmiju�'Hz���g��:�CD#5�9��/�=�M�}�����]�O��λ ��m����9���n{�c�;V�E�UZm��3��3���e���8唓��/c��/Uٟy�Yj��>���TK��JR�������}�y�4~����?�`P\��wݥ$�"N<�C~���>��%]x����>�#��vst��z�����VqLxND����Q,��#�T��3� ���Z�,��MSs����^~� �L�C��j�'���`�]v����Pk��{�*�ƦF�Srh�\{-jcu�s��e7���N�~�=���D
N�
�47#Tä%�k)������{�����_�z���p?:j���~�al}���b�+E��'��Фj���F�t�~��B2�!qLB�B��\6���0B�g!3��h��v�����){��l]I+))�q1f(�Ax�m�$tq�S��vk���^�����y睯�7��9������I�1cBa?Ǝmǝ������x"�b%�����o�/��>B�F�����[O��/?@��eh��!�R���#W�a�}�@cS���GQ){��&�={�m��/���Đ��e�����o��xb��1:fD&�a�Mn��Q[���d�g�<�L��`@�V�ʈ�q&���7!K��u����.F��)���#|�׺]�5�`���L���l�Ĵ�&�Q#i������B�A��=d�O��|��//A&]@sK�z���׬Y�M���Um�>��=!'�t���'�z�!�N��@Xo6_�z`��FC��w_�΍�q�_��_��dI�Z#�s�ʕ���Gt�W��h�0Q�?����
�{&O��_�}�����{�k�x��d���`�����|���D2-�/�'�g������U��k�k�&`uM�|�,�[�|^P	mx�-�2����}�]x�o�#��,�:�I%�����'���㌳���]�HW�4+��{셓N�.�w>�}�!f�+�r�-��˱b�J�����'W�M���<&����H�ǿ���U��;��c1<��o�[#Wz�u���_���<e���(���M��*�5�Κ`������7��<򈮱��&,��:q�x%��s"��Z,z&����w�q;���#B%��#���;��oH1����Q���nD(L���<�n���`o���8���p�a����$��^�Xm�L�N;�t����˓��3��Hg�"���kwW�F��͘�.���J4�����c�j�*%��;Y�9�sf���{����NS[�_�뮻_}�}�a��a\ӍZk�s4�ј)�2Iw���'����N���ի�tI���'�G��n�	Ͻ��Ө�@M�HX�F|�FԵ�c޼yX�z����5����d�`X�RI�#��?B!���V��o�����v��y!��7��;�:�4�q�Y�;w6�3���7` 1�`4� �6o@=�j5�k��^���_]�]@���My��7o����r�^�+��/�Q;o5��A��*X�b�z�\,��X�p���!^�%q#�D"7UIV*"����?� 
�%�fo�3�F1���4�Ƹ�$�3b��c(���A�QLؘ��´ڣ��U�.���L�l��ǵ��1�CKk"� �o6Y���_���S�c���ۡm��u�#x��Ռ�(�"�ɡ÷Ht�)A1�B|�-mM(yJ�{�\=��V�E_� ~��c���fN�����o�
b�P)��4ȝ��F�ۣ���T�y]��._R�rF{�e��V��v�8!4&2$�I������r���U79�E��v�AE2�9>���
ٰ�Ȥo�9�ဃ�Z�fr��V�Z�9sv�g��o�}��~�;��4b�$rL@X�Ujkk����^\p�<��Nx橧q�����g ���R�y�t�����C.ˤ��~�v�=w�9"��*L�in7^~�̟���혠Ġ���(ƕK�z��p޹��g���%%By=�p}��B��}�=̿�nMp]rΛk���wae��؀��n��V�U�4�	����S�Ҙqz#��uC)�:��4~q���������#�"�aVo7�p#�x�5Js�����Y\UD�A�s���z��Wp�������sq��7Hy����{.�lG����9>�@,�=�ޥj�n��{�Alͺ��?>�|�L�չ [��U8�FIa3�o�B�]&/&��g�U){Ƭ`�|���aA    IDAT�d �)����BV��$�H�>�TG+0�����"�9q تc5��<O��s�x2�1�:4y�� app@I��O�U��_-Z�9��F�����B����8��G��OW��>*V���]'ǆ�T4�-�S#�B��9�����瞣DH�5��� "Q\�]����c�-f��SNAc[�H�@wo
��y�Y!w�9M�-fl1L�n���y�x���%�hR6��A����ǟD#[z�f���FK������A>�Lv5�i�?a�����9"�×�l.�L����fD�x�m���TA�;�����?�p���<us�^�^�-��
��PE�����6F�/^v�i~�G��ܔ_x�AWtn��qe��h�1ܹ����~2�:����kW��B�`�� 	�20*�!�Ǻ	�f�Ae֧�>�"N����]�
!J\V��Ф�*7"V8T_#DC�O�i�Ce��rc1ښ�@�B�<��8N\���ٝĘ��U}�O4��rW���3$���߇/�;N�l,Z�-��X���ga������8���0���̚[B(f�Z���h�D�G�H+V}��fL�b�6�w�/=����	gwܱbt��*%T%�S��V̨��v��qR�g��
(f���drsC��TÜ� �E��(�u�2y4���B'�����mU��,,��J=c*K^V��;���)��� ���y�������y�჏?REqܱ�K$�k���]U���G6SD]}�O���6*�`b�����n;c���R榛o��u�- $��; ,/{B��>hd���,�l��LUkW���a2����z��eK��mhjVbJ�s����℟�����=�|�M��O����X��_=n��v��a��	H9J}⏠�z4DM�� 792�)�Bh�'
���h7N~M�pv�x|��Ֆ8��`�iSu})OJ=r.��j���G��$���}vY���h�����'�]V�o��.�|�v�����Y��[��0F���f�l�q1�S%�՚+l��|o/6�a�&0>���$5�����
�M���*q#H�%=�i�$��DG�Z^K"T\ol�����Z�Ye*�9+���E0��� &ut`�Y[+ rP'�g����:������D�Bʧr��z\r&;9�9��B����I�p�����>���S����՚�sӘq��'�<��&Z��8ɬ��qF��`´����#ͥR�gQ����	��:e�$�����Ŕ�[E>�x�O<��kX��ψ�(��&��#~���yCS�Ú��H�q^w>�|o�oYْ��D�R4�ud�rB��h�T���Q�،B�����I�k��&�ճ=H�h'S�4������-J�%mc�����H�r�+������ƈ����?��C��C��?��M��ŷn�F�W����x?��G�ذ�L���v�	�AB^,��c,Y�í����A{LΌRel��?�.T�D��<�(W��a�F�cg�lh�҇Q1�C��U��������Gg dχsߔ*�֘L�^���B�(����6�b �����p晧c�}vG6��"��� A��nMmV���|��x{}�@�˼���}��s`�у,�ׯ@���Z�y�w#	�eb+��5o��&�������}b��B��Y��*�{��C�����5r2n¬G'ALN�ڊ�& V��w���������ـΤ��Xo_��v����DD��3���0U+#n$k7tb����eW\��\�����><���[������;8� �������(�:8�w����T�1&f_-]�]w�7�|J�V~�u���]bR���ށw����t�\����$o��I4��q���T)0��܎���|�J���X�}l��dE����B<�VM�"Ι g�!V�LNm���FJ�r��C1Z�B}D*~1Y3��P�ؑO����.�3:�^�>��E���$��v�y��!)�5�6��B }Љb��N�1Ne�\D|���ԉ�G#����ᚘd��:�G<oLPf�3F:B@��Rl��(�y��׵���#�i��ӛW�TZ���u^A��G�5:����b���|� �2iͽS�_L8ҩ$~/B>/J�RH����=�� �<m���54�">d�I�9 �z�*����o����ͭm��J���d6����Q�3�"�w�t�i[U�%4�4��X&�6a���33�r>׍��d�\���L؆b��I��\{��sm)&#|ny���~M��g@�*���.)`˘Y�H���"BK�wmmz����$�F2L&��`��$�	��e.�����k���O�L�@
�0�c�ԢB)�*Gv����R���'��p��^6��W�ƅ�燾)��ۗ����߾y�����fox �ލh�	��b��5X��B�����a�|�T���c@���,�T�{�;{�4�}*�:3Rnb|(w�iw	�|��ڸ(���NK� Af��]���D8�s�n��ׯWe��n��K�yl􊩿�Uu�M�f�����QR�Y�𮜫�s��(EeL�F_ǜF1+PǬAE�`(buDAAAɠ�:wu�\��>Ͻ���������緦�N��s��g��3F�\^t�r&>3	��o��鑙gf����2���֖Vds�v��`(���6�����S�ByU���[�X=�p��T��΍kP�s;j
}�d��[Mh���Y�@YU�����M[PU\-�W�˂���ʬ��W^)��۷KbLs�$?D8d�Gs��b$\(
z��YY���uKP�M���,�Q!V i5�S��P�ҳgv���v����C�(�\+y�(���sC�n���>|��;P����L¾�ѭGw���ly�}�����{�AyM5�l�!!�""7�����ڂ�Ε8���ok�3NO0�'Ӗ���fl߱����Y��y|b
��Ĭ&�M�ga�f�9��u���!o��$���hW�J��HD"��T����	LH�^%�A�U&Gj���+�<X��R��.U�^]*+)���&<+�xRY��e0�8ؠZVr�RIq�(��� ��f�ʍ�'�����T-��N��RѩZz�<W���ě�>�Nx�� �����O��b�Z�E�j^���u��ZR�;߀C�Td��Z��8���)"
��<���l�H�!��qj�k�O~h�5+���[����n����:�x�*6*z=�y\�����Q �:�����seI	��؎Qw�.�w��7d�F8}�H���F�r�Nf�$�6Vk�&a�0�Ո��YZ-�0���;TTu�����6n�Od�r-qܖ\��%@�2U�P�}6���B�ع��`5#�PJw�	&���.<1��}"Y�Z>[R'���8��U�p�TB/4�I��8���I4�
9���	+r��)�."&CM��Br�(�w�}'�������ZɄU*sJq�dD�*��x&+d�	��w����N'��o�H�b6X@�Nzu0Yr�
�6����M.)v�y�Q_>���?���:a�%M��o}������̦X8�	��c7D�Ӂ�=���Ѝn]:�������>��
�o�A��0�k�; Ai͚ղ�8o�@��_*�(���5k���E(.)��"��(߸\�0y1q!�p�CvN�}�r�
V���V����ʜ�M��	��9t���_���u�֭�T����:U��*mTD�ѣ����._��m���Mm1X�>�.������!":�Vt�R���.�����+��r@��}p8�EN��R���^1�ڽ3>R���}�b�[A�k��O+�^YkY5���	P�D�F����7����ڦ��km3��oq�b%t*�4�mf����=���x*���G�>0��A&�9Q(Ŷ��� ����3N��͸������&�1�v����*� 8�O�D�����+䆲��Dc��<�駟��ƍ_�w�|�w.F�~��~|��gX�z-≌<��y�<�9n�YA%R���E
���u�	o�U0O$�&#�3����%�j^'>&[����r��+4j0�],�-I$��	(��LPc� N<�xL��4֬Z�@��p^��X
6�L�����!cC���:kjnD.�B׮���3�D(�GYq	\.nh&��j��ǅ?aۮ݈PX�S�w7۔~6{���+,+��b��-���D5�x��1"��qR��f�� r%�*h�X�e��.��M&	x�09f��%1�M&��Z��Җ���5�����1?]���Ɉt4&�H�r�_�Ty̅J��W��r��P3�҈�`���B��d�@*�ù�~�g&MƢ�K$���*���@%/��o�^�)8iDb�v��o�ŗ^�7�,{��I����V���F�[Z[b��ٓ�/|&'��ױ�b�
�,3|@��R�Z �M3��]+�9���ЭY��vl޼_�� ��j9�:�AT�栃�%�������y�R�I|x����;�1�S��It#$B�i)�h2f��;��qa��%�6}�W%���q��s����1��7�[j��?�!|�ŏ���3�w`��M�."�4bcv{d��B[i�
�Fc<R��W�G����Gu��?����4�/|��s�����Ę%K�0��@��F��t��B$D�NŢd�bE��Qy�� /������He+kQ��k��C��'��߈�bq�JĔ4'�M�#'���(2�xԢ�&�T��D �xnM-���c�j#tB~.�k����-d����E.���!r1@�18v:������ohjBUM�;�OqB��B��u�^+��>�G�/@�=�VR��ߏ.�:!�#�p���bB.m��-�ѹSg����O���Ǳ��M���T�=�
T�&��\�L�϶�G�����d@'�@f�5�+�	+�Q;ɮi�C�
�z�|��r�����!J�����BV\�LJ��b�>�b�<,	C�`�u�4���̄�((*���,)g��4۱u�L�4�T�{��ʁf$�2p� L��(�͙�pF\���g��H����>��~߈��'=0h����ˡ����*�����Q68�:�[f�|�6nES+�fKE�����v����3
���@��v�(��K@w�1c�`�Ͽ����Y�2Gx���F:ǝ�SHV��t#lV�f$"1�z�����-,*x�1����τ���1��X��6D����#��K��x���X��g�HFc 4Y�p��Mv�¢R�);-&a��s���շ���z���@-r�$�����V��a0P׌Ra$dO�Ya�Ո��h��¥��Ȏ��/o'Đc�>�ۛ�<���4�E{ޢ�~�1��� {�d)0a`¯�ݳ� ��ϝM����}�}�q���z�������
�χd� ��a{"����>���H��C��Z�r�1�閛����,���+���� %�̉��r�+a�"�ucB�c�*P��$�����G8�Z�����0�IgP��`*��#Zߜ�sIf�.�'t�M�	�ص��n�D��!.�D��җ��m/%}˖�=�P�2��c��WЧWOiW�@�~��w�h�W�iuM�>zG��b��M�E��\6�/�Pr?|�@ȔL
R����3$ձ�6}��X,�YL(�q�]�j������{�е#��9���yK��3�3q�����@�}*���a�ɱ��
M'���qK�T3]:w�{�o���H��[�n���ND�޽1u���R�G� ���ǐ!��7�Pu�	����K�%��0�͛�3�|:,&��̀��k��Dq�U�l�{���T:�����L�M�s��'�()*GkK�E�ƍ��Q4~!D��[ҒYd$H��Ml�"���A��̇�1��o��ݱ���G��;2� �LR�2��҈��q��a:�4����s��~���]Ke)���p���qy�ǫV
��33�Q*����-��Z�<�L\�y� ���N��\Nzp܄	���X9�������I��u��U��u|�T��6mQ:�F#�+	E�E�иUP =5	�m�w��^�|�c�C�r{� H��X,�ݛ7���n���'|���by_���C��G�տ��L~^�g�ر�XǠΊ[6T��`)�1y�d��{n"TA$�(��\��LN�[��3���N��H6���c������c��K�V�<��HL��*�[2��UR���/��o۴�Ņ����4,r��s�[���27T��r�|a��x��G�o����}�ek��^f��q��Ew{�5�b�u�Qx���q��c維(����X�R�AÈT�U>:�AT�i#���m����[��_�fB����渚�u�s�D���]7pQ2���~��^U�@�6[��Լ�)|����#u�?�x����0e�(��|4e���O(~�{q��:�� |:�M<��d,��GQn�uN��1�;r(ď^}�����*m0�4��QR��xy�����;4���a�b��q�W�3f�PZ�ڋ��B����kimy/����:�<�|�M�Z-t�����`�k/�ȁ]�f�&��� ��gϮX��
<���r<���b� #"�`NM�q�<��8Q�:�����0v�}���o0~�3���'�ƛGa�+�b��=�:<���@�$�8j�/o��`�%C��֯��;��K������_P�s�-{!���dBJ2G6-�5]��HrK"	�=!��T��dX�[�b��M0��0K5������� ,�$zv�"�?��A���C�=2�D�a����[	��}�T)�=2�Y�V�O���ի�JOH�۲j��	Ӹ5؆��r�	��?k�`k(���%No��óR �Dn�b��*��;F�d���eBʨ�銆�Z���ߍ���^]ˀdV�Y�X,GZK�dD���g�v��(
<.�t�	"ky��cdѬ�m:w���P��*=mr�QTUt�@��H%�+*�7yA|Vk�DN����EƱf��9Uޗ���ܢ>r(�V$R1e�B��*�q���J�	�0h�4��q�fAC�5�R��+&�-F�`v�ٯL/������i(�>jV�^�W_�)A��PDqx�9�؁��+���b�J�)�h�g�s�۳GTʸ��~��$��t�SH^�Py��� �r��W���A}}���yK�ə��g�M�l]�$u��-++�&�g��T|���7�h�*��d%���U���h\+O!�Zfv3��Ze�/	��
��&<�G
ʪ6Z+G�q��i�2�d0�^��TV��x�4&9�x�l.�J�#2Jp�3,ʳ�?p@�RV�F�G�@��u�P�9Hu��#��G��oxLt3&��Y��y �yN���ӂ:É��߫c!�����_O1���@>3���D`4��*�V4����ǈG��M��-*��N�r�6���lZ�S��ғ�#F:B$n�9@/2��=�e���)����T�@`�,å~ͨ��{@��;�׫'�M{\pY��n<�4�޻=/��u�lG?��S>o{�����%!Sȳ��������Ϣ�Uxc�L)*�|r4^���hH��",[��>�h��2-�%���
���sѹƂ��>'���O�[o|�M����'���Ȁ�x�_ ����HE:�^n%I\e@��c̽�=��
=o�?���ɂ��Yߙ���D��
a�Tz@'�����)	쪪��W*Au�D^�)�`eA#�H�!��W�ߖ/qy��h u����9ڣܡ��ӆ��ry,�	���mKNs�3a2�i�1�X�I�0���"D����*������q�kG�����uz@�}��s�dQչ�V+��B,]�3L�(
�Y�x~�*B"@9���B�Vd�Iࡁ̕W���m�D����N��%KЭ�])���+ǉI�҄��`K��엟����G��3�M�Ϡ볣��^��{�b��"ժ>�����LS�^`>-��:�NFaȶ�� h+���6l޴UHB�jh��\|�3�����-ҝ3    IDAT����莞}z�y�ĢE?a���6�!Ɏ$V��������S���[o�!�"� .@ѿU�r�}�9"{��/����wa�����DMu¡B~+)�R�=s�����X��
X�c2�$� Q��K���m�YhFyY�ҧeD>V�4�#\�ϴ�(��+.�"�pZ��=^��~�= ���)�u��x�Е��=��K�?���L�l�Br�H~"]�hW����
���f5e=��1p� ���[2�E�����Ѕ�G9������(�+Bc�!������m�=.�H~�z��W�vܱC/V}���^}�Yw͘Vz�PΦ���.�]��[o�Y���7I����H	k��?����IJ��⦼���1J��n�^d2��������ڗ{5����q}("�v�����gIN$�Q��*���9��&M�q�Y��
��i5�'�~{&�1^����ש�����W�܀�N]{��NR3�c�Ptk�3�i�Z�y�a�И2eF\+V�^%�"H]w�H� `+D�Y�E�|���$p��#1n�X�Lf�۳5U5"�L�I�nx�w0��Ũoj��������-Z`wR��%�,�}��ݷ=~�1=������������%���~�`���PҤ ��Ҋ=���@2s2%|"2��d�q�a�s�fV	8,�/5IROD��˓�I��p�$H� ��e3��0#l�!���`�ݻtF�.]E��b�Jy�I'"`���Pb��RU�^�N�%΀fѩ�
���^��4�p�fv���FS��Q8�?K!E�UxB�x=��$�-{6p����dî�}��ňN%N7��Ք瀣.-M�BZ�5�l�!	J���o~F6c��a�q��}{�J��&\�|2W�#
v(��A	���Q2Г��*��w΁��&�9��	 gV�}��%nP���Եyv{J�2`��j�	��}�w�`�Fn"&��8X�-;D��6Ie${�ǝ,��GA�V���u���.�u�����G�8^GD乡�3җ��>��>J�V��T��b��o��/��0�	Z�-��{�"����M�]��qg���q��n2�P��z��f7!Iy��QR^��H\�wY�q�Kgg+��V]����:K�9#;���	��2��'EN�6?����r�>5y_C�\��)��x�G�����u�b�Vw�~v]c�Rc��z0W�9���b��p�@�b� �^����)Qn�+��>��RB��AB����+�����+�\���\���u|=�됰���Z�$¥b�z]ٻ���w\+�QMĈ|i���F���)�v�|rM�\��9�V��au��6��f�%���l�B�Bg��`�oAe*�	2��9O�g>$�R�
�y�����&0xK��8���d�x��wa�"��D���Ηc���˃�k�GG ׯ=�s�qRH�Ҙ-Lx�2n6pP_��nR�6\t饘>�Q\|��v�+��jE#��BW�W��P�J����O���=�@K�$�N����|��s�EH���1�I�N����&98�`�"���m��	�W�w�B�.X�b �=%�����3���� �;��i$RQ؜!�p�����M����s�8�6V9��1��B-�~$��+$4�ۄ-	�!���SE1�uH'0n�K�a��D�`�O����~X�^b�a ��*/X2n��sL�}j��^=��B���b��&,Y�;,����i�;�7/>��&�ƤU\�f#�����6lZ��:W����ڴQL�8L�������Ń0X2����4�}�,��{1hБ"t� Lm�SO=U�^�?�x�צ�g�eC�f�IL��j$=d�����C�Ś5k��Ҭ����3�38����+aei�b�iO�%�"����ޗs�22����}&m@��������P��I���b����pD�>BZ����������1�c��-"
Dd2AŮ�9Oa��m���M6R�꘠:D8;vlÂ���A2+�t� ��)�3߷���l��hj��M�?G�����1F�F��;%m��3��5�VO4�qDjyٯf> �-d*S��� R1���|�Ck��x4����o���.!j^D87L�Srg�Q�GV����x�͌��0a⳨����r��`�{'Df�~�B�$�i�-2��k�h��\Y_Zw��_�r�G������WM揾������v��	)�~�������R�§�ȈV�3���>3I}Y�Hh?KI�L�xD:�MD�2E��v5EC�@Z3��%��2��1��&��kR�}
���W����l���b�F�S|�<H�=l_�tg�X�*�����i��v��`�I��p0$��:/�jQ
�C�ȕ��={�
���]��p��]
V���$�>ZZ�p�%�����}�>��֭W��Y3M��cP~�D�y�O�I��p��v���6�Ww������/>���Df�s�]�"ŵEn�g&/�o�1�'�U���'���o��~���C(89�V�����d��̉4i%2�,�/,��4b3`�đK�PRH�vV���.��}C�[�k��H�q,f�(�"��'b��,��ҋ��';��4���1��#���eK�a��[��19^@C�3�n(�j�{�#P[׊�M)|�p)���EK�dq�N��`\���3�YN���	=z�����l��ȍL̏P�.lߴNS��V2�ɚqZ��)x}�@Vmv�C�t��Xq�u��jie�d��Ѯ��
o�⢪���}0�f�ق`�N3��$(PC�����/��5{�ܰ)�I��[t�S)q}�ݻ��M�	a�gR��	�j�A	�d2��1�>�46�a���b���KQ1Z��B8��
Y�g�}6�=&�5]:c��/��N,��l��F�����*�(+QJEr���ǲ��l�:nqT���+��M��N���>YQ1��iim(>N_u�'���h6`�s�yV�Jz�&�6��(����|�uK5�m�z�T�&���Si+�\M���J1�@ ���[�%����YTuRc6���!���e�3DYq��n����	Q�4��C`m�R4�����"c�&ɯ�U&�����^������x�#�=��6}���?���5�#Y~���FoW����3��,=t�B�����g�eu��?�wF5Ä�;!r�yS�G,G.y,��*��pPo�#��bpf� 2�lOqM;�"�+�m�O�&����'�����ׯ�N��9��w��qˊ��\�����F��
Y����;�� �{b��{&�B��jl�X�>���2,�w/�x���(�����}Z�NA�d��� ���짓pM�����M#oļo����Γd�k3C�����Ԯ�`$!�:V��$CUE�ϟ��?�����#��[�R�'G��v���4v�L�L�dpr�$k��hȢ�"H�j��n�`���h�߇P[Z������U'��PRZ���߷#�#�B}c���]V���pYӸ�Α�ݥ
V�<�q�54I0j�b����n}}�������N4��.��@��M�6a���8��s����~�z�߼�di���v�n���huA�-C�fd@�~}eV;��c:�ӌ?;{U��v'�
�pYmpظиȹ��Dכ���?��PF?8[͌��[o%��r����1�%�Gf@��COr�D�b�@!m�ۜjs��v������F;K�+�s�w�2��8.z�Zd쭰P����)��S2}���O�@� /l{q�S�De��v���`��5(,)��rfѬtH2"٨���kkQRR�ʚj�r�ip� y�}�9V._%�"��J
K��uS��.@�bH�jm��b����d�t��gI'��}"Ra�}b� JկX��5�-��XْpE�Z#�Qe,��q�e��f7QA�}s�X���:�4-�g;��U����x��w��g��Ků(Eo�Ra�!��.-�!e`ʨ)7�t2�N��p�T�s�(I���#u8n��:�4r���r"���m��ǽ��e�I��*v��4�`{�նT=B�ˋ!z6�oA�h.ljF1u���H�������.�=h�o'r���v�@%i5�yt��LJb-�;=D����'�����Ev�P�f�RY�Y%-���oN��IU>
�p �cj�`�B��st���~����TA!N3�u۫y�ӳBm3�e�D�W�3Q�Cnz?^]�ڟ� }An�O��7�y��%I�c�b�A� �H�B��� a��чsd�"I\C��J�%9`��ҳvt�*�0%��2�D�n�L���1dfi�2��زڔ�+v��-ɅՖVZ>��[��).��r��ݯ/EP0,��("��(����Y؜�0����m���Vc
U�����O�QU^�݌�}��BIq�doNwj��ď?��W���x�&��?��Ѓh�NK
��y#���ːC��v�D!G��Y���R��7�ܰi@"�\�?�/2~����.CUU'\y���v��c�*l� �昏��A�탌P�*C�B�Zga���̥���#�G��V���H�|�~��F�-��B�Z7�b�0�.���jt:=���1����pDϮ�ׯ�lDtTc �Bf����_|Y��)P����iMK�
�0�2�s���B	SV��a�M}q. V��8���X�1��>|,��������i��V���˗K��ǋ0F&+��Mͭ8��3��Œe+P^Q���u�� ��mO�b�N�W�Ed:C���3���b���{�1�RUΈ6�_F��*�����8�F��H�gz�NDCmȤ���(�y�������L6��;w�kcS3.��JaǞHQ
7kB$�E(�F$�E��T�5r���B&1]R��B�~X�0��#<b�$�x���u�dCW��#i�퍑��g�=\P!�n�UA�q&^�I׉���K�}ܨ�����+زe��2U*n�<�zUO6�{�R��!;�UR(oq����LojEfbU��8��C���8�?���mD�a���y�_˃șH�u�9H�R���ɏϯ��" ����q&ˋ�`eg����ᶀ�;"=MA���0��y�Y�g��h���<	�T4۩�PcWV�<[/."���RY��V5����'&F����X�(�3h�8��>��(�Bu�q?"jĄ��u0�ywJ��4�����]$F%d�ݫ�AW���o�X5�����d�Җ��6#6���r���Q\Q�V &���bi_��������t����4��jCy�OPU�����a4�)ށ��뫖��<8=`��6�	6{&XYh���;o������mo����W��<�1�b$4%�e*!��)2l)@`�!&�͌h,�3N;�6�Fs�.T���e4��/=o�݆��V����G��.]�ɨ����f×_-��D'�-����X�z׭ע[� ��bƞm;�+X4���/��'r��Z`ߕ�U\��$��:K�۱c~��Y�ɧ���G�G�|�e�!�a���"�ؽ�Qrl���DF��*�nK���;���6�_��}{пGWd�!Lx�!T���7�E.���B,D/�r�$"� �;wF:�Ä	Ӱ|�j��2�B����ˬ�L�����(��~?�����3�s�ј����b'�̟��<���K�q0�_�Ą.7u2������XI��DV�엋���{�H�|y+5�{�������d��h_cs���*+����W\$�$���F��d:J�24-�U�7�2�3s���6�g�z��'p�E�#j��_~B�N�8f@o�a�P���yP}C�L&�����h�ư|�Z����e��S���ⷍۑ�R�Ć!��C��e�C�D���F��!��T�}k��$o�P�Q	q��<�h1V�!c��9Iz��o��e?�k�F8���1�r�"Ĺݼ�
��ꔛf�$՟�h����T� ���_Y���^5�=��`�����u� �� %^ڼ�7�uT ��J�H�V��k'�h�T\�X4#낆'|n�������)Т9)^uu�>:w��zcC���R�H!�E%�1�P˵�.�TR?���)�J�]�Z-��gUo����9N�Y)�"ֻV)�X�3�2[.�Q�ۻ�6طï�Z��K�_I�Q���)Xjxp_�0�n5�6��ɬ��q�@O1&�/&|&-�ƚ�d��ŉ�c��IBy&�N��|]�r�x�S��)T���D.Hf���*�l�/�&�<�t���hGa�8a���}������'�-M�.��0�mͨ��_� tLll	�ls#���c1�
|Bl�~���j� ����ӟ?qߨ�T��~���^�|�|r0m�LN���6��-�it�!�O	��a�
dRZZ�ݪ�j�"x=�؁������x�س}7��_��z��'�DG�]{��D�Z�x���W�,"�X՝�q�Eg��؅���8���h����y߉��?żￓ�]1%!��b��Ƌ�n�H�bu���uX�����S�Y��f�w�Mx|�$4���A�t�ȥ�h	$QX����L.��ݻ��a�.t)/Db�18�>��9̹R�8�VE$�̄�1�q���HήZ�U|��G7����F�P.H�c�ͺ�)��:��N������ggo<W|^p�_��	�=-o�ai]Ջ^�o�e�18ݾ� ��+M���4m���H��Ѳ�k�
'Y2g2��L��%�߉c��'�NT��(���
�g_�Lwyfd����H&�x�������b��eؾq-�z�nR!��k������D��m�0���I8��x�2�3�c�E�x��������K���͡�A*k��۵�s1jH1a�gkQR����K�G�h����-�K�V����{�j��7eK��{ꩳM���3��U����+^'_iP�x;$�j�� �X��5r�����v^��^+o4J�k����VsJ�_gb�s�;v�y�3HХGgt��� �{yO�L6�5�G�~Ҿ!���y#M-͂qm���?,X��z'8�s�&�<�ʋ�K&�ۦM���o�O�xh�
J�*���<G�Wt�&~%J�"�W�xL�v�����tNg�u������8��6���4ௗ_�G�w�������hll�k�[�.�l��1�&g�nv�dH�M���G��G	�lυ"ʭ�B[L�v��e��l6	�}�V�q~�����c�b�j�WT
�ɀ,�Q-��B�i
5e>���X�r�Ywn߉^��D�x�
6遷i5(b!et��У[5�Ly����y_�~y�1�\�/̘�ݍP$	�� �xNz�S���9;�6#�.$�����rT�������h~�����������;t.A���&�
��C�=;�x���+Hm�������j�҇ۢ���l.G<US����e6l�Y ����G��Ո��سk#��>=j�M��w�Х��p��nİ�@u�n�ֵ���b��a1��^�.Ł:��xa���oDYy!
]hl8 ��&����I�ɸ�Qj���PJ\<m�~�>�	�u{���ǟ��S�7�Fλ�z|��|���R��uBYe�o�Ũ*\�S1 2xP>��
�еg�������0�!� ��o���U#�X��[7�h	!�%��@�JPS�s�~�����j�X��x�oeE��>7� ǣ(#�(����	����U�1�TV���g�f5M��]���A�^���t�cp$�M����y�	=��w���NW��M/M���p��x�2x���FԄ`Cc��i�HX�fM��H$�2;��d�Lk�ht�*�},"� �Ŕ��\4
��	FC
/�xs��u�v-G[��"-�ߵ��u0��3�.}`c����w�ĵ�݀ؿ�'O=��5���J�T�Eߌ���jUc!�M3�����:z�P�k�l�K���GΤ�]J���v{G%�GTqv��M/���wi�R����$Dj{�gR�O�$�p�܏z~@��,w�{�׎Ϫ� ��
�    IDAT�Z��O��'�_7�%�^O�3YP=~����{�T�H!�����W^�T��$��)��Ѓ�bۦ=x�ŗн{�����_~�s�=7�4�
���y�F�wX�|)&=7A�1���v�B�{�E��2K��IO2�;�#3�<GD@F��;［}�L����W6����b����rd��'졛i������V�	t�ta֬���e"<w���هT�����^~�e<��XA��xc� n�����j�{�}�V�����J+0~�xIB����q��!x�GE#}݆�Ȥ28r�@�޳K��j���Ti�]y嵒hs��k�Wϕ����4C�ŴI���?�;ｏK�zn��j|��"�0}l&&L񔇀�G$ac[��{,�c8���x��{�{����̬�߆?����E(��BK���.�^�]0��z@x�Ϟ�kē����\.gmii)m����g�	��dʖ3�r�l�(Pu6�1fsY�ɘc�L�R`���`0�
L
L��%��Q�`0H=��l4��Y��`0�T��Y"Ɯ�d��r����Em4d�df�h�-Ƭ1g��2H�L֤��Ig�t�h̆f����_I�.�X��H�UH$9�,$|���P�q�����8
��8P��\e�^dA���v�B�*�Z�4e��D�F+r+*;��S�B,��[جN�a��+��h�^��[��&D@����y�5�y�8"Goa�0o�+��HX�rV%]:�`����~�B�4����
Wa	rV:YQ\�E���B��=0["�J�Y���]Y�����h��g�>8�gR� \��� R�zD��.+�VEeE58���GΔEQi�T���)�Zŗ�������c�b��~��$����䣹Y������r�� �6��3wme]!._z��E�:�G��)457H�A��A�Ǐ�#įk@KH{OM�ǝ�&��ٿ��3��p<���V���D�Ge��dBaI�l,���VW�9�E�p{KDĄ��J�2ԓYe����'�����:��X4 �x������3ѫ[9��C܏�][pp�6��A����x�Pt�= [��bź�H����ñu�~���Ǩ�y$���g�,$�f����T�7���Z���҇���w�E����fG��R�zC'*�뤳�:R�������Q�p<_�:������٨���ecmW*�搵9gn�H�Vh����^�h$@�g}̪�2Q�c�̵&�����mtc��?�-�t&�z-���q��K��k��b�R\}�p�I��D��W�ٳ�ºu[1r�H\t�%x|�}X�z&N|';�<t����<� �z�x����:���Jq�ॗ^�qO�q����Ǒ/©��#F�o�ï�_�_�G��?��X!Ͻ���X��7��+���Ir�������1B!{g`3�p�ȋq�e�`Ĉ�dΙ�>��lܰI^���Qַ�z=�vE�^=���˼y�b��0��'�3O����r!.��4<>�yѝ�:�t�UW]��F]���;va�ț0l�1�D�����8�����O�p�㏧���ǧ�~.��H�J�U��D�d�>�@6�*�W^~65'��f��[oφ��A0B��,$C&���ǠnH#� ����ȋ��|UU��E1m�t����.����C$�0�s2��ᄅ�j�Ǔ���ƍ�����2�\�Kcc�9�\t��f�hmk�F��X͔q�V�$mS�k���TJ��RRb�oH�(:��si��|��\
[9��`��*��j�q ���\&���r9B����ɔS�w&��L���X:i0d�\<�3��fOi0G��}������t*.��<��dNf�M*.9%�2�8�6����C�f[Q�u�����f�6Я� ��7�"�	���o��g����b	�n�{����v��E9d4�f
��`��hWI��
r�����N�xm��v�
��6ذ���o߉ʮ=��&f�c��Z��?M�06lڊ�nR�+�B�Q7=���F�~}�}�6�ڴC��Gs�~\;�|�pto�Z��D=�vñ������� �܃E��h����Ǉ~���\u�5�߷&O�(˦�����hK�[J�s�������+B~n
�P>�ߓ����^���:��MCg�r��<;�q���b�
�&�=��Ѯ񮋚0��F@O�=����N?��/��[`g?����^$kXŚ[�u���"�5c����9 �J�d�r����*i�HK<A2�D���d���	<;�)8l9�Z�3�����иw֯\
c<)�'E|��G?�������^��ႋ.��)/`Î����lK�5�BV�mN�8xS���Z��L�(V���-�� ��I©�i��.����L^��g�E��$	d�^;z�J�71?	��LM|>FGdt�@�l�b��+l���޵�����o�U镾^m�W��1�����T�yd,"-:�P��zE@T2����#�ಋ��#ݎSN:SLI�Uw���>�܏~������_�`�ʕ���1�7D��.^�u�{�TWU`��a���|�+��ާ`v`���ĥ_��S�J�9a��"#��	���z���G(*2`޼����޵g7���#�b1�r�(�i���J�w3�2�S��5��P��:���.#����X�t)}�q!��7�N��ŋQr�u����gr����xp�����[q�gࡇ@��V\��a��������㇟~��w�7� |�xf�$TTc�O��#q�������ba|�YC�ys�T�k֮��sM)λ�*͚;�d$P�e��&P�⤡CpϽ�c۶Zdf��d>��6;ij��鮐.������1�������'0�����\�����K1y�;x���`w� ���s�;^��4�����O��wۓ������G����͉d�M�7T��߿��c�.X���&�!d�[���΋ݦi5˚�c�7k}��_H�}����<)�g�#��� �|��D�*C.�d.��Y\���iM�l2Z�q
�$a �E��g��	�4�6ʖC��1���)�F%Ū0ɪ9ح��$;�&��U5�}�Zح9�z��ػ{�XV�y|�JřP�(�KbHڐ��aC<����lG4��N#�Zd����sϻ\r����L	[��!cs�h�I�NA���
TF�s�:��$�t���qA�f0Ӥ3RM�nؿwZԡ��N���0�^#��vl݀=;w�fs��p`��hh�ǱC�ŀ�G!��c�3S�r����_���V��̅Ւ��iA<BQ����Y�L.���FYT*���Һu��c+B�vd���P��bk�g���r�c����*�(���u�oz���ͪ��W$I5���@�sޅذq+~�e�xD��H.]����$XUUVK����$�sziGkR3�K5�frJ�M�A:�%�0��-�EC͸��K���{�~�,�u!:WÐ�`��-p[,8�O?��7�
���M�0�9�=�x�?��p�t��=�����$�[p�>U�ֵ�%���|�}j��DV1�����x�M�Ȅ�,M���t{�J�j���� �7��o���h���U�H��2vFAB�R0��<���7MGHn��?*��K�h't$.�S�zއMK�I�j`m{"�ӷԧRGQ��JC_c]�0�����ߖ�k/��qw��F}�47�้��=��oǔ)S����?��w���^������vI�g�V{�`�|y*����9�g�0�T|����������~D��/���w.��pD�ATWw�%�\�l*�׃��ǣ��#o�M����Ask�$���\|$�g��[��.�FY�_������L�w�y���xL�:�~��B�z��+/��3��/��w<���b�_�i��G���O��v>���0c��n�u~�m�=�"�~�a����+׊�Î]�eO�ҭ�#V�4����uמ����M��Jj5/�3A�k=�U�w�~�M}�~�N;��xd�=X�|7~l,,�E�3(�<V���7�`a@O��s�p�U��-Є���b�?`�ͣPѩ;f��6,�b��T���AV82&M5>#{�&x=��BGj�S������k���xޝ�֭�:��c4J�:u2��` gC�M�\������l~�>�ߥ3����;]�*�o�'��n�ڕZj�����􊀋Ȝ5Km�о0�D���ds�Q��b�"cȈ�i�>b��˙d�I�h ��C�M���6���A$�X��bdSc"U552��G%�ljhT��i�sr䌣b$�)X�)����!��~��4��B1F ����otq�9!��{�}8n�	��T������'���(��1��瀑#o��Ͽ���z��?u-(�j�a��qWf�MdE�z�xe�ص��E�ݽ��>���W# ���DĆ#S�,bZPXR(��?���}��8���T_2�/眉p�	+W���
hQUQ�-�0I]"&YIb8�F/u
�P��9��9#O(]�r��rI�����8�c��c�A �F�w��=�Y-)�]���(�r�Yg47��/����f��7��4�
YF�t�p��7f���"��Ը�M�v�>V��	�3K�����]*��2�>9G��~�k׬�$��IfV;�h�����VTv邱OO����������&$�l?ЊpΆHʀ� ecbY�kIU���ŀ�M�]1���@�<&"��$��ﮪy�*���,�Z�M���@��Ã�^w@���4	���G�u�\�:Sf�b`D�K�+UoY%��5�\ޟ�H(s�������e,��}QWS��{�9��9Y���m"��`N�]G8Ý=�	 n����ĵW]�;�{���h�_��/<x�m������{�0o�"�!���T\�X��w1
)*-�}�R������xﵩ=�9���k�v�J͚5�7lO�E�-��՝��؄W_~A _�fL��c������;v�r�҄DDO,v�ɳ��SX�X��I��߄�a��f�;�b拏������w?�I'ä��`׮}H%R�Z�ҥ��(�~�ilݼI��t��ڭ���1Q_�jn�y��46��qceͿ����9��}b�'���i31��O�6�����hT��-p�U�q�0��q�h47��B�zb""��).�ME����عe{�t���w��W�ʚ#�BT-����l!W�
���%`7�����G�E�ϊ]�w	Jx�u�1m������a� �2#�c+N�sRЌ�t����͵��>����/�ו#�G7����j��n�~�	'0��hh���Nl_ɇ
SZ�Ω�,����������`�d�Ԣ�F�A��P2�	�C|z�|]}��9�//3�t*	�9+���V��P��$����G����C^'���U3G��v�Y愔�]%h��Mm���(`��`�_�q�&�v�0�Dը�Y3<��
Z�27�d2&��j1�ي��Ѳ?��BaU��E��}��2�>e����}�>���0��4���w�>ralؼ����G}]#Q�M9d����ġ��
�M-H�S�(���5�����n�!����ؼ~�8�Q����Ԉ6��%"�p{AY��T�D ����W��O�.���sX��wh�7��4��)J����R6l�m܀�[7:�j���Dz{۶���m�$ �d8
00#g�D(����>��߰r�*�Ƙ$���v�2����l��&�~}��s׮x���d���DYE5��@��Y/�#V�v�ڔ#���MM~��̲Ͱ{\"�ʀ��{Ǆ�5h����+���	�`�� ���G��)ִ$h�/�e����T����TV���f:zܾ�ܱ�X�����`rc_]�⃞�	�Ey�V��\���4�y[M�L���Y��w{�� Gh6��6�59 �o�җ&s8d��=SdEޗA��HGi*�1/{��).$�l�׸�����d��=J��5q�CF�4��Z�L�<Mruj��)T ��^����r�c�ls���׀!��g����뮺UZQ�&?��4�S�N�ͥK���>��9��7����1��!G�;y��9X��b�1�EL~�E|��������"%�ǎ#&>D��zM��<j)"c�����^�ĩSJ�1���d.�UX
_i%��܇@(&�U���,�s�T>K�ĭO�N��ʃx��Y��/ѽ�ҋ^��rlۺB�ɤ�n;�mC�_|��S�G�^GH���cp�e���984;������z���z���{����8�Գ1���ū�qc]J*����s{\v���ǨQ��;��ŗ܋�`X�O��SRVH�5dHOF�ܓ�aЀ����U"�ZRV�@8��~�	��(��D.�V�Χ�z�e0����٭��o����QL��
~]��i'`�"��)e=�P�k��٦�;�VhO}���7�?�����h�����c��=ztw�Boij�9Y��%�j:d�����@����/��JZϘea����U����ǵg܇�[�p3i�����P�>f#�\U�v��Y��_�0��'�3���y��{��yce9��Y>�r1љ�J� ���q�1����>:�w�f��F�SV�&��V0#%n��=;��t�S&a����۽��i�ՠ�`v�R=��|)+YB�U�bwʪ�g�&�t�	'bǖ��E���e31��Sr�܀�.>&(<޸���L6�|=�5"���ݸ�ҋp�Y��Q_�_6����$N$������X�r�|n��>�@��U�{����-m"�Kz�|�ǳ���J`1ۅ%O�jqVsP!�.� ��#2��B�bB��_n.��2mQRR�E?.���DB��PLn�\��]�h��*L^2Y�8��\F��h *���L���!���V5ϛ��ew�u��B?r��7R�(��D�M�h��G�AZf�9���B��>�Z����>�����-n_	��bHՒ@0�>�W��.o�K�'R �w=���qk�l;����b�ʵ}�;/`J?�0Z\{@�E��J��-? K�A�J-����^���a ��}C>���t$3cz�e�rΥ"?L1N��3ٙ��5گ͓Am0��q��R���=c�W]~�0�O9�̚���_�ѣGc����`�7�����ʬW$�>���رc��f̘.�ٵ�\�!C�¬W�ቧ�⋯�G��.�.>�;˖-�:��];wb��c�ͷHK�a��Gd.��}�=�u���BFG�<
��0���\s�\?�nd��8I�A�
�:�Uh��5x��G����a�s�p�I��I�����˒2����V*�%�!\uť���+�w{n�u$�=�l�u��8x��]v���x�L�2	����w���oaƌix�������'�BH��D�C:B�ۊHK#��f8n����-%2HX�[`02�Vm�ЮSx~����͇�[��r��N�6,������ʂX���b%k�ŀ�L���Xk/^�w��7��0�w@�?�t�	�͇LΎXJC��;1�Dn�f%���~�9����xn���E@߳��X<vv����.$�75��R�ސ������zլK�x~�:�Ԣ����rxeߞ��A�|}3�zk�����3O.P4�(�Grr��(Ly%`�î��RĀ�h�g�'8:�+�y��y�8(�	sW����2�B~f�s����&<�������C G�P>,0�<Fc22DE8��2t��C�-���*���T~Ϫ�/��T:�N�R��a�Ӯq_P ���nij���ď-	U]9�F.����0s�t���A^Fs���t�Ba�/m�&/F4ڌ�b��c�q��/��y�e��z�)RC�9-5�����Y*�
y24��"F7#�Y^�l�H8$3����{q���Q
�;�<�̳X�|��鰹��}6_6�z]f��$�Ӆ�3�ND	�ťEb@��G1-"0C+^�>�.,ԏ&o1�� �Z�(�!H�W:)�?C$�����F�aeJԯ�`�i�bD2�Z��"n��HW�=    IDATm��6���3��SB-kIl�jTƹ�1�MD�+��ܮ����ɇZU�V��A�<��%�I�R��|&�|��~�(����?
 @@������s����K��������:�7p�������՚���䉣h:�szA\u�E��Y���?����p��+ѧOW�u�(-UʆL��~�)����ߋE�~��ٳq�	Cq�`����֛q�=���+���L��n������l:$tP��"M�WA@B 	IH�
��|���"/�HoR �l�}fvz���9��������u���3�����|���p߃���CmU5֬Y#�*v���p���2_�j�$�n�Gu���o�~ӇX�䧢 ��OaWK7�?�d|��cp��7��{@Xl�m�=�F>���jj<x�����Ã?��Pz�x֬~����8�cQqk4)�BcMyp	vo�y��G}~��2����p�7�9�)���s/8K�/�d慗���>�<��#���'��[0��WV��!�����4�\ ĕW\��?���Ft�"�|4;g�.��Tw[r�b�;��&�ݎ%�2R-���h ��'�x��N��}��!6���=��vҙ,�����	�buc��mX��>��a�^�D5�,�FEɴ�ܰYM(��<��+��l��T|j��i�ukk�_���g46YЇ1<8Α�2e�N����(?ز��� ^8;�ׂ�4���V���y�u��e&��	���_�C�����CS	~�d@	���?Y}1s����o�?�����W~��˷A�p��݀$���o_��X�t-v�t�ʟ,Bp<)R���Vl��(JS<Fc ���񣢪�hB�F�&��JM��9�L���양[�z��c$�S�дb�	�VϬ�.���Iǣ@�"� R�(c��م�xE䆓O+�T��i�Hз�����/����7��S|�qJK��M�bZ��r<B��x<�D���!�L��ȬD��"d3g�}��2ǯ��B$Go߀�}xn>��#�r՝������?DYeb�<�"����� ��{�\R����"�N����!+���~�ߥ�������y�y�mN����Q G������s*��DLdq�Q��!+�CFdCXD�*L9O��������%��B�5sV.~j��orO(ĩJS��Ő"��]��9ؼ�����򜸦���.�=u��_G�����L���O�ߩ�>&@�!����kc��7;x��2��s��%`(~����Y�� �>�{8����f��,ʋ�ر�w�Y���1<�QYIP,������o��9眃��:��f�����{ｇ��޷̃����O~�x��8ꨅd�b˖.���+�5.<�dYo￻�����r�J���=12�@e-qD@4�ƕf�i�0����p��������,`�F#�^/�)+kK��?Ɯ�M8��'`���Xqǝ������G����Rx� sodP��lx��c����������w,�3�}�?��;��y��p�%��C�-�\�3~x	����X��A����%0Y��h����ݽ��p>{x�~#��wҬ�M6d9�$��sY��8�̥1��^�]wo��5�#A���Ѡ�w�N��N��&��M�a3�ȣE&�@8Tx��v����W�;�7Iv���d\����䒖{��4�6ǟX�蒕�ͬ$R�?�2�ٳ�x<����F�=G��O��+�)�S�ISr�����������)]f:��w*L�ל|��^@��,蒨�j��::�N5!���O0f�Ȏ���忮�����ֵЩ7/�i�J֮��u�X�d%v��ĕ�ވ����,��.� yc��x\����$A���xJ���0 0��o�C{W��ѳb���7@^/��8�G�aʥ���Di:��ʗ��ҭV#\nb�����j1�߇��(J�|�4���!A�f��n����kǅ� ���W����h۳SE>;�`̛3[�<'o���(���pi�gnd�NDb�����ۄTb��(,��y��Ȭ�i�,��އx�ŗ�n0���O�ŗ^�k�_���zV�G69���e�E
�R�;��I�؆�H� >��%�L���{$)�E�r�>�bX�S �	G�u�Z�b�� ��6Sn�S�V����R"�+�:�J�ē���:�tx�ʗ��I�J��$�/7�V��*��)9ϮT֘h«/�H��e'�����$��NS��{wR��=�0��?v�u��wQ�˓|�����3�����kL�,���BP�唖����<YcT�ȗ~����WA=)\�\6!4�``�E~��gZ�1�`���l]�y�4���{��Ő��{��)|v}�G�%��μ9se}����]��P�d��W2_�]b�h�d�)��r�����)�>ܸ�%�"���k?�����Ȩ�������.{�{�O��WO����382���*	꼏�����`�|��u�m7`fs��>;;�Q[W��sg�ޗ�����?^{��;�����.�V�o�.��S��W]8��g����Uk��G�>���B�@�3��7���*X�,�LY��}������
v(��ؔI[���� ���݆ǆa��3�Q���h.g�'L&���
�\�	d���`���T�#ns��.]��zKKˇ�X�Й�Ͳ����D�� ]�VԘ��H:� ���D�8/K/̴�V~~П�`)����6�$ҝퟩ_�}⏅s:m�>ql:�o��ɜ�yxFk�k�'|Y����"c@Mf;���~�sC��`L�<	����3��@' .B�I�����{~.��ϖ���=�3�P�4{�)�"�OڴѨhw���vQ&gDQi�̂�v��4�X^^*X r�㩄T��tr�D&ØJ<b� An�r+�"�!#��7fNdeɣ'���9��|^���F�(��5<�Y�?gc�R��1��/���|��?|6S.��K.>���T�TɦTRR�g�{����}3Kل��N��xNcCg�v?�@��B�1��Rݏ�p�-K��`s�['���N���nv��5H�ZYN)�-3x%Vc{T��/לB<��Up:]���=j��x�>̙3OLr�{:�[�sU�'{",���8�lS��Rp9,��ME��y��Y�n�a�䧫���,,�Ɍy�P)Tp��k%p3=�|����{�<*���=d�U~@�V!?Y37!�_�ɞ�Zt�����׀���f����}d�x�!8Ӎ�&�]�y��~d�J�����il�?o7U�Vh~F���N"`8�9g�g���4(�e1g
�����$Y5fY#l���Թ��ޤ^:�#�~��PD��D���|&w^�[��o�T�\�Dcaٗd�a�B�N�E��Y$"C��d���+F��"������\'�K��I#��T2�`�˗/�1��3ϸ�hB@�I��"�E��BC�g�|��'q6��؈ te��䥤�N�GFP\R"	i_�0JKke�d69�=��qTW�c��Gr~��b<��_q��{coi���X2#@`%[K��E�lu0qm	x.��,��'���(�w����{'�a���#�sx$ �F�W���.,��ҹ$҆��&��X�Bq[b�/��%k>S@���� ��X/���C����T9�6#�/�3yb��t}��t}�<]�>����ӵ���Ѓ:߇7��-��)_�Y@��x�
k��sfi����)]���F ���5�Wݫ;���739lm�&ss�Пݢ4ƙ,���nTT���W
����n�H(���˹H�R�r�L�ZO$���jsIv�ty�ۛ|j~�|�a0`��~�����4b���@9�e�Y.7 ��D'��L&]��e�8MM�̞ǃA�1x�����>�wFPdw�����X�W_�3^|�Yu�<��i\}��غy=6�_���<ZZ�<�&��âEK�ߛ��tZ�Gav��Ӗ�1ڏow�w�7�}�f�l�@umJ�*0:8�b�[ 07޺&������n|��U�uÁ��\kOn�:Œ����##h�h�������):�D�}>��$ҟIA|Q&;�4f45�ɑI01�8����QRR���4�FG�#@����n7L+eؽ��@H��I]���K��
 (��u�	�ԫN��
gy��Z �gÓz�y�(yɲ̢��gvb�����\���!u�?.T����ǳ:�:z�!�-��OR\ճ�	������oD���?�	������&��'�	ڜ$9�,D�!�Yq��15��n��gBѰ�GV�|.�LΉ1�}����P��L���8�7	.D�TJ��"�qaE̚�,j����yf '����)ɄtoH���lV���G�n?1[�;M�Z~���@���� �ʘ�_r�Yx��-X����b7Kdq3A���U$���U�l��.�:�N�︮D���C
Z�s����	�]����7�aq�*�Ddl�� ��^R:�,�BA��`
�x^��%�J�_bbUR^! X&UL@D�Kc��Hg�ZXݯ�|-��,:쎚�&I��D�Y�����C��n����T%6ɐVn��63J<�a�5���7\���YUCA���������p8����Ad_o7z{':[�
]�"p/x����Rau�W��G���'���M������N�@e��,�K5�5�9;�B���;z��6; 9�r\X:<6�A?��	�i���((紲:�G���ڻPU]�e�WcOg/~|�b�E��d�N�8�fRB��-�e��l&E��H�Ehq�j�p�甦�ǩ�y�� "4�Q.Q��(�I>z� ŒɴBwGc���0
I��lM|����|�́Ɔ�ܶ] u�e�1�����o��|��w��q\t�ipZ2ؾ�c�t�"���N�bǆ142���y���χ��)�f��C=��h*��+/Ķ�`�֭8��+1c�<A��ba���X��?�g�����ۏ+�������j��kw�&:SY`�E�$�"7�;R����S @���nˉ%����>�O�D�c��P�l*�L"�+.� ��!��#�Ҵ���`�PUU�\&��*��f�R�z��!�O>ނ���Ϟ��p���;�e�IC�˯�
�����̽�l����&ɬ _Z���64�.�	H��k��"Ը���w�^�� �0A�¦|�e?��f^�o20�G}��!��J(��~�E�$�g�OJ�O�e&��O��}@�	�-ϣ��+iZ �������J�<x;��
��ː�m�x������I/z���M��yM�oV�l$�B�s�A�߫J,D7�Sd���/-u>��M�Yr��F]u Y�DGh耉�����������\��P삼�H2��S���I$])�a�w��( =�Ș��	 ~J@ ����8�Ig�x IB$ �����j �`t$���: B֠H�i"7�v�x�R�u����"�P�7IwM ������#��vo]���.�cÔDŔZs����߽9�ؑ5�Et�T�
����X@q>Ð�t�O/��3���{v�b��sf5+Q��>eqɶ
YRI�yk��T@獡f��ߪ��t�����Aaz���A�5_gF��������e����_tqD�8���3�3���N�.}��
�Wv�""�CTi�Yx'�h��7Hƺr�j���c��;��݇kn�}�䣇BqD�9��� �H���_^x^���=)����h@P��"ɛeF><2�<����b���:���ܓ����8S�$$r.aK��0^��1���&�J���2y�^Ax�=X�+QY^.����e���;��Q[U�K/� ������_���_;
�?�X����|�4|��@�+�$+%G`|C#1�^�k�۸%�37�OaC��N9�Kx��_b�M���nr&�\���it����۰d�ݒ]��k�q�.���	R9��2�w����,�l1��b@��186$��W,mC��:�KM�Q�/AmU��:���󢹾U�>�{�-�"ؼ�C�wc��hoۃ��J�ҝ;�^��8Y}�.ǹ|IY�Xƾ���p������}C�h�9��	á0��1<�v���em*�I���EU��Ċ�Kȵ@�M�&jГQR�����3y�'�Z�z_�B4y&KiZ��V�A#=�fկGLM�M�;�%��S��ǉrw^�}r�Rf.�Em{jkh6�F��|y�x{u �9�LV�z�N����,8~�XbdĕT����T�.�O��v��P����7���s!��{CY1�\��vI +���{�[t3$�;��dL��L�ŦU�ɘ��%xv��k���؁�6�ԅ�� ��^!�̊�=,�V#R&R��y-ɾ�DX|��G�?�(*)C[;U"�d_`T���}��Z,��#�+�٫�X�r����b;�V�#"�q(�.�{%��kQ�D����9�I%	H&X1��@f�8���"���ێB�h�F���Da3Z '�B1+�_Q	r�`x,��^{Y��Mx�Y�اS�`��6��}�kN>��������?�M}$+�ݑHd��z�m6�wP��<t�l�^�5q�*EҪJU�)��Ғ�K���^�8�h�s�`8��WPW�A�m$�$��F�#�-Ɖ��ip���� ή���
���`��2�d����]�
xx(sY�FSI%�~v��o��%�/G��n\|;Z:{14@��BYYF��BW!��Fo[��#�/q�f2��������~"���7�[��ãҬI���|c�̛�6���O����։Dڄ8�h&�lT3c`�"��u�����EÜ�]�w��DPSU��r2ֽ��y�y�?�g��u��ḯ~��̀хT(��H.�KfV�X��z?��`+��U���p���ߍ�N=g�b���q����~&��2!�%���ų�;���G�s�;�<����>'�=e�u���O;ܑQ�UTHbB�ζ������-���:�w��U�@/����:�d_�� ���@׮ݨk���C���������x��׉@C��-mF"w�0��*dS'��o`H��6R$hwK��|�	�p��wi���#H��m]�$�0Sh)�(����&���(�K\Z�f�(K�%���Y�v�u2�4;	S�L�%s,ԙ������y腵���>��*��;���,{�TYZ{@ъ'Z�:�]��*��l��e��)��y��菂\��%�%u�/9}��Qa�����Bz#�5�^v����p*-����G�6E^�\�),&8cKZ�,����@q�_��QM}M-�����P��)�$�e��Bc��ӂ��N��#�lI�yR�d�2�016��7��%����W$��4%�UIY#�6�����cTnc�Y��F���п������D"F(#�_d#��ɕ\P�����|�j��F�2f�'0�
�:�q�	��΢P|�Ԧ���� �{7�F��3&�K��]���Oy/p�ּt*yZ��>K���?��������uOKg$�c˝j^ݝ���i��$mG��j:5��r�[�����֭+�`_x����S*�O�p'v����.B�C�
��tV��4�F�s�l=hS�����W�\��9�礚,l��^��N���%���q����'�wcx���fg�(0����iT"�y,&�o1jd�C�2˝=�	W_y9����X�a3�}�����R\Z"-w�ϏM3�0�m��غe�T�g�����D�eg'R�����=0:
��)U��XP2pFI��*�eo�b�ǟ��2�jOa��Z\p�����Ʀuo���M8���j�U�]*�����2��$#Q�c<���ՏakK̾Dsid�Q3Aw�����c��MB߉$��j8 /}�cA1�i㒫�g�knX$�<�[�U�cp(��/�-JC�$�2�(.��[�C�P/�QU^-��H�G0@4DyE�����%��%EnT�zq��E8ha�Ԋm��H��Ea��D�_���ؙ    IDAT��<E�`�����6oCS]3^y�M��3�꺛P3�W�x7�۴Y�9���6ߕ�ȃ�b�Ō�͈8�A��dri��F- ,�e��*>���0ata��lA� �g�*\���������2��2����E+^�^4Mv�GMnj������f+�kJ��f�T%`�1J&�if��=1�)m��`���jUf����|�Hh	��10�؅�|7r&,J���_�{��ס�.i���qL��������\�];V�Ľp�a��=��K���q$]�#��!&��Z�do��K,C��O�E4>#Ì�B[��D�� ��I��2�*��L�4ͮR��D����<�Y\�:�@.�v"�cwFy菓j[/R5Ƅg�b�c�t�� ��er�@��HZ�B�adX��oLRx츤圱(����8lF�\(�&^q���L�mOkO4�f�Λ���M����E,т�F}��\�e[����X8/�[��',��I���8��7�{�O�����P��3������_���1�ǪW��f�М����7�.p����&7��i 4��P٩լ@d�%fPX�����X�b-�lۍP4�h� ��L�q�9�/߇t'��\�5�'�ܘA502��s���SO��p�x�e��0	`��e�Vy"�C�(���c����i���ƛhk��E^*���7`s� F� '_�S�X��<��E���ٽ~T�W����[���~	�S��#|�ѻx��ECM1N����ױ�f4�o���#�+A%�1�p�i��(E�`���*ה��Ȉ�<[7��1�/�����Sh#22
y�x�OXu�/��dpâ[���[�׿�
��H���7//r��l��D���B?��lF�����K�PS����Vt���n3�Ŏ�xC#�;\p9���rX��V~�$bAI�I����k��]J��a�*!�� ��{����dKk'>x�#\}�5x�����_���=��{���c��w	,n^�u(�C+P:e���O�@"��d��/�Bs�^���$�u�F9��*Uk^yˍXg��"F��/�����#�<��MEۏ�j�Oe���(3om��m���\��01��n	�&�3�M
�L��8�9�t݊��0�[�tdUM��-۷���	だ|��J	��ڵ���`�It�s��b��=������������EbِH�.!��׃#ʗ��R�v�����>����=R����bP2"�I���/A,�Fc�L��eL�:�d�8��Ǫ���Vu+�0����+!6mt�V�ĉJ������*�MmT3е�/�vβ�'oU��]��Q���*p���hז>_�{8���i3�;�K|ץQ�N���m[��絤@V^@�/�$^z�U���o�?�q����X�bfC� a�ZZ���G����k%���e�.f�SQ�������0hO���u�>�ԓ8�m��K��N7,��Bt�>kS-��V��������Mϖ;�pӓ�V� %S�����s' �-�TZܸ��45������-��h+�܍���D���5�Ջh��6� T��o�Ę�g9Ӓ�7#4��ax=N\v����ظ�-D8���
��/�(�pԀ�k۹瞏��-������g�Ǳ�}������څ�`�#!��qY�v��D�Z��͙>?���//-;���.�~�3�q�����_�6|�&̹�Kq�w��=;���|�f�=�P8,�F��_=�$^~y��fc 1���� ��N�����c@[�v|�����Î@��L8����ض��W�=��Hgr��k�3۱��{��X`��^��v��"��lj����<���;؃��T��av�Ld1�ر	u������Ǜ����b�o����K�KFQ]�Œ[�����O6}�d<���2�cA���S.#(�C=H�C�B����"���Ӌ��|O��+~���0ڰ�/bp<�g�w)F�H���Vi�Q�W\>�s��̥�rc+�3I�$�,5�ZYS��b��	��IȽ�MY��ȳ��93������mb����G���?EJV�vz�Qͻ'�5V�{��UE�7Mmo>�:O����c'>�x&��� s%�I���M���ĩ����=��C���o��{�����H���x�5�u��ߕ}�'���i�O��F�7/^���J�r�ɰ�lx��g���+��d�<���Dv�W�e���?���|��/�k_��M��⋘;o6.��r|���x�G��X��~���z�!	��l�����!46����h�1���7����loϐ|��'m�D2�h2%���t��Y��� R߼xW��V�[S5��뢮a ��D�,��:�wT�稧	 M�*�%X@�N�ܙJ�C�g���Oڜ&g�)�΀�'^G���`�P:XY	s���-��D\Y8-p�^p�����#�o����>C@ok�3���f5�:CǞ���v)�қ2i�QVk[�=��h��W�>�p��d�(� =Q�U��c�g\{m�|y���y�j]_�����ԍK�kz3�󜟴p#d�b������M����v�_�����G4���I���?f���}?���7�t��,]��l�	�ӍP,�`8�����qʿ�kb/�>���v��ȍͥp͏��Ք�G�^GY�_�7�����b�Q�u�r�a2CO%�ظif͚�o�M<���x�����
��P]ۈ��a�TT˼������XP�o���Dc}=��u���.�?��2<�����+/���`_Ο�#?w8�n"���Y�P�������_Q߸ 6'eN��ƀ�s[�������2��7۶��gIe�y7�;�����w	x,��7�$\���<��J���a48�1�ϖ~4���.X��g�i�E�X?�v����s���v��s7؈���6vb��+1:��@�,T�[P[��O���~��Dq���B<3!��!-ٺ�9n�O9��RHer=v��aw{;��4>�ъ�p�;�x�����Đ�R�#�h�s\�0X�1Y�YEiE9�t��qR�vҹ��I&�z"=FN~s~@��HM�G���(���<���8�N&�·�l_u0��
����̪����u��i��z^�����f��{�!�2������nE<B&G.5�1�C���x�Mh�o�s��x�g�����Vg�{��.�&�f��K����.�&�#��7� ����"��_=�{���K��_��[o���'ǃ.�����wq�=���G��f�a��S�²e�p�A����I'��o|�8\{��]}�2����FAu�X�k`��J!�����O=���l���a����0�l0Y�m/*��p`��A\
�-�3<��R�~0�8��@L�L��!��
��5L����\]��MD�	�$%뷶Fwd�J�)����@�k�Z�&��y�D[_:[2��}E~�����鶭��q�7b��n3����ۓ/��{����?,�)5��)��4CZ?��m�ϭ������QZr��I�
�-�T9�Z�2���������������wZ{D�č�_��U�^�7�r}���b���nZ��.��<`���@�D��~��;Ż�'�� ��ۖ�®�.�-���963^��(4�Vg�jNO��W��j88�˥�o|3�j����9��Q .����8q���������;����fs��_�:~���������m I�Uf��GeMbsXZ^+�K�ׯ��Ζ)�T�:��#�������̟��(�]�e@.��n������������͆�nA"�����M?FEe#�F/rE͊�vD�.��F;�u�p�!����Z�w��Ƃ!���߰sW\p��hUS���%��#x���b���`��%f��Ub4Bkk����W�T�ݝ�t�ݨ/���w��Z���*|�m'��$�6���#>EEi��q,��z�"��.Asc�(�uu����Fq�W�.�e�ȥU�r�F�%eU���ǟ^�+�>'���9�O��AIy^z��`G(�F,��Ȳ�J�t�|2Y��'sF,x�^��|y��_��ed�!����Km�z+Y�^����ҕ%����&7*Cf����u#�W�.���}Dp%\&��u\y* L�E]pm_��@Z���';�x>�G<���=.�y�Cc�:8��/��$I���"+۶����/�9�]�o|�زen_�s����ŋ�qӢ[1���x@0 LNibtӢ��%����o���n�M*��{N,�|�5�7����֭{g�y&�q�����o���QG��?�ֵbɒ%8�G�Η��gKnV�-?�U���~#�CR�74�c�����������֯߃[o���+���d�.1Iq�#'@��銽"�>B��LUe-jHr�M�+'[�23$#�L8�k�)��?ђ�<1%�jO�����ڿ�^� �dVM��1O!�?��J{��0��3��&r�f+v��[�W�-�����;��E��Rt�>���cl���QI
�RS�s��5	�*{��M�A��(���t%�}���Q�Ӯ�������ؼ���6ٺ�w*t�(�N�{�΀���$���'ש_:z]��K�	�(Z�:����r��n��wŲ��o����k�?<�ۗ��x,��[v������(�BA=b���qFC�
ߏ�r[tU�fX8>��#���Yi3��lݺJ�F9oN�\���R��8����Nъg�y-]�
�Ī���L( �:�V���Aye�������=�Yf�t9�b���A}C�.�?�K��.��߇��A��p3��&�w"�3Ȕ�T!���f��쎳2�,v���!���bDE)A!��H5�*�Z�Uu�B�۲�c̜9KW.��M���O �� � ϡ��ٜUU����S���DuC-�{:��@֊"���A5��G�������~�lʍ�x����$��~�r�	�;-�����,E"��`/r�Tq�DC�8�ω8�Ə�����3瀅͞�V���Q_:Fdl�cqG��G���3
���hͳ�I%΄���]�H�s�cq��IQ�N�k��D������H	��r�����|��)sJ��X�L� �]����g3���T,�^�M>6�瞧+��_���
#�~m_a�F0V�Ң�K�="��0|n�ԙ@
�dg��8픣� �	f͚�SN9��W(%E��Rd�0 �]^TTUJǏBBd@��c�={Z%ГN���$����;��܌ݻwK��䚂H\��,���;���@�
>���C)���� lٶFC�������EF{E%^|��TT�▛oā4�տ����A�������|�2��a�~H�(����rƔ�(�Z�02R�E���I�l��ڗ�K����?����?& 
�'�t�T9��ϻ_�������zr�{La�� Q��P��)����),c��`w�z{��h$Z:�j^fz:��:��r���K%���:E8����tA�7ߧ���u��^̧{����c�7���m2���B4���˾F\$�s��R��� i'mMF)%!����s�E��y�۔4��ދ�3g��.B Ŋ5w�.puMZ;�Ő���=�}��>�x�=�t����=����˦��-]R�8c#o�����gޑXT ��97��P^R��s��I�>	�>\���~W��:a�^r2���2������Dڐ4-�����͚�,� R刬��w�!����܃�y�q�~�l���Z�D���AOW� qi�
EdN�%��g	Gǅ׫@�،f�x�عy3b���y(.-C�h`g1�l,[~�oX��/�A�,����
�΄!iDU�)�ܹ�O�R�fԣg�_T�i�����2�စ�x�5x�Ý8��Ka��g-�P@�1�ӌ@hT ~t�c+��H����C��~\�OL�����`^o��s�80E�]EU�X�p:��J����fua�����ݭ8���PU]�?\��� ��J�����<�h��(�)5b�@���u�Q��M̘]H��_Mj�3�����������c���{�ڟV�K"A�����ǝ����TY�Y/鎨�i ;���t�R�qX�ߝK����v��i����.�h�w受����k���D{���!N�,��J�l��i����^T�7H��4be�b�׭+�eܒ#=�u���ՀT�����b�)A�F  #82c�6���h�s}��̎_80�,��w,Fq�>�}}](/+ �-�n�1����4n�����J�cg�IJ�z��:�	--�#��cX�k�?�?k����_/����d
%!_ݯl�Of��Z�n�G
mY	��t���Ǘ)��H��qW~�@�z��PNi{��#Q&h,�)�ˀ�wa�ؒ���n����\�G"��9�r�=ݝ����A���( �����{���{~ ��ZP��`6)B3�B�?����tp�X��D[��	SA-���w�_��M'm������b�,���:��c"3�) ���%���<=��p30�->�Bgv����vYz�
`X}��Xp��A8�@8��`�Xv��>1`���T:#�@W�c7��P:��
����e6OSf�l��O�3��'7s��D-���Y����IX�U@��|�P\^!҆��2+���JlٲE,MˋK�M�B.�@�?��K�-����ozC#�����4g���A4��V�LL�6�oFiD�)8=~q`�P��aE:F2D:JT��#A�<��֍3�q�yga��X�����q�I'
m���w��6oo��W..l}��ho��������>�����f����ؼyV��o�q���%�a��v+vc��"��p���
�6%�uv�M����?���/�k�1�x�pF�&���Q�+<6l�Wmm6m����Wpŕ'���`_��| �m��H0�ߏʚj�f#ð���iժ6T�5U�E������7�}rP��F��T�vz��L!HM��u��){�4-�B���C�O��s6��ڊ�"�D�[���n��8�a��(��R�Q\��8��y���/���/�x�W������K�Ĥ�A\��(�w���&����%I3�m.M{V.e��i3�1�k� 	�Q���>���n��LNx��h	�#��U�(FZ�����M6���a���fA2=R��Q�-.�.�Â��12[Mdǩ��'���afc�=�Pl��&�Й�
'R&�V/Bq�O����K��f�XJ���M��V�M�ϧp�՟&AϓE������$_b�O��%櫖��/q�DD$])L�;�R���\JzS��{c��&3b�4l.'2��=��!��]�\v�~�zgG���gϘ!���)Aqz���^��N˂�z~ �Za����.���n�V�X��1��6��
�{	�L���0?�`pQ�2�t=y�[���A�ռ�].�V�3�s>�z͝�oj�m�ݎ���Y��?�K����x,	i~��?c��vx���"�L�)�!3��u���a	���E:�_��RHb4�j����mu�T�J�����w��L�Gt(�Q���q+´9������7K�PUY#���۷K˽����~�-);���q��s.:^�19S�f��~rdH��&�&Y)�p������٨�DB��"4W����<l{���q���A��3�/@�5kV��j10�DY�����ᗏ<wQ*���?0���N9�L,���;8���4�V�l�Ԅ��m"��g����D.�椃UV���p
c��x�s&ID���j�Ɔ�E]e� �,V,���C������}�ňfrŐ����UP���ED6�K�QWW�u��3�2.��+� 7�_��O���g(�Á�g�����(r��R0�-�t]4�.'ia�:�6L]�y� �[P��'V�t]�O��-�k��a_��	O
�c��f��&��>@	�P��,-^��P�)� ��7�a!$��hj,���]����C	    IDATr���pݍ7�QD������U�:'���PU,I��(�lp!â*��I�ب���}�
��B��� ,T�L'��!�4���aDyQ�p��������qI�����G`x5啈�"(� ;@Ŀ��H4�p��36�	آ)�H�-�K����ݽ���Q���L�G�6#��8V-_���=c�����2I)���-#q�N8�Ƈ�6���W6Ѕr�oզ�w@�N�T�;���Y�Q�ۨ0��)�]O���:�ru����lZ���o��uK�=�j�i�葁,�>
]�Q�u��3��r��k>mM��ϝ9Sް��K�	Х]�g��lW��p�h[k�i=P�2a����8诧'�����ga@�[��զK&?}@�B�u:� �^���L���B{w4�G]�@�����bfϛ�E�����V�Ɖ'��=-mBWk��?~���غm\n���7�5IqM�
�����M'��l�ǈ�0�RF��w@:p��-��t����B�<��:Ϲ�d�������f̚��Ʉ�6n@qI�t������J2�-S6�C�n8��&�u�
̘Y�Ì���P�+�t�Ņ��0\���	ꛮsV����F�0:Ё�
?R��-��T���t��Z�r�t'�g-���*|�l�@�3ذy�l�No�j�����!��B�-m�r���QY�C:BO+f7��[�<^6:���>�w��G��)��D*�ёA�w���Fp��9�+8����qZ�{�v$�a1a�;�+*����a�;
��m���_�Ë�9�ɚHd�5�����s�((���(F���q�'c��Yx��W��� �c`((	�����}l<�d&�����j�]���ѓ
�扁�i�� �����9]�0]`���	�^�~C��K@�����	�EU��["�f&S����lFGaȍ#���,ĉ�>�>؆���eؼnd�����pc��Vn��3)]�B�����+�D��"!�Op%�iV~�>��J���͌D,	��#��$�ŕ~	�0To�;)[A&ƶ�_�L�H\�E�S�}. �_-o�F4@<Ĝ�j���p!gReq����vi��·������*���㿂��!�GeU=�yg+�Y$�%��y��KDP]�G,2�-O���"U
���u���D~�s��LOk	���y%x|2��.�����\�,:ZQ[]�`8"V���#px}ԬE2@��<T�<����<������ƢѲ9�3���:ۜҬ�P8O%@������醆"��0��7|~��n�N;�GJ.ǣ���}��ra�0]����&P���p�
[�zR�":y�o��rg@ׅv�q+)Ľ��]����~���;w.���zq�Z�b����}�Nq٪���Ǟ��P��g�:`��%[d+���l���ՌD<�X,*z�ۃ���	��Xn"CYW���w�Q��:_v��ԅw�WT�`p\9���
n���ۃ�۷	r�-���&lܸ�X%�b�C63��y
~x���ϼ�U+V�������&��Y��Y�q�ܵB�K�i���4�I�h+��eN�q���\+��L�����A��p�mK��ւw�~'�t���ݾb��������ꤓZ���в�C��������Sغu3��n�~�f��x���\u�%(�o��w�{F��1<:�d��̓ʪZ�@C�aDB#�2(�8�}�7�d�=�l߹MF]�_�?:���=l۲w�� �a����G��B<kE&m�)g��dAy���0�s���n�shl�D��Ũ���[�9&�Ǥ�PI�4-�f��g�.��4���zkjbC����^�.'��0����|��,4�oT��&Ļ0���H�#�W��n,
�)�/u�z�hmہ��~�HE�u��3H�#�z�v/2t�E$�LdMp�|H�`�FL�\h�dC��G���cQX�v`��%��{"���[�Xʎ(�}��(4�b� ʊ<0��hiEY��e����>w�t �~;F���[�p��p� J�������d"!�q	��.X-NX�6�搵1>>�!���j<��2�>����꾇Q;�`�u��g�� 9�����Z����DuF�=����V�Ч��v�ˀ���<~�.��x2�'`U{�X��a�tvvc۶v�%��`��T�@2D��4\�3<v�kWQ��_;��#�q	�T����?t��.��b�i���
��WY`�b�;�O���2�Me}��<M��	�{�Ч��'�n�?��z� F�{���A}�
�`P*����f��D,�Df�e`e,$�h`=!�`f�R��\�Ɔ����,��e����~��[��ze���'%P��i�9��!���x��~h���83���H�NKQI�܂��<�	�:?�B�:"TyP�����h� ��V\N���00�F���� ��ڊH$���/�����Ѫn�kD`�����8�ԯ��'�ǣ=�Ӎ"��s0��������k�G[�y�$SX=&��U��`u�����Aس!�,Q�x�������#0(��-���������OY�����������QQ]/nv�~��7ϕ꿬�C#A�ٳG���ڦ@�e�hj�����p�����*�!��oŶ���3 _Y���5;������`6d�Y�=	%n+�6����εw�Ï>����Å�1
-�W�|,~��3��N8��;���.������F2���lGh, ��P4(�T2d�L���[��	8�~T�TKEHs�h*�Պ%;i~�5��i-�lʹ��P���v��-�b>̀�0��+�+���<pӔ_�c�^8��7#~��~m����\����9;M�`Jq������p�e���5 �Ջp<%l	v������p�y����cD��O�+�\:%�W��x3��$Ey�G�p#cx��אM��r?d�|4����>AG��X3
�l�B�=N��j�Jq��Gb˶=ؼ��Sh���Q�,I8����`�&1���rZ{;PQ[-1 Kb��[04�If�6d�4��!
�_�F`l�� �^}!������{�P6s!�b�gu�h`L���y�X#uUu�g��diR�i��(� ���'p�̲w@�������1��?��2�b@0�Ï<����D����V�YTzMC�̓w�t��cfy�s�Ԏ�ցH$R>�y�h��vu���>
s��B��˅G�m�;$S6v����1I*5�u�9ӫ\��r��յq��+���A�z��E{�^���S,L��婖|a�N�d=���K��Ø��sQ'�U����t�Й�3��~� ��ε$[��1d�}�2����K�ζܬ�`��;��;(�.f�Kf��̴���;���{���e-L��j��3(z�R�b�(Bt~R�LJ`��.�`�c��"��������1z��L()/sf�;��s��c�$U|ow�8?��L]9~z˥ؾ�cܽ�>X�@�׉��eTU��5,�
�=��lVvnn����r�2��~8KkeF���
k.�*g
Mv\rΩ�AWo��er=����5�?�4�\�6w)��b<���x藏�W^Cw� f��8�؊K+14��O�����H�AyY����Cc8��q�E磨x�����__DGW��o'(�e4#M��ɜ�ِBtt���Z̮�D:�J��BGw�T?��M��8��3qꩧ�����Tg^x9~r�����8�H����0[�nX�6���H��(&����G�>cr�/.Eum��Q���]��Qh��$H4���$�J��c@��xO�dN�'~�����%�}������#��{ײY���&��n���D8�� �)��f�ᚫ/�ko����&�q`0 v6��� ���<�u�A�G�kߋu�섿�V�,l��\��v�2��@,���8	g�u�?p���b�ͨ*+���n��Y^���.���a 	_0�j���Z|Ӊt�P�3��;nGC�o�ۉ[��9��2e��� B��X0.9�8�&���p����(J}N9��>�,^��ۂ��mș�p��"�DÖ���,9�W�����mm�8�B}�XlH���n�=��3v�精Hi���?���l��ּ���׸u}�"��,��O��"	3��|�+G�g�N��d�?��'���F�3�	d�f8\@��%���\w���-��������6����E���93�Eű��C���YL�lZ�̜ܵ:(�����t��km6�5�}ѫ�R�s> n�ٶv����'|U����#��s���~�t���Pt+"��C� 9Уt>�p��[�M��e/H�^�+��]w�#F	��X) �e�W��3����6�X���Pܶ�)4Α��[�j�A��*z�ج�q�N��P1�-~rVu�<7�X"��.��R�kR�2'R�	D�������3[��c��ې���Q��X��C$I|��3QY]��KoGmE	���jսx���a~s�:p6f6�"0ڎ�Z�ƙs�[�������bëo|�Ǟ�<�s�n�h0�����I,l����
�����+P��(��ln����O�����k���W����G���PT\_i��#�J**�Vq׮]p���٪����с�xN�V�	���`��DC�����@Dw���kA1��p[�/}�4W�bݛ����H��������b��{��]�W�^Z��;���-B<gF<c��Y�h(�����[0	�WL|R��D`��`5��M��D\�u�ף��Ҥ) �P״�[֯���=?�O�?ETF_SӭV�r.�h��z��ݾ��{��U�5'�^�ۊT.���*f����c��٧�￉7^-�}�Y����1�
�,86*x��p_s���~(��X�y�R�sfA�+c��������O<fpǊ��/�G�5+!���y=�g�~ių��[Q�Sp8|V9�.��b�Y��m�#̙�b7�[?��'|?���:�ʻ|0�@��O��B�z���5��\+��1l^RE�����)��-��nEY�+�>�W�\�݃A��1�3�O��������{Quf����:�)�=��-wpY�Xu�r�/�؆���=v��A6��f� c7��%;�;��i�}a��K��ѿ����ܝm��H���y�н(n�m-�dKs4������{�GU�_�gz��$�$$!��DT�4ETĵ��Et]i*"� MA�뮍��bY]{Y
�tBBz�dz�;�����M&C@��>���;��$S��{���)�s�I��K)�I�l��-_&8�zo��7`O��i#J/��4�l��]3?� =���*�e���'�!�%w��HrTS�jE��E�G#�n@��H,�u�6p6�n�F4���G���+�Dcc�zW�?+W��?@*m"��|w!Wq��}&�	��^�N	R�H��M�ݒ�<����ԯ�.�����eD���\�Eq�2�o�^��h���¼��1g�=C,˗���W\�I�Fa�Mw@YV�>�O=�4>��SLs&�^o�Q�Q�#�#���@&�	--�h�;�Ƃ˶�+a."�6p��Y58oT?\0q$~�r;f�xr��y�-A�$����ÅO��[���%�Ϻ���O>�W�C	��Wr�Mֲy}
��q��!��,3
��p{�J�:���)]w���>��I��t���f��!qjWt�K�I��ÿ�S=r(NR���~�DB�:�>�5ܽ/�K��iU�4��	P����B0,�Gi��>ۍ�<�;�-Q�6��Ck��(u��o���k�1���{J�R�Yv��ŭ4�{�c���MD.���K$�*��X��ϸ�
Ģ�����C�H�����H*�����F!G�;n����ڽ˞�_�1��H2��&*ZE��;pӕ��."�^~�]lٴM��eK��Yn-�*0���8\oG )g!��;���>��x����G1��{�Y���e������w݊�B%�������=l�k2�p޹S�G��仮�����s�����-�ɀ��'M�,֯�/��������C+W��l0:�~�Yl�B�Z)x3��|I�/���_2���Df>Q��{��\Y�RE��vM�7p��OWM<������Z���t�5�ބN�-��\p��m����_@]V_W�����A��_I)Ψ��� �2=ڜX�6�ўH'�`3��3�@�D�M�� k(syiٴL�$H�2��2�'�䟙�S��VD\���3ĠFԱ��B]֩��q�<�?9�I��b�B<�DZ! \��Q��n��8��+[�j5.��R�`(�¾��܋��29�iY\�"�n��I܅Z �j�m�M�ZL().�^������,�:�>��&P��*���70���f�)C���F[���	0BB{��5�i�J��/�>|������w��˯�j@|���8k�̟�w;�U�b���X��9|���8uH%��y��zL;w��A2
Jp�fgۚ� �n����EF�����>�]�]�|��Dȁ�O�'�5� �`��ulf����U�U�nFX �Yxj�Z���1f3]k2!�H�����u����	��;�,,CzD"�G<* �p ,t�󒜯�!1Q����ѠV�
Y9��b��3�����~����Xݯ4�6|�HL�8G���ٿ�]^1bZ=(Mو�Ԝѩe$�#�p��Rw��$�g� �$�ĘM��M�h6�b�B�ס��f�+2�!�3i��|2Z��e2=mi}u��S�N]�/�
��5�IjMc�Z��	I�������@'M_���$���Mjc2ER��d�i@2�ǀ�|�x�.������+�G�%�A�0�.s���A�@�^���7�<� p�ʭ�z���6DJ�C�t74��Q�QDݍ�s�Ř=k&"q੧_��W����������	������_;1��U�*��H_>QA�I@�oǘ*6��:�n��߻��h.=�2���W��!&�Ć'�g�a8�1d�塽�&�W\:sf�@,L�Y�m�a��'`+�(�I�Q�I����:}K��ˮ_���Л��+��[�.���XJo���tz��t�N�q����ɒ���)"�]��M�D�('<�:e�\�`��)���D�̇ !#ZtrP�T�#�E�/K���2�x��S'~�E�:����*�ׇ��~$�������5�)CgY��Ǖ�H$�j�RD�t0L<H>�$�����t@��v���`��Х�zɮײJ/d��@��4hP@�sI-ХC��"U8T�Þ��e�%A�ޛ2t�5��c0]�v=f^�.�R?��b�x�yT=ƀn0�pɝJj$D�7�����9T+�~�T�-.DQ������{ly9\��x�K�NTR�c�Q&���F6S�>8e�����ݎ�س�rm��tyYg��ۜ�N��z&�����%Ky����_��	��W'{�ڬ��z�#x��W�ƶw0c�d�?�*�cGb�Y,F>�2�F�Bn���@�k�z�[�~W#ƞ3{A�Z��3��'��3�p޴�%e��jTj8�+�hmw�׃�X��)&�,\�?�ڇ���	��Mo�*�����v���(3UM����lKs�2RfgM	�bԫggq��#�۳�f�4:�$�aZM���\R���|x;���@~~��zǏ?c��8��s����Ͽ��������X�#.�")�@� ��$���hqh���缘e�x�J	�Q��7R	��
���Hֵ
�����!@�l���R�go�ԺN���k�M�7 =�ω���@�u�N\j��)���O�~�&��0�ģ����$�A% ��@�4r?�T#�5#B�k4�`Pu�`��[q�%cY
������Ĵpj�XE2ƣ�4NU����m��d@��W���oc�����F�    IDATj�=����Y��������{x�շ�קn7Un̬�v7cL?�ܰ�m�(�,\�Vw :�
g�:w;j���x�ٗ�g�!�9�IY��N4�J�/��?]~�u-X�z=�r-K�&�O����0�Qf\4g��O?�}��,xBIˡ�R\D)X'�L������6C��7���N�k��˔=����)C6n�v�F���e	
�Ķ	UZDyJ��l)���*���68���]��Vm�|��׍�g�_@]VW{�6	�3�+�m�h��M:-~1��a���͞�3��)�5�3{�|�"���8 O���L��N.-�~l��袦ow'���_н�ܽ^79:I&�&C.u)9\*�� ��H���UZ�H���D�%@�,wӦM�E?��J�}l�&\|�Ũ�o�����r6n~5���h�f���#=�2��Ak�r6A)꓏��=#�E��ÿ���Q� N�d�Շa0��5���(��[o�ls��=(�S�n��g�yYV�9���;a�ڸ�M�1���F�u?m�)�ⲙ���/�駟�����x
Kʰ`�=��b4�
7��������p�Ё�~�iPiSF��j"�b�uR��D2Y]�+V����(��1�jjp��(�X�����T���ƃ�񆫡����j��je����mB�?ށ^~�7�9wރ�u����K\q(�[��9�&KJ���^SS�R�b/EE}������ I�KQ�B�@G?�2O!)�Kiܓ���b��m�B+Gñ#�}����(��a��2(�A<�����O8�b]m���/�����C44wb�%u��hsT�lD�*��"�F���/�(k�� ��#��D��m����qۈ�)�A�d�C�6�����a��p�A�cf�����z��uo�������MR�S��uU{�Y�>m:�}w���Ԩn4RI��4
JY4�!̺Ꮨ4n8���?��k��f니@��dU?%��B��Q) h?�f��K��������Z��yl�+��;ۮj���Q�q5�����m7����_�'&M�U���x̏���D�zx����V���V�T6�\�9��7bˆ�V���aν+�F�|� V��g��$�;���A�^�ɤr�1h��G:�z��5{a� �n^�A��yk]��ox�o��f!S��w� t�$�m:l}b����?�c�҇�	u6|�(dL>�l��o�� ���lћ��� =u��%����xO��zk鮐*�]2�	:6v%�B�Ji�ӱ��H��Y��tU�
�h�$K¨�;����cb�=sn|��3��y��� ?��`0XQY^
�R�%�NG;�)[$@��RJ�WtQ�>E�Ie!��h~]��t<�'�� :o@� :l���J�����%���t�n��}���]:�� ����[��w3�8 ��,W�F�7	L,�(��	зn��e���{���M��`��騫k�>yAi%6o}�$�p��PX|������p���CNf]x>Ə;{�@����K>��C�ڲ��D�;��31d�=�2?���x�8r���� r�������C�3�d��@��X�c�3iΙt�s���mo���DXH���}���3�	��Ͽbђ����?�oQ>���<r �Y���q�Ö[$��&����҆o���ǐil0�!$ı��_P�m���}p��3�j=��J1���,A�T���`1YP�Њ5k���_��5Yq�Ms������L�{J��Y��pP��ɀNeg�ٌ�%E�{�hlh`{"��"��5!Vhh�FRU$�2=���F�������f8-;;1c��<v�]��p�d���G2 ����z|�ٗ��m@I�R�޽qhpʈ����o���ԚX��2&Y�n%�PV���"�!;�T	b�^�Vk�J��B���]�:��+=�'��@��/����R����ĥ:tFF}�ƙ���~i6�H�=�r���Ǘ��.`�����q��6�2(h� y"���������fϾn� �܈pB��B�#�lә��@��q+�f��'���+7�˝5H��Y�UA����R�t�	���F�~ݹ�s�Y-�ɧ^���eQO^>�D��	�`�������1o���hr�( ���g0b�#��Q)���1�ehh���8OmY�«�(���u8x�j]6"19\n,��q�T����h8��\<+��������֗�Oh!ȍP�����Ѩ~�W_~.�z.>�������F�cZDH
��-���O�X��RI��@<5����o ���z��6YU��C��&���/��XT`C���j�����6A�{�����3=1m��O�;��w�9d͍MG�^oUyi_i�o`@'~�F��{~:��F��]K��Q�@O��{~�x��G���/-n.����<-��'�\��i���^KJ�1M�g�.V�Ks��X���RP#)�q����h��ޗ�xt��U�U���h[[��>�h7mzS�NE]]���`Ӗg����%w.Qh����\�f��d:���̸p��ݻv��LO,$ CU�>��#6:�2*�.��3���S�?O���fg�׶����
t��Tht���+�Ɔ:hT2�^����@�xw��8��ojGG���y��_���aÆux���0r�i�8�q�m7A)�#ۢ��jCnn6�Z5�T��'_Bc���B����g��*�Vc̨��y��}�P���(ַ����C���^}m;�F<�8n�s'<��x�@��L�l"NB�ρ��`W+t�>/))���BC]=��Ձ4�'�/��O6� }{$��i���PX������F~���c0�b��=�0�T�}*�+6mz��(���x��ٽ�5r�(45{�Ta�-�WH � �P�I���doLǡ��"t<��V�b�Cո��,Vң�>�T�� ��$Lٹ(�S$������+�t����`lMJ�{�+ǡ�z[+m$�7�@?n.S;6����ޒ+Z�:�������~�iyj�S�GF)R�t���J3.>�'����/����r��Is�� ���'d�a@u�������'pϊ'���G!� .(��6G���՜���	�<����i�u�e�
��ϼ��^ygO���� UH���{X�P\�Q�W^��������'C�߉S������S����ݽ�͸��Kqˬ����m�=w��>�> �E�Z�N���<�^d��}(˒a��E�,�Am��Vn��c�)��h�֝V�m��ހ{n�GV㻟B�U�� ��1Ϥ{�(�t�ѭF:[�f^���2t2��q]O x z�wAI��p��#;��Ż+]�C4��pJb8�i$HvW��j�h�	��"ɨ�`y�KW�<����i�-P��6�r���J��i�wvv:�y�Ğ�FQ
�=�|����������	��� ݮN�Q���z�EM�$PtԻ���Hg���@��� ��\�w��G�T�L?G,L�*��S������S�ƍ`-Z� K�N�J�N����#���-hhjE0D�*�E'@'���i&>˨G(��
�3q�W��p��!^�������ݷ9��`447aƌ(�[�2�MMM�8m$>��44��_�a<s�ԙ�ao�Sº��Ъ�W^|��6\�Nl��V�Z��'�/3���a�~X���x���O�C�%����bn�f&��k�b��p"�õ���W?`��_Agȅ�Z �5�H������\0kRU�R�d�J��dCs���؅^|zC�r-�{=�z~�u O>�W�\~���6������Zf���MIY)���c��hL��و���մ�+䐫U�F.���`w�����hzY�O��cD#W��hf�`AA�
������a�)��/�ѿ��-�*S6���G�4d��R�E4D�VtJ$����H<��n���TZ"�Q_���z�{&���ʣC*�}K�XC���I��w��e��n@Lw7K��'��*`�c����{��%)�����U�ʄ���QB�vh��S.C$D:�9����Cr�FY�F�Ȍ ��C����\{�X��������EH��P� L�R��)l�!��|�tܞ"�=��x��w0y�Yx��;�j�p�q�M�pތ�1���8K�U+�?�FvA	܎������^�D{g��]���,]p;��}&tz�������>�L��PRo(�N��R��\�I�A�>܁܁�'�d��������!��BR�[5�0��\9�\̺�bVV\��o����0V�
C��}8�f'�J��Lm��@O 3m�NTz��H��)`�Z6��d��HU�T0�n�����;j!�~O���w	���,��ju�ta���p2��k3�:�O��v͸��'uY[K���5� �X�T>tt�����i*�^�)����������鯣�'��+��zzf.����Yz梕2�t�$��	�	�K�={��$@:*��Sɝ���$?N�<Z����Kb�����D��6l`�Ѕsƾy�t*	?�n܌�ѬE��2P��;�;��F
i	!H��Nv��Sأy�)���7߰������M�\ޥ쁾y#�;�<�nյ57n<�=�\,\�Fc6b1-��f't�l^����r���� �2�-���'�����]��=�M��8x�j�Vk���3n�}n�����>��0�2	��ɀ>�����C�j�񵼾P�(ӷTe��

�ߟʜ��� �Њ���Z��ÆrvNi5�m����:�S/�\|	�}�]|����d�p�J�W^Zv����������a��@�橅��	� �R2����YYL�:ഷ�(ۂ9�_��e��+$����S�hw�B��1�^xѥ��������~��#N�w?��_k�P�y�T��,�J���@w�@řTv.�
P� �jS&��E����`B��N�	�
�e��4��Pٓ�����b��@�C�}K~����a�� =x-g~�����ث���{'=I��-CgƳ��yLE,E���q�%S�G|����&@fb�aʰ�=jzS ��A���x,<��B���k�1#)Ƞ���U�4��iB�[p�u�Y2�g��k����'��#�q!���V�u�<��I�\�(F�*E��=Ҍ{? �1.WN��æ�k�S�`��߱�,�?���������;k�۠4��	B����
ǡ1[ B�:`��q�W��K&s��`����=H�r!ǃv�x~w#f_wf_}��}�m����`�; m.R�;��I�3z��=��>���� ����Y�V��y3�@/Kpqi��q1PY��QI�B %d�� )uz]�$���Yّ�z���A7LfR�	:y�Pi���?^rλ�L�t"P�}���,:	w��a�����i�b'�ԁw��J�]'1UF>��O�[��0�H�͟���{$�~4���:�R��=2�a������;�iK��=��h��	��%@�2t��+��tp�B��d�t�9�H@��r��ЉQ�`�B�-[�Ĕ)S��؈`$��Fa��'9C�I�t����EF2e\ԯ1�T�����߯�mG��=������XL�����e��%e��ɓ�{�U�u��!���[��9��1�M�t���+�N����Ŀd�<2�j����
�N7�Y9�n��X�n�K����e;���Z\w�5x�����_"7ۂ�l��D�~��Vtf+	P"&�����Ʀ6D#q6�!�ɢ�"�6�#)D ��V���`2PTR���b�9p����.�y!���b<�ʧ�n�^44��D��k`��V��q����}��rrPVV��N;���Fɠ1���q�T�J�fH5dG��%y��<⅐��\�L�A�yj��a<�������ŗ�a���<��r�1���嗷�pun�k>�<�?�=��>��������@EJd)�?*���:1�S���MA;�����`9,����
�\�R���)� {:%���R��(�?��>�@Y
����R��2ei-�t@z�p<��\�G9?5b��}M���É�ܵ����GC�� uᜳG�M1>��7x�ב_4��I;;;�'/ ���Z��7�W�����g����|�s5��B���*��Z#�SN[�*���w]7�͚�p�J�oa�ko���j�HF��N7�]��M�0dV�z���O�{�?����������+�Rh�r'0w��_<��b"B�������v"��ADm�;�JCR���2 ��<��tI���;oƵ���퀻�<��~ڋ�1�9�o�e1�T1��m����E�xy�vdT�T@��sɝ`O2CI��.m�b�L�,�8�@� t�B�Y�MH���{tK���_tg��hI��ě����ZꕓV��x���IP���P�~�Q�˸�G�>Z�
��ɫJ�

�
e:U"lQ�(�<5s�ď��:���;e��].�����Uj����l4���Դ�w��)2�Qz�4n{��Otr3���O����[�uc&�w_��%q��J�3����7EL�\}7�J�T�R�K��M?~J &8:���N�!D4� )#4�\ɤ�?1ł��Q�G���7���P	e�/��"����K9C���&�w�y��N'��67=ɮ_�(1�I���SEP&"�B!�A����U2���j(胎��#��u����'I�r�]�@cc�r��	��h�� :m��QA�Z�t[�B�ml��Io��	�q�_�b�x�F�=�ݿ�ǒ��2�\OQ=�tJ��ڱd��첱����o����=S�P�(G�l�ՙ`��g5��C���gRPBY��ӎ���0�P*D�<���O>�a!�������&`�O`���v��	Ag&�=��啕��=��O����ep�;�o�Y��S�]ͳ㴰�J-�����e�Db�S���w�����\b��;�v �DA�����v�Yf#&L:��8��Κ�Ͽ��}ϭy�x��� l�i}���k�-m"�F"\gl��K|t>�8��?=>��i��]�EE(�[�j��$�DYy%
ۜN���DT���^�F��a����"=З~�k�:)���W�V"?nCNӖ��������/��%�FI���MLT�3z|#f0'��h�ryX���X�:����݊���9�ס�B�/��B�F����8�X�1���X~�-8w�p.8ݺh����e���,��� :��m�Yr,p����g�?Mg����/��2�O9�,�3���'oi�b��e��h���uW_�+.�M,�E�.Gm�QY�z�J������Ýw.��Ӆ;f݄���hxx��뫟��)A�/�@"�>�q��qD�HF�(���U�w\{�s)[�'^|���9TfT�,>w�ܦQD�gUcѼ9�'�Xr�*�ߐ)�ڝ~�D'������SfN"g�j���=�Y.A�j"�2%��j��T�H��P"gʻH"&te���/��K���m�R�_�{�{�S���b�L
Yy�erR�"LeeK$>�8�^А!U��F�l�"w�Tf{�֫/��%��j2WY�W��p9� ���	3i~S8&E>��%���i�z�z�t�w%��^/���~ף7�
0���(��S ^������qd�T���uq�����$����a�˵�$������q8�r��щ��P�j���ي+yl���Vr��f(C�q�UCGaӓϡ���Yޑh���3��ˉX�z5��I�6�0L:-{%�tC^8�L�,'����.
��X��]��YL�� �C.�"	�@Q	�ʣ��y<�����$��ƎŨ������m�e��ƺkQз�A���p��'��O����vq��7|�y���\�`$��:���D狎��=�>��'\�"�W�
MM�(�,By�b�+x�p��YLf׎}H��Ƃ,��e�*���@u�&��\iy_t��PW}�'���b>F��=0
��.[�&j�BIrI@E@���y���    IDAT4���r��3GV�O���!�6u���-D�+S�{U,�@ݱfx�~9u,�^Q��ф
�( ����c>�0�m9<�J��emO ��xz!p�H�L`+,DEi9�;G��Ɂd�T)��p"AJ��T�Z)B������^R?>� $@ۿ���u�;�čD��"��u�b]��޳�v�j����'�n��Ԩr�kˇ�@,�^��>�RU�]��|[�0BPٮ�Q�F�3�Ѱ�z�Vu�C?��%�%�a@�m���#��V��@#�r@.пuĔ�#�cΕSq��?�<��g���7^���c��w�����-s�CSP���M(�ec�?�E<�kG5�;���r X[Oe��p9}X4o.�6�+��ݿ��"�� ���N@��!�LB�e���I%�6�6hǒ��b��c+{�}�#T�|�I�*�^'Gg�1̙u��z
r��}���Ͼ�	_X[Q)�^g��d,�"@G�be���I�Mjuvf��q�$��Eh���HZ+�1$"��`Q�]L���O�t���]�ϓK�dQ���Ci��+��
a9�`�NbU"���~��oB|��L	jhQR�R$!���f5�C�XE~���g�����t$}�t��{t1C��
;��:R�������xd�,���'[șs������{���� ����ل���̢�u�.Ni�N�СCy����)3���w�8%���yӐ���T
���[�d�#�T-�������G��ax��֚�%_�
�j��K��?��t����q�V�z�aoŀA�Qٿ5�� DE5
6h�z��a���e ����u6��#�BLYmʑm˅��bB�
��pۆ� :/�˖-�N�ŭ�͆�bf���L��1�H8��c�b֬[X@� =�"`���W�RS�V��M�A���A��2�7B  �|)��Td������ޤ��oo���A���#�P{�	��(��/z��Gj���3e�%hjoB{S+�Id�����h��`� �#M@�1"!W���'�y1+�McaDC>X�jX�J(�Xt2��*�5B؃�?z��%0�/F�>FC6���ر�0L}*`+�B �`/����I�����E#mP����r��tp넀�*�y��Z���ˉ��T�U0�{�$�ByY%z[����g��{�S�ڞe�̪��z��e��K����e��u������ғ�L@W��f����!K���D�m����Gmu�GRk�ʘ��[�h�J��$̪��{����p�ecMw,܈ow�@a*�r7��i�P� �j9<!�v̹l
�r�5�����]�I�f�|�c@c��@{���\1���,�YGz���O�K�SOm�Ũ��6f͹����o�W]>�P/�������f$�Ehs9���LM$^?�z%1?�a�Y��X���%/���v��}�Jy���V�a�Ʊ���,����Q}��e�p��Q貌�"�69���b
�>S��UHC���H�+�ⴄ$�"��������}z4E-R���38���CH~O��
�8�)�/���x�� �,��Ŷ#4�%a�|(Y��F�I�IA���a�6�~2�V�(���3&�y��!G%\$@?�r��ؚF�Ie�\���:G=I#]7v/cc]o�aF"��Ǣ��#OF�c���Yo���X;I{.�c�{�1p0�*�H?O�� ����P��H:m��Sˀ����$���Q���3�$Rm�LY�;������	�	�h�6�Տ<�I�&u��S�ĺ�O�X}�L%W+�^:	�Ļ �z:��B��׈G��`(�3ƌ�i��¿��ovr��M,
�QUU�.<����_}�7�ڎ�%�������D���J���:�.4�43��rr��g�O;QP����c��x`��8p� L�,�N�0:O!yy�1����{��'�REX�R�������Л�ܞ��ж4��@�J�t��*-���@Y?��J��<X��V�`�+�R�摰���քl��M$P֯
�k�r�C�]R^������$�A����.O'�Y��ݝ�uf.���������䘴�9ې�������$���#x��W��ן��Wͭ�u��xƥ�e�>���-�9B�7Ι�۟@\��^o`�{5�'jąA/�9�^8(�\�)����DU������N�aEy���!���3��w�k�����{Coy� ��8��=+l��2J�'Ҕ��u� �~�&%�cߑڀS~���C�Q����f%.�h
n��,����kq��АY�A*@���Ick&Mr�/����g-���7����LZ���.
z�*Ba/,�:k0������K�2�����m�aʔ	xxᝐ'��� ���0�7{Pз����4�}����ic��xOl\����0��'��沪�E��;n�%�wo5�-�
CZ|*r=�wCB�Th*֤�C���UE<�f2 5�aܹt5�u�6�"M@.#��T2Ǝ��B^}u�0 ��B���R�˞ꡋz��� A&r7h?��#�J��˙����oj�M�����2F��w��9
�s�I�������Hz��H�EM��ʉM	3��EVQ�T��+BD�$LoPS!�bitj�=mG�5�y�/x�3Gp�.kmi=�v����,>��C���9�D�R�ɢ��u2@���vj�u��N��dn�ϬpQ&��+�K�I���9�Ө�F�`$�~��$@/p�6��n��%'�|�H�]����3H�_�gM� ��7F���5�Gm]#�1����$0�L0�K%w*�R�O�N�:�@�G��Ղh"���8���?����b��>�VCҠI�2�6_|�-�����7;��[�FY3��"'?N���@���ΎN��١R)0j����=�y�N��������r/�)(R囘JMZr�K��)�ڢ �2v��&~��a�{����T%!�6)�V�A I�8p�K�4�U[[���vTTB��{>�P�F"$�b0è1�y$@��{:���Ir�յ0�T0h���2�hVAc�����5�uZ��-�e��R��dQ�2yVf]{%��J�Yx������<G����w��y�.�'��_����z{�e�=��Ί@��g,�,�=N#"�l�V��)+��
�.����OQ&��3������+˺K�t�++@�R��N;�}!.m���w�)��33�㞗��@�V�i�n�7��,I�q3��T�~��Cڨ����	�]�DX#=��fM���8�?`��hq���*��N�¤(����$��f�9�2\:cr2���^��!,y8X�s��C�Hn��G�ߌ����1����_���>Ą�n�]�͂�n�m!:=4�<�ChU$L�#+`���:]�=��ȳ�⫟��z��p�Ŏ��"<�a,�=�������
C	��<�H�0�۠V$���!ڱ�?�O�Oca����-6>�:��FZ�:�*�'��+����`� �Gl�����8�.���O�&:g��Z�*�KS
]���E��'k{0O��R7���r{ﺮ"�����=�����R�'��'��K$�ۅMRA6*�S�]p���].�Y ,�M��4��5P�E�p,��H�D¢+��޹����6yP���ٟX������p�J�bϨ{δ7POϐ��d�G�������4.m ����ͧ�>����%�
.��&sȜSty��M�1��M�z@QBI�(U�5�{��D�Q�U�G�$S2����'�w�W�����7s�N����`�)�q�N,w���C8�1�7YM�wR�����o�1�#}��}ƙ��_���V�?{�e�95L�z�%cȲq����)����0f�$47�ؕ̒��@$��%�ܜ.@onmጹ���{�>��ofևW���@<'��M(dP&V9�����3� �&bəҵ�s�E�c�e����ft8�,��ϥ����{��Ͷ�׽{ѷ���l�=_ ���? [q1*����EI��HV�w��	�I��b2�����:�;Q`���%�(��2 ��w�ԮAC�;2q5�r���桠 .�N�䱵���9�&�16��:��䖍�>r��Yju8Z}��*�t�-�q�.�����*��}cNL�Ű;��*g1��!�uO�-���<Z(�T�SZ�{�2}�٘��������GeE�������~��3t�K��P����@��+<M�!}}�����=}h�g�c�ǵ�zW�9.CO�ȏKZ����h&��z�B���
S&���ώ�~�2�	�z"q�i"�%��,��{q��2�^q#�J`��-�g���&-S;G��sNj�$��;0q�@<��[��jBs���~�ڏ�FŖ�K������=KW�S0� 1r�tp:�b���1��0(����0�Ԑ�u�[݊����W���ubŊ�8wBg�_~��Y�T�P��$ࣖ���{x��p�ð�/s�o���V���څ8i�'T�^'������:���x���ﯿ�%2U���g@'bz2����	D�Tɽk���L�$P�*	�Y@��.�KIi�q��R=�ަ6�@�!:u�2��!h�~O�$�$�Jrģ')��C�:&ѵ��hI�S "|N�z-sdHjת#.��X^����}��������:�K`����E<�d�Sp�9����!���h;]�%3��(���3��Ř��9Dס�1a3/}S!v8�*O=�Ԕ]�h��-�3[tl7�'}&���1HߏFŨgM~� X&f��6>��'�������j�?�M-���gq��Ir�2�͠��ba�����>*�ʹ�*W%1h�@��LM)]�#��ʫ����Gka4��h~�e?>���逭 V[�{sK������h�I&c�9����;��H�9�wt �l�Ɋ��� IP�B^G��_G�LU�kL�6L(�l�yL�#�o���Q��Z�����F�{��CaA~~�a�,p!ۚ}V6L�\^,u���KB-#���kU%Z;�8r���L��g�����a���TU���B>���7�x�k�q�������$�T1�S$����Ձ�Ç��FT�7j(���R�c���*j�\ڧL�ig���?��n�����a)(BvQ��AD�c���uG[=Ə���xZ����ÇH\O��N%ٳ�sU-\��N�N=�(R�����=FՓ��dk��>I3�Gf�}ҍ!��Le����22����I�4�^K)ٝ��h�[,&t�5���ZnDp������������ǟ�����"�w�F���I+�^��u�QY�"��Ͻ�7���O5V���C��69n�u5.9,�2�������
Z\v�w:֭�Ң!o��k��X���Z�Y������c�㖫q��AMx�"	�و���}��*�TU�ɍ@����������w�Ƽ����A��}s,���?a��R�H]�Տ�,^�V_�K�P�9��qR�Q���P���|�ï((��'�?��L��REr�"�s����	�{��}p���`�UJ��EuQ1G�k�%E�t�'��c�V?�CN��R
q"�t��%Y������!�I&X1N����&��2�#
@g�!(��Ǒ���I�s�z.�G"�=�]��Gd����N����4j5g�T"�"�;}a���.5�3Pv�K{��3K޿U��D.z[��Z�d.��T&e��������a���w�t�4wiF<R�yt���>l�0vA-�ƢK�KX������`1�)?)�F٤�So� ��������Ú5k1~�xVc�c�7x�n،�6V�"�O��G�%;�������̉4
���z=>/2
&Dt��N{'3��(�J�
Y��J�������.d�f!@'�pKN.�������o�R�4x��!Gii9�;4���F3�F.�R�H�
�$SjM��>�4�E �'�M�{Q-ɟE�c2Z����A�fn�����Z�=��/��m�|H��F���m>�tؽ>��٥�*�`6�aЛ8.�_���6���V�a^ ����ʱ�#(̲�E�s����n��8md.�ﯾ<����5����GLH@�v��9�{{3Z�-��8�(��b�F��	!���4�RA�nG��.��F=��
m.t�\Qw��ZeW-��ò�����O�_��t[���^V�+..d@w:���GyY���
��3t�`[;�LJ�+��.��/���@ti=���ho����`Kz�,��������/m�'�O�������ra_�f3Z�b��p��3з��/k��`��J��7d�א����VŵWLōW��)�#������_���`Igkv.��Y���'�̑zc<��쾧�펝p}�q�y�o��e��r���YP�� ���FV�
�P;��8�,_���'��ر�+{u~�s�q��E����Oa�����?�;�?D�dl�jx=.�����Ŕ�C�j�q�;����Ga�h��xZC�UB��_��)�/;¡Í�h���r`wRk��-�h,��"��\tq!�,�������K�.fPi3���,F#��k���')���i�9����%�TI��uQN���������zb� :�e,F��"���
c�g�&ID�7D|�h"��,4G��6�M�<��#���֣���C�g ?Fnk�vd[h$H�ĩT,$���/��*��VbO�߳��Kf�,�Oϒ����XZ����x����2�Y2��S����3��,�ʻ����\Q�S*�M��6����h&��QI]��d�JB2�]֭���~�̙8z��G�D@v7k��V���P��)�����}���L&��!��ea�&��Z���No.t5�r4j9:���\��8�Yrm�h��@Ss3
K�"/�g[{��+**��k����:v��r:N�@�D`Ӫ�io,+��׽n��F�j:V��f�\�m���k֬�޽�Y�n�ʕ���od��k��O?�4��7oތ7�|���v�3�|L�6/m{���{��u���2e3�R����/�:Zp�� T%
rsP^^���j4=���,���k��T��7=��mа�0����?{�T��d̂���〤$E�W5���B0�T�:��9��~�P&H��,%8r��QA��Ag�g3W0��dB@"������ 4k�Hb���q�h���M�!1t�)���4�Ú��R� �ny<d"�n�Icq,�K�:��յfL��6�=_���|��x���M�ܻ���7�4�{��;�>?��G��Ϧ�P
�eI@!6���OHBU���ɭKA�K�<�}�k�j�c+��?�Z5��5��P+b0�#�w�M8gt?�\qdg+���P��e����9�@(H�/��}������c'��5���{��-��f�CXf�B���W�2�L�a��~L<c8V?p#�V|��.,\�&[9:]AX�t���xx�<�U�B7�w-M.ĂA�i �ӂ�>�멲'狯�/�};�Y�H�h���ցR��N���G�ǙC���Q�\���,t:��Zx܌4Hݐ��P��l:3"��W�rMp{��u��eBI�%d��Ҟ�d��UBy�%�e2J��B�����)#���)�-�@��ɒ͊�d]MID$�dɄI��S�*)�W�V�p�5i�DE���!"�+S叜�I�"(D����T������c(�sC"[D��D;%F�5������ ��%@'��*�ICL�l�??	��ONz�.E+�{f��[ =�����t��LU��6[�%@��Q<��<"]0�}��r:�Uӿ����Ϩ<,:�����M�D�������՘6mZ[���0x�(<�v#��.��!hu(Ԥ��2�RG��lb����'Ű$�v:��&N�a�N���/gO�����E�����%�������~�BL���� �m�N.��))>��&��H�8�Q�+���D���8;�\�b!    IDAT��JI]-�6���������ASS���)���Ç����'?��#W=H��6�U�Va�̙|�/^����/��"����cs����o`�M�`ԙc��K��O��JeB��S�H��vACr�%*���p��(�NM:5J��oY_��2��3&��AKMM5���z#��^{��ۣؽ���!Vkya+����b��$�{��HT����դ(�������?�\�BJ�_ 1�js��q�`��iǀ�R<�d.I۶��}�{XwzB�	��� 'Ǌ`8��$�C:A�����A2Ǡ!#��2��Щ�����ꉂm�d��z��g1' �� B�8{���1���i�H� �Ϥ�m��v*�g&� ң,	�R@Q�*�����Ғ~xt�V���0J�d��A��P��ШHF�y�ذ�~L]LC(ĕB���t���Vp;�x���������Чo	�ۛ0f�(<�� {�3��.C��V��(��'���:�kp��+q͕8��ag=�-]��҄�67F�1�~ �|�s�,�2���F&@��� SE0$$a���mO<��m}9�UH�-p�b<JIKN;Mu����1r����/]��>e���P��,x�F��cZ���@�����
|�
caq�*9��"�)j�566C�"��$�dhI���Xj���0He�x���|���ƅ��x=���be�,	D����`��ⶉR�/J�!ݏ�ۧ:�eB�\N��t�H��K
�
y(		����*���>�Z��j����t,;C �Ѓ�OKd5�4J���Ͳ����������d�M�&��*w���"#��gÿ�d��g��dFܙ���z:��/��O	t��CF�M���J=_ Е��s)��*����h�fO%���*�S���'Y���i' t�zޜI)��j�ëx�z�$�rڨ1X�f=���rW��:�dZuP)L��R;�%���=)p @����_�u[�z����{��U�_�gz�����B5@@� �H��X����)!@��"6�"�H	)��ZBzv7ۧ�^>�{���Nv���y�<�ݝ�������[�{�a�g����C�����E�i��p��_�ld�~�mۆ��1gC�G���.s��:��xޛ>�,%w�|�����<��M1�(��ȃz���DA�0���rl��#�y�-8���E_��[n��׾q���3�jw�A!�b͚5�g����>�H&Β;���<�r�,X <��O<�)c=��#�<�(�(�I��&�D34wu�b����5w��,ݎ���uv���|��L��-#&K���B�v8�{�wq����G��1�R�����e�h�1���xM�9��xx�����H$&�i�|�bɂ�H6W�����KY�6�͍��p�3Y�FQ�ف��]���F�t�K����-�����+:ʘ?o�@�r;�$?��^�6w��M������=U01U��%*8W�~�=k�A� �o�7o�<�"L�D'�Jd�Ȍ��9$c#8�k_���(��o�2�ӣp7��AQ[�t�w8�$����Zm:�����7������k��
Dg=쏢g�z	��z�e������l��gx'�f�✟� �l�#{}�d�`� ��A�=��2j��At�Zq�/��^�7/�{������P�٤6C�|�p���P�6�m�q���d^y}^y�M<��*4�vK�X�7��d�|h��0i	�b�}�@o?��p9�e�I�C��X�u[Ŕe�h�l�n�f��� ª�ю��v�a��=ff�k�[+N�V����=��Q�v	+�:=�d�Âl.�\:�#��"��ɏdĮ�.��e����w�#�V</�t	�~n���J1�"oIo��B����̩���/Q�F=Ɉ�]��Ƃ���f�+�Ka����oqY/���l�ԜטZS�,��Y�59�HQ���ŎdLt��Ҏ�}{����Q�4f��R}��}袺S�x�����M!��?-�O��Yjz�S�ϧZ̻d�U���7j	��P+.�:eYR&H��.�K�����Rf�R��RX��?'��3tf���y���%��R���e��c�$�G��>����%�l��Htz)�Kt��H�k�0�9�sM�b"8sđ�a��.<��C��`�����6����	�I���ͽX��'(���-hl�/Ȟ�(��ۤ�˾�Zr'��F���X����n&�PØ$K��m�s���x]��G�u3"�!_���2�FH3��!m]-3Lzu+�^7��	�����%����ߧ3)��vJe�I-�qc��P���!G@�G^�ôysዄ���a6��XW'����ă�X�����}�g^��������������������hl��X,�����%g�\�⣏��m�a��{b����hl�#�ʉ�I�\����)'j�ظq�\�L��	洈�tشm;����;*�kٌ2i�v�?0
_  �s:������~D�
p#�E�̙�`������/3j�S䆀�ҥ�.NY���e����|��\Ѭ�-�O�R[�5>��'k���Y ��Yc{O�W�]��߼�z��'E_h�1�G1�R6m!���	fϚ�+/��d�b	z�[Dcl��C98�n����H��+g0Է�3���� ��L���Â>eJ�]��ւB�(�l�׆P< ������1�C�8���Z�+�0�`��PH&z<:��Ff���'���P2#�����
����ؿ�X�&J��,^�r	�tLuH���v``dN�G̗�����y�����wN>�;���Ӹ��eذq3۠�;E;�΃($𳳾��VF���&q�!A�/!`��@�$*�z��"�ɥaw�K�e�dP��ԎP(�M�{Q(R�GC+n��Wp�5 	a��i���_����կ�['�(�����W\u�ϱa� N=�t,�����qݍ󦺆v���P�F��P�=���Q;m)�"�d^�9]��G���-������?<t�bSSS�e�=k)8K�\J��k>�ؾ�w�}�>�H�)ꧥ��mu0����p{Q�a���Δ����P���E@�K��у����!�̌`�|g+e&���B��V�pwe����T��T����U��OV�S_�vA�F�j�a\w��� �D>U}����	���z�ʦ�8����
�������T�Y@����]}��HW_s-���W�h6b���b��7!��P��ds!�e牪s:-&8�6��1)[7y�t�l*�eRJOM��A���w_��^|{,��t��� \7RY ���h��d�δ�HT�6�[[�ibB@g况�A�K��z=\� ���Υ��$��$��t<��&�*$��e䅝��^���)���Fb0��2�Fu;�g	0�
�ډ���"����$���8jd�!�`5��H������у��?N4uv����n� �Ɋ֖z�)}}��C����k�~=;�q�_ĥ��t<��Q?~p��ڛP�<K>���t`��磭���ٺ�MM�w9e�?𣩱^z����OF���A�F_�v���tZtN�ｿsv_��7��[����hj�.��?��>�~�!�;�6�98�t&#<���8H#�h4.׌��̤��L��NEG{̱�6��Ы����*��`���}���a��K��W�j@Q�LT�?�P��=G=Sr��Ⳣ�� �b�L��l"�� �hmi��O�^{�}�
u͘�L�js@*���eB48
��}9C��b)�\1-��lt�.���ff��d���v��q��D�"c��P�+k$;-t�j���ڗB�i"��f@2V\K%X�&2R��5 ��~�\��T�H�&� ���bD�%���5O��R��|:%��y瞍���^/p�������hC0�R�=Q3>ܶ�Ry�<|�v=F���h�}!���!���(Pԡ�n�9 �M���d�JԪ_��bN��[�	[�q�W��w?ބ_=�G��u�x�w`����2	���;W����h�t���Z��:q���p�������N���Ơh���2�&�.�v��Cho���+��q�@"<��C^��?�^�1�b65�\.k�~au�ko|��֞ѯ���ôﴲ���%�5��f���54þ���_Gx;�� �K��#W{j4^Q���Xu�L�f���W��RG������.Hu�c�I6�����(U6��ҿʂ�� zu�]�}&�D5��TԀ����ڨ﫞��T4�Yr'+��[o��w�U���c�"X(����5�o�H�}5�Ij'�H�E*�FgW;� vkC��ѓ��F� z,�٢�@X��k�hnl�NwWּ��~�M!�x�[K�`�7�l���C8@ojk ����F�}J����&�%�,Eq#4��0��1�^[���C!�F"��2����0HV�d�[�Y]�
f1[��X/eK���Szo�{�:�^Wn>��v+±8�:��ؠ�ZD�-/r�6�L��dY��?� �ɂ��Na'ϙ;�7���T�}+���xm����04:�[oY��h�	'��hFs6m�E�W�+.=�������-Q�r"�����I0��g$
����R_�λظm����Sy�ݭ8��".���E�.[������~;��Z]��
�>��Ci)0��a��M�5�9`0F?�(�� �tF �s�ٳd{g��v}W�����5��5�׷�f'��&zmy^m�=��ڄ�v�7��M ���p��0$/�����X���fs�<�$.��B�g+Q����5ￏ"�x)�ɬ��l���m�ȥ��&9�@�.���T�bZ�/��6o2�Ln�TuJżI��s`�=�-�
4e���y��F)�M�d�B���E�B���e�#d�JKߺ�텗��dJ�'��	�Ztgd��8�u��҈~�4<��SX�n.��Rlظ	ϯz�hV*c���xHo:͸���Á{�M&�_x�M^�%	��;1�};��hj�.�AV��J�K��W^~U�����v��_<�h���W�@z�3)�u�m◰j�3��ފh`���.�2	�~����o�ˮ��]�_=�"���蚳�XR�-��D@kT�$�ԪG�*�Zd��@:���m�=��~�OK�;uJ���P��M�o|���������?xZ�`�[284ܛ�0�bu���=4��������M�R���:e_9�<���H ��)����W���L �O���^��`;�{V;��f�j�^��3���?Ɗ�T�^]�sȴd��9tt�������7��x�V1mپ�V��s<�.�\�l�d���yr�<��r)�9����_��^����ER���"_T�����$�[%�����\G%5�[�fdR1�_/>h��k!��9��f���嫹���n��瞃p<�w�}�5�6���z�V�G }xt��-c��jA��Q�����qC�@����DX0�|Ab���&	��,}��\��U�lMFO$8h�̀�Ş��)��c���:�gÙq:�^�2P�к2��"gJ�r�r��9d3E�;oꚉ�P�KZ��M�����݉@d �`?{�>���G���a�80���9���x�a�д:a�6�������_��M8t@*���􁡝���).x�����46�D��h�k��˯�wg|Ѩ�һ�8�ؓQ�܂�n�^X�>`k@(ĳ����´�2��F`����R����<�����;ޓs��x*�P8n�t���f��U`�jO�]o�V5W������������a{�`a���.�A�c�^�vt�y�,I��Y���{���6+he�nС�\F*6���/�!6lN`�5�b�=ȸ��ϼ �ۃl!!�ڒ.��^��U�f�((����C$J���v�,Hg�(4��R�u�d���1P+r\���L�X�JЛ��s`8���fC�U��B�t:M	V�y��	�V3�$:k�Bi�tˠ�j1��gPʡ���{�7��Ųn� ,�ǋB.O]=�9����A��p�%?Ü��uF����l.�h���Bl�'���"�I8E$E����~�g��ln�B ��W���mN��f._v�f�(��|��c<��ߠ������{�Gkk�?�|\q�5��y�����'�|�uh�n��v��ҷ�}*E��b"\�C[�CSHō��;�n��?<�w���1��s�O���y�������`����ӝ*�a�:�;�c@�����tM�(D�$�S�<)Wܔ�Y��Qq킛ꐪA�?�]6��l{L��
p��z�Z��U���"�JCS����D0��٣�?��C��I_���3JW���C�]�S�]�j.��S�W,�
Z���q� ��W^�����d�>���o��`�$C���%KA�c�8�YFK؃n��u��Y�o��,;��{�����8p���rY�@�8����c���Fl�ޏ}>46�Cg�!M�7�(�-<6t�C$l	�,�s^�׈s�̎�8�TS3
��Ib�n3�B4�C>��k�8��+^mO��J4
�A/o�f
�P�_W$����n�)��Ҋ�DQm�ى�h��b�q�tA)Μ={��3��ƭ���!WТ�{6�Z+,67�������(�������?�O>���_x���{��UO����~t%>\��/>&��l˯���m�����g8,�tN��O7P��n�YD���o��Yx�����������+�_�Y����8Ͽ�O<�:|�2L�6�(���1鴈��@6+<-/��q�W�ף��v�C��i+�^���Гi#���ger�.�W��ϳq����Q��U2g��E+D:������	)t�~{m�=~,
0O����~,P��?�b�Qi���tN1X�yg�j� b_,�S��3(!���k�����"l�1��i����!�����x�׿Fc�2��f��hVN��^�����&%�(Ǡ�6�3y8D̪�@4�l�|W�}�e�:lm�cQ���D4p���Kv44J�i2[dD[W�*-�RFĩ`4�`}	҉�%���E�yoE#!	��}�)زq#�y����p��<��6�v��H�Ël�~�:a}ۨL����A�S�3��UѨ���R�g���4��w����Z��0��ر��H�P���Sxm��hjj������Ï�S��v���w�y���x����/Q����b|��'�ܳ��?=��r��8�3�mn��oDA�����'�F}K��L\?�꟒��P.��'��rvs!���3�}����_��z_^�.|f�Ea�RNg�O�52%�{��/�����P��2g�,�2�vP�uT�**��}�:�Q�r1g3f�b$de��Z��醠���V �!5����#�M�}b�}�ܔ�[�^���a�d-Z$_�o%ZS�['���B�cVK�<ՠ�@��s�="Qz�-�3�ǹ?�9�q�&�B@Y��AX�l��R�"l.�Z�A���%�f��F�T�!9�`8���I��ދŋ�^{/Ċ����ւ��pځ܊m[w�#���-�wb�+�!�����#ėQ@�6n�W����eYO��'����b��x:Gc���G���|��Z�%S�}V�� ��1G+IeΓ�!3t*�1H�(���9 �K.�A<��bV/���Ns�;f�]�����N� x�q�W��ى<�
Ͻ�*Z:f#[��`s��mB]S������ނ���|�q<���8����c�%w��7_��k�b����	������y�:�i��F��؀��V����PP4�y�0P���|a�?���6}744�c��o�u�n�>o_�~���;`�#+��$d�2���3	�3�*^�֎v�%�(���&o��͖R"�|u:=���q��lYMFtˎ�Hk�f�G�J�Qq�R���ul�W?�f�[��5�i=h    IDAT���J#��{�����Ԏ�)��W]W9yE0D���eB��$�ʀyI��J�[Mv�M�\w�"�t�Ϳ����o��+W��Z[���҂��}�i3�8�EkaGo/:��*j[6*n�.> =��ȹ͜�!{Q_�(2�fN�R��Seq2�6�E���G�- @@��f�Y��Ҋp�/-�ǅ���cQ�A���Vc�=���KG{�\�����&����p�i�
/���������Ҏp<%�!ie�Y����ˌy_?�:�Ã�s�ԁxw��ٰǂ�D���0#�Ć�HU����p�LF��-M"K@��;�����Oz�gp�y�u�`�-w���"�ˣ���-�&y��5����O�KZ��<�8�}΅�"8������oO���t&y6��N�U���� �2�Ʋ/6��Ń����g���¾���g��=��K��n�D�lܧ���P�äI������á����n�h��gB�Q�Sa�@vv��>fʢ��A�Ʌ�Ay��[uOk����MO�~�*��(F	8V	Ϩ����@$m��ઁ���c�ߪ�>�LifMj�>vܕ]q�T3N�x�J���.փ�h�m�Ȥs�뎻D�ছoE*��E]��q��4����ދp���đ/�a�;Q���4���7��)34~nd�'	d��\n�a������3k6F���e�6��d	k��0��p8=��Л�rcBa�B��쎊V�c/�77
V2x�qN4���Y�z�M�0ط�X��wB��K��g* ��ףl���+��\���ßЙ�R��%�DT1�QI�"a�,�FfV�L��,G�6c%ys���Z�0�h���#�V-�ӑ. VO��v�����_=�(��v-��h�Sg��?�f��ݝ8�;��o��uk�E2���Λ��]�D&��鐙Ձ�;���n���lf���H'�$bI�(�b~��o��}:Z���ݍ??��&�t�o����:�w.d��Eǟ�Re���d:���&)�4e�� ������A���.؝�
�`0V�tT!hE:y*P��9qh��^�<�[�5k�Sk�ͫ�z��-��G-ɮ��j�]Ԗ���W�Ƙ7D�PE��\��L��a2ka��P*�
q�}�b�=��+/����q�|�]ۏk�Y�.� G��}w?9��Xr�8�Ѕ����K0�|��S12\�t��'_|M������[o����X�x��⡇�[n�����s��b�
t��X��L���K.]zfΜ�����Η\�-m͸�³�~�+�X*�Ng�}6�<&�y���������&N;�$��q�wbG�\�&d�E�r%���P�8���Pv��\m������C{�B|��GhpYP�&��Hۂ=样o��#.w=���A,fDR	��Z�f|��F�d0k��cy4u�į���\�/ԷuB�3 
c��y�sϽa���s�ѿ>���	�^{�M�]vz=�k�E���$��~�V�&�٦��J�KEB��p��ߝ��ɏ���G?�-��O���o�z��w.J�N���ʗ� }`p�H �k"������
VJ\�cr�im�k�#������`U�T�c��$�>ipQ�W��j�^��Y�|n&����ѢZr��R�Ϧ�r���
@Q!�QB�:C'谏y�-�I6D@�%�X�d)��җ���F1g�X��zt�?&+��(�P�d1�onl�,�=T��	���$�R�/gMʏ�
���L2�B�Vι�7oq���Q��"#]2nbs"�
8R�H���	)�3��y���Tx�I*<��*M1���=[7b��u�}�\C
[>	II)CKPeelM[�Ziu:����5�Ye�{2�v�$�2�,,6�R~��l�(�:f�f;�e��ds#������@gr��5�k���e|�i�lj�R����I�%�� ���=`S�B=���ۺc;�0����/8��p�.�pU �����}��T��vJ��b�4v�}��uK�����V��Ex�+�f���ȕLB��8�P���|B#;����2�H~�s����}���<I��^��BB�,��eO��J��˔I�[�^��H���Ts�*`��`�'(�NEt����}:��*�K)TY,+o��2Ţ$d���i�9�
qx�f��m�l������w��ÿ�=��쿯�7dq�����݁�38������n��u������p8�Œ��{�M �v��2���ģ�<��<r<N����ƛV�λo���ؼ9�s�9��U�~���ہ�����8㌯�lɒ��Ձ���ۢ���;Q(h�l�Oŉ�e³�>���n̟� �l?�"�WF�]rr�s�Ti}d)���p�9a5j�O�c7�G���n�K���w�����p O��tr)�&s�De� ������-���ς��F2���GX�} <�t���xJ,�WFFF��>Qf�[���M�nF:	�Ū���(J���.O�oZU+��|�8�`,�,�Ļ�^��k��c�{O�wOl�{襷��擾�����|�0���>�n3��zpt�/*�'d�J�������^��V:��ܚ9R���Y��؉Vz5P������{w�v��{���:��򅜰�.\(��1VYa�r�>&�[I�Q]��	P�[n�E�M7ߎH,�e�o����G<���،Ysq�M�"�@c0���P:�����vf����!;4Ǵ�]�1�/>�C��R�%���������� >�d�/�6m�9�LV�l�$`K�TVH8c ��5���߯(�Uj"xmXN�zWG3���8�;'a����^%D ��7,�q,��. ���C��[,*��"�(�#�S�Rr'����:\��4������wN�[����d�4���9磩�O=�
+n�-m��3;e���W}##hn��ͅ���&��>��R6&ɮ��M�x��w�Ea���-:�6��EA��Ԭ��-vH.��f������)A��xώ���lHg�(괰�dζgЏ`</�#��N2#q��1+/HٝLf�����-���GF�5�e��c���g{��,c�z�B�����V�ke��B��6��p�M�6�UB-�ͦ���X"�y-J�z��P�Om��$+U�<���1ѭQD(*��"�L����g�:\��E�Ll�����+F�C1�0���ւ������;wʄ�½���m=ؼu�ڛ0sv����{�E����?BOO���3��r�B�|�q�/��c�$�_z[�l��y3p�����AEj90���"����w�qb��OH ~�I'�=��Ǟ+ؓN���ܭZ�J�<�X�&f���pB�5�6�Ao���hTLo�ed1$#A9��F��0J�v�6sF��dto�����Fᴛ1<ԏ��F47y�O@�D��z�۾�G��c����:y�:�/��6��F1'�X&�S�\Q�)�`�����O�����]�ޥh�Քg�]�(J�c)�͇�?��=/}����7��T�f���WW~���6-Mk]{�#3Vr
�}>���`��п};|���R�����7c���To^-3Y��Z�Vs����ZRۮ���%]��W�V�F3��L�W}.���{����!c����P[�sx#TOH@P�(*��^k�y���c��(��n��7�_ ��W܌y�/��:�h]�f����/ jLz��Y��F�Չ�0]sy�4x=R¥n���EC���͞����z�m�,��4�bڴ���{�ц�x�w��K@�&�(kl��:/B���`��z��Y�%��cFN�&0���ݝ��نt2�l2
�͈z��|F��h,,@L�;�gf�ʜ���m����{�V���d�����_�/G�� &≘����荍M��a��Lv̜�F�1@k@�����QV;:��K�adp�$�]8n�B[g2�"���,	��l���)׫��l�s$��.l4�I%��L&�����&�[v��dA�<&�'r��,ۺ�~�kl�i�m���F�ǕX��	�Vf�#� ����Q��d6#��\� ����8���F/=	d�}�,w��]u@+��/����-�Okە��DW%a�Ț���+S?c�,c,� W�\�j�ܳ���efM��wA$g����Lы0����wRTC�B������2���y[�JT�8l&dY�����oVT�e�b��0�E�Ĺ���:�?A:�J�M?(ZI���r�"�/�>ϑ =HXc��l��u/�sH��k�9M#�X���
��L*	j�7����f����|6�H�-*+�!�XPO�M:���I�l.��7�2y8�MH��`k�4�l��쮇�B�L���$0%�OX��&Q��5�|����Ud�ſ��jW����u�1�b>��)g?��N�r���Gcj��8�~ѓ/�j�e����t�8�>�H�7:�9�[ }`G/F��QGh1��@T#��z������f۵�. W�"k_m_�'[��njRꯔ�k���d꟥]YE�S�8)��G�a���C��ƴڹ�V��m�n�tr��"3&�F� �=�7ڍ+n�|���Fp�h��F]C����Ԇ'��O�!�S��Eb���5��X� �`�I�����B%1t�hl���b�1��� ��d���Lz�[����a?F�a���C$3YxZ��i$��(�Q��=k�D&��$�\�Ã�?y}=h=K2[[K#�� �6}�N��8.��Ee���#i�O׸<�ו���S�c@�k�kG�^oE��(�
��1
E467#��f���SI���!�H�h�cӖ^��N�BXr��"�V�G� z���D�nr��Q�yy���.����T�K���Zс�X��Dю,"ѐ�֨@+�`�/s��G~��X�s�.A�,�j2Y�7X�3��'�5مG�mj���A�X�?�k���R{.OY]�>cP(k�N{&�H�Gr&:�) ^��,3�	���R:�j?�d�g�2�������]ZxU8�f�Q;�cr@W���*�J�=�`��+��\��tZ����{��o�fhijF`tD�7>��$s~~�.� ��D����Ћ\G7Y���أ�ϫH�2�ł�����SM�RmaՇ�?~mljW"e�HWs�q}q20Q��ȹ�UG�)���Z� !���Tc�Za�3�e�*��"�ʽȤ2B0g`K�&9�,���ݾ	3:[0�s;�]Hƃ"�L`�q��aDS	)�;]n�,V��N�eD��k&�u-�k�HX�2H�K��\:'��l�L����+�<f�f�5d�"�@�I�xDo@�+�q�@>	�EΧ}O��g-���Ń�����|������FR��S�~W!��|#�ё�,t=z�]��+�#*۽r'OU"�>�I�S�J��M�
���'��K  ��]��Tp�<��Yz�@p �����U�]���J�����k���3��sa��0W ����Y��W�$��K/_"fm]]�A]}�Y�bфd�
�hi;X�V�Qe.���E���2��r��� �z�Q�O�э��v|�������n!�����z�O~�P4�WV��C�8
Ͻ���-��H�|Q�[��1g�N�e�������F�u�XW��)S��?>�����eW	��󰡰�k���Jɝ�0�Q��F�������\Y^gY���%2� 9�sf�����8�e��d�'�6�P�l6;�_q�]��/���^X�z��xf�K�/IDDh��S��0�a��ǖ�ۑE �^��	�L�N2����a�ٲ?0"nKV�Q,n9��Q6��==��J��Ή9�kh����x��px����a�?��Q�����5.�'�����F�8I��_[���%�i�[�B�TM��P���*=C��S=d�����tt����w�T������iR�{���i+�d��(�s�$+�H/��!�Yr�(�:: �Y��V
�8�Ť����=4[x�N;�e��/�y��� �uu��@�A�n�}F��Z�:�i����uf	ny1��|�Z,��T?�o8��H5�׊Yz!O�e�d�±`i@6����g�)js�i��ב^G����yڹ�e|�{h,UH��<L��9h�Yh�i4���;��O���k�$�I	�#����X
�x
nO�(i��4u@g����L�BYڔ,�3  ���,?sf�hO�FG�BI-�Q�B�o`�Yz�fť�A)�۪��S����g߹�S��:?����עg��h�h�rT���E	stt862<�=}���>���q�e��,�q�����8�?`����DV�x�{j���w��k2�Z%��M�������_�SmNc���������
�qK�"�ʅ�z���e(,}�(T�rt�=�+�w�{;v�b�u7�v�9瞏�7mD{g7�}~tM��m���2�A�g��9ʫ*�.�4�	�TBX�SbF���~�b̗w���9D��-���މ=}�Lظy���b֜�����q,�݆XL�R��*��SJ�J�j����A@�qjj�Ⓩ?�������Ö���L>�3���Ҋ�Ug<�M(Kֶ� ���IO�I0g���=ߟ �Ϊ3�	�9�ì�$cX�9g/��kcS;6lځRق=.¶�Q�G��-v�tt`$s���!sY1��3q��Qf=P���z1i�0�5��N�L���m����W.�I+՞z��X\f�l�̧�(�!�+Y��BVJ��`Z�M��;=��#U�\�$�,��}.Y��haV�]]c�h�s4)�N���p�og�"~����VFˤ^mN1q���SքE��O����{5���R��5� i|o����~ٓ��d-�.�5-w޷��0n�)����#��0��z$ SD���I��{��#`n�Z�CCH�Zet,�ʎ�c����Лh*�EY���┈�h@2NA'�L�eD1��fwK��6�l ���+�_��CY�
O�砂�v³�
�9�'�Y�rߥ2���f%:��X����B6�1V��1��{�p�$�'�E>�{��Gm�b�����LqI{�w�%x�}j�;0g�<tL��<�,�]�u����mBh���Y�p�7z3��,��8�0p/�G�-(=uUP����l�	�3���lf�E�0
by\�'H�哣����o]r����/oj�ܯxr�������`�yx�l�đ$_���hdtd�%�8��۶#8:���zrY�l��R3K�Zc��!�F���ˉՌ��}J�_�;���	߫6(�C���A������ZZ�����^�s�=���eᩜU�s����J0����x���ח����>w�y7�}���ۤ��d�2���:�\���ՀX")d�S5��2T��(����w�m���ʕE�rv27�ʢ$�P����(e>�����V8���VdI�ZQ�j�'D�}~f��|�fs�����C	�|o�))�<\0�Pd�	x(q�� �����\�� �����0��(Y�hhS�Z/�G�޶m���̟甌H���|D�A��ܘMl��l|�(�ju�q�#I�hi��B�@Wf�x�ZE�'/��%��gF˲(O��"���&Z̼(�S�ge�W��Y�3��3jE~5�����?�L")
�@m�-R����0C�Q�%i�z��b�Z��a��0P��n5.�.���r�v
!����g�pY�"������?W'Q&��t��F%'�55R���Ɗ���E�}dVp�zmO@O�A��%Q)LU9T�ޓ�&�|'�(�c��WS�]��一���O^Q���5��tsIHYJB�4?% �(I��S��GU���9~ɓ(�S������]�-ǖ�QѧU��0�x?��r�R�5r�����f�E���T����V	R�(�HR�P�i�>F� i!Ѓ�Q��mfttu
��u2��v���O8�Lo�C{�sg�c���������]��I�����p��/��7��<�T�()�����47���E+.e�MT    IDAT��Az��+�M(Q)��ެ�왳W^�o ���"Iq� ���\6�� �6�-g�o�E�����/��69^~{�_�xǕ��e������h����B#C���A�m �ˮ6í� �/�����R�U��)����k}��':8�
��X�������)�{�����آ� s!�����U�4������1��.ǵx���bd�'Lv��\v�Ux��50�]"�h0Z��N0��D-���Bf�2���Xj��l�,k�Y�c����(e?F�����4Hfs�1�*k������L��pC `F��>�<���V�`pB %83���`��=�w*���܆�owܺ�p����U� 3�mc�NV+?f��J@%X1���PH�p�L#G���v�R֔�ہ�=;D�u��y�����ǻk�㪫W�s�<�5������"�L!�ʹ4����>	*tZʶza1Y�q�@j���GD7Zg�(�q���eػ,"En_�ؾm�����r̭��a@J�v�CX��P�;��$osK'��0:ź�>�;k?��U���ftL�s�a���!�L��\�:�*�ʶ&�(�'`.xEϡ�cU�
�Kս"̤��	�,�������:�2�%���T �U�#�B3�r���cF�$9/z�y�'���*��B6�'�L�mP�U�`>gˠ�����(���2'�S|⪺oTWA��$�r���BS��?>�T
�{��,�T`�\�1�0�ʘ`�p��|����q�J,4hA�+��8�&^|M!��2b���X��;���~ه�w�"�D�R�s���"O������m^�s̙ք�o��G�����1� ���]�܋��i���_��s�p|��x;����}��� ����>���}�)I�T���MS�i���*I���K�*�X�K0&נT@����D�x~Mlm�o�p���_�o__������'��aL��(��R��P!���F���T@���J���fP�_eUAH2�J4:U\��n-���Q��*���Ы�����߮�?u�[]2��P"J���0���ﯰC�LW�~��h� ]=>5Q�ߒFqYS�S�c���{��v��h�����&�u�H��ЛlrC��B&5}�Y�c��J���Vtʧ2�d�˹d����,*�9�2��L����8͍MBh�짍�q�I��اb��
��H�����b{�,���!�2�`�gE��y�]KqZ���|̗C!�Ć��btx N�M6��]!cѸ����:[�pG혩3���0��C!�"�H%�4,z�����js�[�*���}><��Ӱ:�Ηel��؂�`z���։8�/��0������?�g�܁ �,ND�XMV�מ��َ��!|�/�['}]�F�����N����S9�[d2AW{�䰥�ܬ({m��'�g�͉��Q4����oHX�w��[���1�TR�8�Iy�d�=��Ȧ�`9u,�U�s%�-)Sc��E�ͺJ:ը�&@-Q��t]%���JzE�o�/d���eϑ�a������YrQ6�	��ϛմ�W}}u�=t����M�u��c)[�����(��r����v��󭀶$V�ҕ��X����+R�H�Ch%`�B[f儿!�P.)J��eO|5�'jV ��9yME�N>S-����Ub��TYC(+�GʽB#f���))*�<9*�)�V�ق�ϯ������-�>&�TF�\3����ҡ��Ⅾ��YmH����� �Ϡ���`w��+!��|q5|ᔈA=��%,>�|���P��x�M�� ���S�]^�2υ�q;.���L�׽�W*�g�h�TT*1٣aN&!-������G߼��ӏ������k���\�,�a��I�EE�����5��N��N����Q������(�;̤�P�:?ρ�E95Y2�d�Pg��f���%���m��w��
iG]d*��{��A'�t�Ac=t�"-Z�y���A���׶�j����i��W��X��h���Exi�"�K��#��s�l�۶�2���8��	�̾v�d|$��7Gw3a6EC����\e�S)�8�6���1�Nا�Vau:������tc2���ˤ���C���t̞9�.�[�F�h>H�����+0Կ�B��u�<��v*�u1q�e��a"����3[^�ȡrc�<�����.	#��"�S$/��������@�ބbQ)�m��Ö7S&�6G�(���yQ���{ԋ틫��#�Qa�66�c�3V\�gɠ��7���� f�	_:�h���'��k�B__��#n��|Ի��� �N��`1����o��m�&�cdI���p{��|�m�BQ�^|�#��������������p��y<M�z�	q�br��O���J{�*9�*SS,@Ռ��e^��Q�L�*����U����W�����+hu?�LE��\T���\_�ngiv��rTJj����*)���N]BW^;��-���Gy�j0(��*��-���j��z��-:��f��5�����=�	V%�B��=�l�U�
��5p�i��,g���|����=V��˺b�NR��҂���%8r+��J�F���اf�^���AP�6���	���Ȧs���DX�g��ͯ���ߊE{�ö-c[�z�T ��fw��c���r��-j�7Fs�h�.��I5�sv���z����I���(6��B�K��K Ȍ�Z
��z��PV4�sI8-�|)�hެ�+�����;�R&���|?�ݫw���������,�3t�vћ��>����P��
����:�_E�X�Z�1Y��EVn8��4V��a�O�c�_��0���,pg�W}T�d�;�k�z9O�ѫ�Ku��:˹��Yr'��d,��N�^�U�
�Oþe�5<01�K�N��e׮P ��K������؂x:�ь��f�w���11��@
3s��9�>���@4�9t��%wi$�R>&x�������TN�W:�E��~qU�x�?��ᖹS�:�74��}���HVLF.�����F����s9l�sjm�G�6\u�������F*�����j@W�O�;�A"7�6ϟm�T0��gB@�9��N����::��*{ǥ�0���(Z;:q��~�կ�����лsNO3�f;�9F�zq�:���q����3NC!�ApdW,]�SN�.��r,]��Y��y�>z3�x�=�u�]p{�h�hǒ�/@[�0<8 ��m˨�C6G��s�w���v��MH�3�֍O6m����Co�b����q�1�a�ǽ�y�^� G{�^�>��?����׾���~�ۿ�7��?��9JqJY�b�+ ]��g@U�n��!kAJ���P��Nؚ�(�">S1Y��^'t%�P Nf~+���jB�Osk$pM�=�jm������U&1�����
F5oNI�����`bc���Oʈ��h�WT�,Ou@ѓ�p'��P������ă���+�W��Ӈ��l0TsIX^�Ck0��7�af�PTF+*j�J�p1$V(HK�ewf�ՀN�	q�b��G@�j��|F4:�(���߆&�	u.#�8��x��08�Uȁ�+)����=��?����@�`G&��
���Ī���a���}�~��?�e�q��� _E/���,Ĺ1�i�_q�3hU��b6	�I�r1p�5+�{��?���͟�'���޿�|������9�>���nI�,�P�PM����#�s+Vxcc�@'�(��)zk5}�Zz-�r���՛�d�����V��N��6��9��J�j)\�7���Y�%@�9rQ�</�:Ʀ�guϭ$���S��/+?n�$>�u�=2+L@�d�W^��_{S���P�Z����ɦ��k.V~�\��;$�z�X%��\��U�V�x	��DZ��S� �&�#A��`�ob��}ݑ����|�h$.�Z�,X��Vz�jB@�\@&�R|�\x�8S=�����w�6�Xɝ��%B����T6%�3G{�@AƳ�z��!<?�o��.�'�ل|�V��)��/k��֎#��*�|w^z�-�R%��Ze4����6��t�.��,\���2;n�w�n��W���ׯ@S}~r�YزqZ�[qѥ��[� ׉�_^|6l@*�V��<��oQH�+,q���׋�ӻ��b$�9��x�z����(����ⰣšG������?c4�C��=���up68p�ݗ�� �W<����GWA�� GZ��V��H�
Lq�S ^Y�ՀΟ)�;�3V?_}!Y�U��S�U& &����]�~��L"7������T�`��Ӵ҆���T���s���+O���g[SAP3av����6��
)Nm�HnI�/��!�(d���f��G2vu"�+dH�o���<�n���V��\��\�Wl�YZ�NYq5d�+�e�V��צ�N'�M�	�����نlZ��'ᕤ.��X)����D8m>������1�����6��sf����}oO?�M�����U������{��$r�6wb{�(�e#��X+cv$�)ddV2y�l�1�`U�D;�IH__�\{RJ�I��g�Yrʠ�]�r.�R.]9�E[N�=zm��3�<���<��*��ܰ���+k�}"Y�RZ��d�"����-�8�w�P �mh`pƌi�0�),�}^�SJ�*ީ�Ê��E僭&yN��O���HU�^���k��v�=��\����x5ȏe��Q~'��*��8��D R�?�̬O����V��&�xXA�x�:>�ƅF@/���1�ՀN7�믻ED�^�����d�k�dJB��A��N�f���	�Y&��-�1w�n]�Ļ��Gz�d�+7�2�%S�g�R7N���p��Pz�[߄����LgDv��Q�#>�I�`��5�FzckQG��(�1������}(���mF�ɸ#�w4E`�z5���&r�ҥgo0����
r��;�{f�>����U�^�\��^	����űyS���P�����lκFtϜ-��T"�;o]
��F��� )�O�O?�$R�.�t	�:jo\|��2^H�<�� ���yL�.��a�X�r���G��-H��7{���i�%W�#d�3~�u��K��fn@�sȚN��wH���G�Ǫ�7a�����ۡ�hp��a���(�U/|����*�yF}!a�r�U
���(��$ʃ%V��v����U�I��\�:PM��z�.+{���|������L��ޥ"'�Ԡ�KQ�2�TUN�eW�������$����2��S�Wվ5���+��JC���3�C�H��
�K�U~?v�&^t��Kis	Ϥ����� :8�.�ʊ�� a��'��%�g�.��:��� g5�s��,��]��U��F��L.��xg��;�3�.��о��i�77����㾎�O:�_�\t��5w.����m��N_���!�͘�p�~��E���"Σ>9l��9�8����+*���3�a�%�P���QםĿR&VaiŜVz�R&c��w؍�}��C���3��1�U�V�~e��֭?7�(-����	�����x�Á������t��8����@&����yL�d,�a9�6��l1O�aWK9�ѩ����Yү��Q4%���H�X���}`َ��r<2��h-Ww��F=�U�Z5˝s�
�]}��d�%��WS{�z#E*)%b��w�nA����n��7�B*WQ���V��"���;u�3)��ϒB,�CJ�}�[2c�m�V<��S�g���+��_������c��k��G�x$�X"�����x��g�sy��A���f��+X6'lr-��d���:�����G��H�<�\(�������7W��^[Wf�d�sV���{ls��B�,U�����������%������̞=[�Nc�\.�"����C>?\nl./:�fBo�ch8���yvW#`���m����{�fv�����
���z����C��g����N�6k6n��fL�v��'���W]��i�1���ߺ�w�fYYe�s�=��T�+t�t��D0���qfF�t���Qqt TtPg@E�b@Ā�M�&u����+�[us>������:U4�}����<��<<EUߺ����{���Z���'�(N�oT��[����)���8�d$$��LVx.�<y��c�{�Htcպ��O��S�<�N9��Kxn�֝t�''1>;��%\x�ؽ�E�s6fg<8zx�M`Gl�O�`̄R��J�PչK*Yb]9�g���i�;Q��TS���]e/�G^�HX�|7�us۳���B�t�� �+�}S-G}`S���`��j�r�����PzZ��#�]�k�)�l3AP_��vv/���8��~��&�T��g}���9	�b8#j$�{���:&���řR�QF�^����+H���T��=�L|N�r5��?M�Q-�15>rv��_���B~w�:��_(g�7��Z�s2V/_����.~�ۇ�o���s�|�|���#m���x�"848�_>�8���#S��j���$e�T�p���L`���2q��r�C��#�HA�Q���ȿcqGr"ż�D� <�������}����-�t�X���9'������u��K�zE��ǎw�:�����9�?�W��ڙU_4����	���PoTaLyZ;Za�N��^���-r�G�c&5)$$�I��y85���3�(�Cq*,�T"un�:�r�����o����j���I@wZͰ�I=Z�2�$�8��s����H&�@�1�+`��Y�FV�d63H4!��^�O�m8��Pb2W5�FR\&[��}�F��I|��6!_���B�\��=ΒKa�3�*qS�ҧ����9�b'�[���V\q�eػw76=�$6l<Q�m۶�v��fUͅ��x�%��\#�᰷��U������GGG�r؟��lz�lTd*%kw`��LW�rd�Vay)cZĝw|�1��կ`�� bш�L����W�/G��I���M���I��) >/|��.Z�3�)����c6�����U.��'��w��o��փ�7?����D�]�&�-����ǰ����/|�\�D�\�Wo�駟�w��=������m�}��������?�	b�Z�:����-�X4�+�e'Š"�����5�$���*� ���#�x��O"������b��T��/�A��%V�"J����f �i�8[�?�����5�@;�;� �h������e7)L�_���X�Y�n���Z]m�k&�ΞC=����5�@*	�|輌}.{_��E?�F�;]Ū9w]�	v�PE��X���iJP3�W<��¡�*ET����Ss{����}�z�CH�ck�hQkKޫIr�ʵa�X��lʳE�a�T���	Eɑ�D!3���et�K&[�!N��,���^I��qRk�[���ύ��I�\:'����G�Qr��f��NZ��\x&�`dp?^}�Y�-X0A���]��6�z^��/m���i4���0r�zQ�R����@�]��X�QM����	���"�Lbxl\y�@G!��LS{=���Rl��O�
�E? Z)�ШQ�р]/����p����g�\�v�#'��q�sQ{��sQ%��r��ı��ã��Tn����KR��E���j�
�O��@��r�� �v�@����]cc�z�{���?���	�wd@�v/���<�=�hg���7� /Y��\?�MX�����Ap��f��缛h��vu��5�ݟ�JP^S0�똬8
p��q1�����LG)�������FƇ�Ixs0_�ϙǕ�V�*�A��>��/�n��7�����/~��x���B�&D52�	�����V�^��E�IG���F63�5���|Y��ʷ����DjF�</V�v�~��W���9�\��fvJ�ʕ�'x��G��ϡ�g5�~f�Rh��qt:R��e4��W7$�SO�â���e��A<B�`:Z��������&�D�,�4����f    IDAT%��(�y�� �ߗ���O�V�w��L����r��{���j�r�c�c2�D0<:�cC�H�-�!��^�_�͗Iv�X�c���ǭſ�Y�df�O܌'�<�m۷����7}?�����������0>9�������X�z	�'��:�&#����n�� �I���M�i�ʌ����݊`���N��5��� )@ֿb۞~8<��;c����E��aڰ�Щ
ÿf�1���.�
'"�0պQ�4�ѹyf	(� ��0d3?�㼄�	��]�	b��* ^w��]X��"��'�J=pn���ne�R�e�,��N���1��y��&�N|�]PS�E��5U�oos_����޻dnZ��.�/�;��]Z���{�AM�lL�E����# ���g�$�IzkP�%,�\�T�dq�����0�epD�gE���C�	W�^'#_:��ĠH�F�o 33�F9���(���eq������||�_>(I�?��}��7�B�T�s�oG8Ԃt�F �_�鲁�?���
٭:�]�DØ�P钒�-�҂��rrN>��*oR%��{�J���e&]�׈~�a�U��X̓�����#��1O�Ƽ^;����``��1"�R%Q���*uO�ϊtW��
,��GMP�j>!�z�a(T ��Tf��ȱ��zz�é�a�����̈́OK���d����>f�����z��U�k3p/�f`f��<�dɲ¨R�W9��E!�_"4�ꥸf��=4���cq��I����/��ŭ�����s�V���
�4I6tDf�8uCR��_��]B������S�|O?�Ŋ�L���?�j6
f�*�s����p0(l��Q���N,/�|뛥_�k�	��?�0����-��T���v����A���g���~��^���=!�-��/�Gd%�"�d�;��l\��:�>�[���02<�+.�;�����>��5!�A�T��F��̟�o����e�fB�nH�����$���(d�ր��4��*�5^_P\�hMhXT� ��e�Z;�����lVZo�x���FjzJ��/}�%8�ܳ�^�-��o~[��}����_%�ԇ��ʜs"�a�Q��`��8��S��L�3OC�� ==��}="�ID�HE�\^�{jr��c���8p�(�P1�O���GZq�脨c�AQ�c�EϷJ9�`X�H0"�6׷ �7�V�
2��|�
��ri����2[���׷F2��)�ywBp��Z����O�Z��G��5j�R��D�9�B}��~������+r�NAsg��0ؙ09Sb?�B�?�����L8HJt�#��\IG�w~g;-�y��J�J�]�
U�L�"=�u�v��+R�u��uCa�'a�Yt��uZ��9�4�5�+[�S�7�)&<rq�JT.�=���G���+����.��)k��D�=�$.��bA$���������q�_>�0E�}1F3%TH��?�k�G��#CB�?`IR��8A*(� ���vC�w1ġu��j\���?#	�H�^^+&CD��w21a�_�QE�*�E��.B�R���z�Z+�m�Z��̺߲��c�0�,�l�P|Ax|4ݲ���Â�����SS3[��FN]�Ӌ�ߋ##55.�;U�H`hfNΌ��E�W7Q�L�i�N���H�\�[��ݽA�!ֽgw5��_ۍ��ۜ��<�MLс�3�38�4�����,���'�߀�����EL�J�Fɭ����t����9j�_ӑ�y-�v�]:6��>�)$���[nœ[�G^��!���@��]S1N��%�RU[".��5+%���s����
�}��?��d�<^9W�W-�<�p�=�\,^����'qɫ_����k�~��-I�T��|H�wI�:G�%����L	U�hkMȘd,����j�,��뫤�DaB��r�����j`���c��c�ug�� �9tBg�d82�k��ρ���� 	h4q�}�184$��sλW��,Y��<�����$a��B�!lW())����+�l;��PP6���I���틥d�(Z�tlZ�z-<,�� 了]��a��Aî�Z.  7��d�s�JCZ�C��y�t;���8Nɶ�j&*싚idO#��*U����I�XC�g�҃��5
�p��e�r��Ri�U�8*7�>�U�`��Sg?9^�K+������z�h�ߙ0�2U����ݽ�&z�{�J�F���isV{a�}.�3�/�,n"	�ޜ�qs�3yMj�ñ��Yԏ��;U,D4�i�E���ȕ@�>K��5	�9��'�2�t��|^YwԹ` g��k,�:��*)��+jt��)�OJ$|�H�r��x�)*�6���4��⵸�O߀��Fa��5~p��d�����߇+��3���pR�~��&ء��V��i�6��G�<��mAN+�p��7K5�[[n�N�U���:G��,3��e��dI\�Dפ�l�ay��[d���|)#�B2�}^g\�Vʢ���3����=�N�^�)<Z���=M*�������S��-��~��A�&�d\�S.)�$38~�>�{a/�m��rl�?ֱ>�3Oda��y���ޝ�7����B�c�V���8?7�&��������&��T�n&��OL�c��U2��YJ¡��y�I�`��0s�Z�|����Av�)�n��DL|�k_��c���'nA��7|�l~f�0�Y����Q1n��*cI��Uf$&%��M�)<��S�l�R�^��^z)~�����			q<>��Z�?�8�}�e�I���g>#�6�6=�r�F����	4�5�ʹȱ�%�����3\B�bC���q��g��%��y�B�������7/�YQA.��.���y�Z��0���g�=�'^w&a�'�V���I���i��M�z��y�.^�c�3�?6��̘T�0C�B1AA�tLL��&G�IN0a�g˔@U��Pj�J|�U�)ژzn"�i]&0D1���������Wme�Z̫d���j�d|�0F'��%�����M�QG��!^/=�=�&�s��:�|�^�$�Z*�x�� �{d)�,�^%��|�K�DK�`�95ܪ*L���km��*���ua w�̀������u@?^`}Q�>�MNo���4���P�j�STd�o/�&�id�aQ�pa�S'��MT�΂�Y�5��~��Dp�Oן��Y����s�c�+~���<�8�L�վ�
1"LԹϰ�#��bQV�
n�וֹ��k%4@[�:�q��@�����߇Rf
��yx��'aUO"�:~��O�z	=��E�r���x��G��_�CC����c���ر�_Hq���c-ȑgT�E�.B��-�L�s�(�J���'"RY�!�7�*y���2ҚC��2؎t�F^;��B�V����^i�z2	C-�� ���((�a�l��6��8
��&5d�Xl�'Ǧ��=}ْ%|8�� &�G���MyP�Ǣ��4�������Y�;xK tsP�~4f��,ua5�!)�y��=<�[W@�=1EBqf�>	�N��>g�n�?����as��W�΀����o�%���8 U��U�!� �P���p�P�����٥���A�i�|>���|�8|�(>~�'�w���	����b��ƥze F�n<ph�*c_����хh8�p0"0���*�ǃY'���D�Mu7N*����q�B,�l��'�-²��(V<�D��Rl[���<r�����8���dzj0h���4�F��LZ!>MJ�)���-S<��`���+&<&"*	P��{�{�5��vfY��&�v�g������ �3Y���X�j=JuSY[����+b<�Z^�#�ID���2���`���3���@6���n7�H�(�K�w�dj(���>L���P��k�P'��4�2�{x}��V�6U�*��tH�� kX�^U��\�I[�~�NM{eS͗��D$��(U*"��/^ך�L;d-kҩCs��f��ҡ��]�ׅ���糰v����ɂ�����YQ.H�_�=�v��T`lSS����L��������cq*uUo�H�j�ս7���"�}=s}�DZ�>�U����{0�3E���{;��jU?��:�8ɭ�w�jMqbjJ�I��{"��<86�����&R8d�9&=NW3>��b�Q�9��Gw2���)�W ���Gb�d��atr���wallO<�,�'Ӱ=a���w�`S��0�j���d�mI�;*�#'����h���d*�H�EFT��K��~2�I�@S*�A��2�"g͖��'�*��Y�p���r\��=�(��D�_���g���=-]i�dx�h��7��	�I� ~K
�f�>99�ild��eK��ᐅ��1:ra�1cS���Ct��]S�qZ��Y�;�k�p��ug��ݝ<��D�&�͵J{����@4l���Z�}�@��d�J��"ň�sp�xu �������6d��������_�/|�H��J�`��K�,]�QdbKMZR*U�8����>ě���ǆFqÍ�F0��?|#|���x��٠})����,4���(�E�r�,��F�H�5���G�b%ȬQ�a�U�:υ��5�!6��f||�d��30j!΢�em6���`8$ɉ�S�L�G��&
�4b� 6�_�5+��7����iT���!��7l��d�.�x!��PU����7�2P�H=���y~�>pJ!�'B4���z}�X7�|�u�{m����(���=��h�Y�`�l>_�F�xX���5,�u���N�P���kί�e"=>I�,?Y��ٗ�|HHc�ń�p���[;d3�m��`��![1���ho_��)��w!����TeF���q��̠�y��D�]�,��ׇ��:_��Bs��6M&�y����kR{�+tknbF�1V}�ٺ���~�	�{OY��������:�L�x��E�R����o	t$��u!*�?��w@_��������z��dD}�f߫��ڐuR�*s�|Q�'B�T�^�$�{�jٴ��-7�l��d�P�����Q�M`f'�����c {���$宩x�����y�G3��DHx_[��#��r��?��=���
�
z��^і�۰�s)re+�*�.Zڐ.�Pk��A9_BO{+�:�(fӸ��q�~�������v&�t��~Ë`4&k��U*�Ē6A�|N�h;�ϧE,��9��#�[>_T:ф\�5n�/�!r��P�����6�a�����6��HA:�r�}�s�pf�Ч�R�>���K�Z�� �<$��ה�k�Lȝ�O��HPs��	=�w���������#���2e`V����#���RAde�d��朹�]t���p���h��*P�T�
�P��i���
x�7�݄�	W�EA*&��G����!���1鉰�*{U�K�5K���"	�,6�T�"_ �!����h4�w�!�T7��)��6>𡏋B���r]$)O�/�Йa3�v�J/�Ѓ�6ꬳ����a�q�V�'��$�0A3�w�� �10����[�dƜi�����+��� �53X�t�L~��r�9W>�>�MbgG�{��X�r	n��11:��e
d�^2�b� �g�y�X����A��Dhj�KPr�.�?���Ǯ��X>���7�t���1 ��	�^��֬�}<�g������&���
'��ɥIěIE6����-�ka ��y���.	�]G��㴭�W��{.-�x����t���Vw� Y�>�l>_�A7`{9�@T���� ��r�d�Eq :��I*�dӒ�0��5b��/n����&��FLA�f����[hzIB� �Y���d
vV[�3���-�Y���߻�N���,n?v}�$�M���A����VYR�)�*_/�qsU�*\�	���4�x�S��k���x��o��F�u�����Q����q#�^�D��6��*�
�>�ƽC�υ�OYV�`�M8*A5�=95�a2.��Ӕ�G�	;���x�+TSR�����H�h�8�FM���BG��ߋbf
� ��℥]�J�q���w|��)���l�Xo~˟���6cf���b]H����F�/(Ē�pɢN��Et�%����$P��o�6�FƱw���.#j�J��Z��`z�LL�&yX��\E,_ڃ���:��Ʊu�3���#x��(�?����ʄM�R���1���D�7K������#��D�a�� :�����C��B���蓓��x�����u�W��ۇ����v�7�b:!�G��/6Q��Ke�kJҏ�+%9=&���(��ʡF B�=%�72G��R*	�Ǉ�K	AV[�0D�T�,�o B)��g�����){L�;͞(�"������&4̙qV|�xc���᜞�� ѳ�v�"i{[��Z�:^l.�H�Z�r%��J����NA2т���j���������*e2e5h˃/U�,I���<r�~����ʁ0��_����o�S���ྟ�=�	�|	� ZA�*
�IggEx����]��gO��`OO�����2Յ�f��t,�`�"�u�q3�p��U� e�*�&&`D.�z���Osi9X���]MI�����l���Y��^���c����$;ڌ��ԕ�;7�Zdl31��
Up�:��\�3���q0;�Lx>+$��ΦP�d�H��0����c|j�E���
�a�1x�qT�m�e�$�U��kMW*�q�>�H �ɨ����1OWU�ʉ�?1>*P;�?�bN�ΰ��l=�_��y��
�9%Y_�DW�#N�\�#�ˣ���R��#��D��@0���d��v����Ų>�.(���n�Ꙣƽ6�Ȁ!���X	�$�r�W���	:	t��嬯��Wς*|~%�Ti��mI:�Nf�AĀ�?�Ȝ4y9�TGc^۵�֛T��82�j��(K��L�ز�y�P�MP\�yV麷�����ɏ��_H��܂&��sR.um]| y�T@BH��r=H8�]�V����(r���i2����#�C�<��U�Ұ�e��N��#��hdnF�k���1��1ؓl�x/�R��$�����G!ˇcG�����k/8�q�q���=��_B,D����X7|��{?B0��>�i$[���3�pt,���N�L�,����j�*�Q�%�������w��3��C;��S�1=���;a�8�T�|�0+e�_���yV>��ϠV�#����}�]v>p��p��𮿽��~Z�	lذ�DoټO<����r�v�Rl�9���{�噽864��\�<��Ӹ��C��;w/��m,!�%�?��.��(�J�����;wl{���K�<D��׍z�p��^�
���Rٴ<���{�Zm���k(2�� 2fen���4^�{qԳ���Q��\f�+<�6�0�du�.��p8j��/<�F�|�a�� Ê���X�:��p���:a�O�lzF�~�D���@,E���U1;	ǚ�q��~^���E]$��x8C����
jV׃�	j�t�J�Y�!-n�UI4DO�Ti���x�w����O��*|�_��?�1::z��zlx+NX�TjJ6�j�"��I	ad�CĢ	%�Z�J�KƒjL��㥂|�Nn�k��h$"J�D�V�+X�1d:�c쥩�բ" ��� ��ƙv��(I�âg�Y-�
��A6=�k���G���Ǖ}�6�>!r�^]O a|bTԛ<\�yz����hƶ υ=bD����Ė�RyV���<~8:�"��������9>"D3xP��Q����sK�+�WV]���\�i�K�_��\A�����B$�R!�M���� ��]������S����|^ą�������$[�G�&��R0�fp���M[F-�X8\V��X%	s��(/�v
�S�3����<���(Э���^��suWj��u"�0�� ��[7l/���tK����7k^���Ϝ��"�i(r�b�{�D��E�OuƊ �*����2wol�ĝ������p���^��(��
^�cz���v�ט���Pc! HP��Da2�k|    IDAT�������J��%��cφJ�Ԝ�����1����D�h���ӝ�{��Z��c�D4K���#��f��ܚF��?�	+{���3ؽu�y��(��&fgom�}?�v�܋�=�v�>�ѩ�&��[��r]�5��j�2"� ZA��T�T{ıc��DڹX���M�/<�|.�E��H���A�M?R�Gѻl1V,��֭O��x���7��n�go�ÃCx˛�$$�����U�p��>��O���k߅�����{�/��|�y���O�٭{q���h� r�:>N�����,����/���F�_��3�/���Xv��c#C�P8(��u���te������V �R��ZU0�W:b��\�����0���d����G� <�z��`�f���I�h^�h����!-_�V�4l����X�3�x�zîTju�g�Z�O���D����$�6�}���*e�P�CC<�9J� eY�ʼ�$�#��@1���]np����?��5��G>���F�J�<��E�����]`e�/�ڣ�����\V��d2�����sq��&��~��������=/�}��b�Nx��y��g�u���o�{�g������%��-.X�
��~+��t�>��<7�pxK%�s�3��ș�-��H�I�u�$��8����3�!�̦F:�&�/@��G&=��O>S��D[k�B^�_�h��$i`���&�JdEHd������&�*}��e�vn`���y,T���)�ܩ��#㸊�b&��/ĹՐ�H6?��N������RMi糅��Ǥ����OMNI_���5��U�_(�x\>�}��h<���$-Z$�$ꑳQa����T**A�|���A[G�����i�!�[ԧ6EģVq�euӃ����=�b���*��W�B�7I�L��IF�y
!r�T����;�ꀣ{�����
��Cn���E���ϲ;�X���&��=Vˑ4���	"i�t ���1�K�ˍ���H���N;�u�T�̀=Gvsp��+�~�ﺌ;H��w�]:�M��R�q�WĢ���������<��I��[~0[|\�"��c&=�L텤���ߐ�"^����}�8�C��8Bbj�]%�����I?���	W��
�^E-
J �f&p��'�s���gl���Qڳw}�vԽUQB�Ǣ�>\���كo~�x~�^�2eLd+�[�N���/�eؕ���8���IepE�Q&��l��Ц��Y@B!����pR&tض4l�x���l��0xd���w⪫.�{��g�z�'��;�oA�-[��W]�7������k���d���ނ���*z�:���?��A��(�-�k^V��9*첫��c2�֬��";x�`�mۑ%K:+��	�eE`UO�V��zR��Ql�iF�Uz���eˑZ2�l�Z���
ǡ��h�ʟː"�O�\��m
J���}>_�Ѩ6�Qm�X�4۶�J�f��gؼ��6s�o��F|egN�r�sE
s�����
�K��֫��3���}�?�]���F<B[2)dfc�]�b7*�B�M("@�"��[6#��#������d��d���h�tF<���^ր��>���r�и�}p��Z�!U��O�~5G2�	a��w)�._��Ͽ�����[?'�w:5)7�}-T���:W���:�Cy<LbHȢ��sj�+���WV$=J�L���g�� �VnlDb�0�E�NlS�
�'9��.:�G���H��(Ꙗ�=�xo}˛��ǑC��Ν��V�e��L�%�¾���eqƙ�`���|�n�:y�v�؁�N;k׮�?��T꧞z*��>9���?{�����6�|:�,^�#Gзx1�862��=�$R�<��ؾ �V�O�e��{���hxY�)�=nx�,ɂ�����9�m�[�T����*�\&�EmmH�c���N��#���[23��MD�����$p�ȱ8 �h���$�Ĩ���\�� W`PA�/�rڵz<uA�xߔ}MZiZB��U�z��V�J�N,�c���] m���p˱���]�.������V�;{�2��|��tݽ��W�bd�պjj����ؚ�kb"�M��2y����j���_m$��fW@WCps,y���	�|�qZL�4�H&�B�k	��)Pm��,�/�`�R3��Y(g( qjd��ًfS)x&zzzd�GQ��-H�&��R����ɂH�d�E�t&�ݥ(�gR������-~#I��vMi��$�P�	Ǉ�a�PD4B�21:x�0.<�4��u����h��G��C͠"\�pX��U+��_���<��D�,Z�e�P�����鑪�݈�&�q9�x$.<�d�Sa{�H���9Ba2���jqv�m���H�C�f�p��^��\{5n��ø��_����e�����{�p�9�a��m�R}�?�G����q�ߊ�;v�O>�<�{��]�{�ȕ��c(�l��1�d��*��_�a���߈8�����>��z���(,�NL������>����/��m�pL�1|�ggR0�T
Yy �(��{����ig338봓q�i'c���8�o���uu����yFf��?����enB���{��������
�p��ad3�/��݋C�ajbRT�֭Z!�LL.��=t�.��0XLN���&0��!�hSs��:�n߆}��ɆLș_|�����c�ҥȧ&�+�7(n�D�l3٬^B���3�qB<���T8͵�����XS-��y:�F�XE�,�3��9p ���%�D<�5��avzZ���=�3���?�1֯_����z�y睘�����g<��Sҏ"S55=�o|����p�I'��ۿ*��u�]��|�;طo��nϞ=�����5��~����ÿE._D<�"������U$	�0L�X�FbI���$S(���ȕ��aH�Rf�
vtX�|us�����X������8|�
¦=]����������S"�I���_�jx���=6�#GF1>Q@�PԠg�bE�\@��
��- ��
���/!
#�3�����f�˦���`,Ҥ�sB���0s�̖
2U�r��
�Z�S��~	W�Y��QyQ�������9V8�,�]vؤ�4Kd��i�=����Q�$�B��VK�E��7�Ri	����5�������w����4��h�&�z��\iū�Q]��lQQǀJ�uV�0�D�N�����_�1�����%����NT��"J�g7.�+�ТcD;Ԭ���%������2���1ARZ*]�BA�"��˨҈Y&��ZcA5fgyQ��Q��u��;[U�b3�9��m��Ht��
Ej�x�{%���V"�����hr($�!�a������N��5J�Ve��38��"n���o��������n�?a-����/� �|�?
���?�я𖷼	׾�Z����q�o�-��~��aXQbm(V}�4,�XiFe�I	�'���	&��l����?��o�}$�h���o��ÿ��W�B��=_(�IR�7��m]�]��K��p|��J��^Ɗ%}8���0����El���ضm+ҙɬ"�0*�:V�^��֠sQ���S������Ü�SK[��݄(�ϑhU4!�Z�J�)�ϬP��#��ܬ�(�ך�N�� ��`tl�JUHl|�	�3k���M���̛�0��9N�|>̹tJ~����4����R���#�F5$�V��C�!�����Nx��@�+sj�3P�I��"T,��T�h|~!�����)WLO����X�ՁW_�*�^�
�����~�	��Dp��M7݄/}�Kشin��6�!�����\�٥�t+V��{�D넍��,�Tj�\^�ed��g�¡~>mj��൧�� ���i �*�c�@��c[��\�Q�"��MMUP|<(�-|���E,E><���h�X���G���c"D�Z��9�����x���x�oơ��8ҟ�l�+D׸q�L�
Y��}	�-�#�|N͙{}5�[E��QĈ�˸�r�z�̴#��{Pz���ȩ`rƪ�L��5zu���Jz� ���I��9n�b�!�l�tsiF�iǜ�x��f������A�
RM����yGOCF'�tT���Ɉn���K084�0��!��$�1;�((�������1��jg|��r�ys�L�4�2E���;����Hb+�V(I_�2-	b7iӕ�3���"W�=D�7��r8��k|���<G�*x������/�3��͆$�l�QL��1�|�,j�[��e1�VE~vZ��z�!#�H5d?K�[dޛ�7�h�/�,�;/|���RہS2}RTJI��x�<:�q|�W�:��'�����	4�p䛵J8`�?��y�[Ձ|�^<�⋷ނV�g�lyj���N?�L�̹�o~z�<�l��v9�p>r����ݩ6,��^���h�a���(�"�?d��~&��}z��������v�>�-������M��ǁJ3��]jz3(3��MX��BLD�hK�p�i'������{��Gd�KVmwON8�D�Y{�'g�|��<����VU�@4��%{��Y�0+��Rl�E�7~q���%�`�y�`�XY �t&�{Z���z\+��7��HvJ��8 ��~(g��Ĩ�F�>ǖ����w�h'�_�� ��Y��K�p��B���L$ZT�^�J�;��O�j|�'�=F�G���A_w��yx�_|qN;��a=���X�l���GG�%�)�[~ԔCD���W���E�2�� 2ż��t0A����6���ZjT���!��M��h�3at�}kU�+R�,�%��T�����VqIԲ�x�%g�#��K��u�L���Na����O��D<&�.M�j�\x�؇��^�L>��^}5B�.<���A��#�� �����8�s��_>�ǟ؎F�~��2�e8�Jo�p�0�4S~*f�2���.,_��kز�Go��5�~�����u�za�-�K��E��w�u6���{��e���R�/�w�sx/�%u��Y�+D���XN\�g&��Ab�,N9�\|�y���Vl�;,'$u����Tk$��U �}��؛�r�I��ʜAJW�z��x�f��19]�+��!҂hPYУ�{�u�
�/�lSX!>�^�+�����b���$�dz,�M�N��:q�>�>�U���d]GPk��Xǃj�-H"��Hjf�Т<������~yV��=fZ��>�h��41C��X��
,M+�h[;
6y�l��*7����-S�p(D�|)�Bf&��.��H��a�mQ� �T�	��ԍ' 4�At���Y��\p��(�ӢvI>y@g�u���{v��ʕ�����&'��X]�*��e�򩧷��w���,v�= �9�eS�U/����e�����''�/�sϵ�����S�Ŷl�,P�4$��e5ٯ���+R��E!���$ZcX�l1J�4�>�t?�ggd�S� ���E��[�������h?�	��ég�-�$$\)'/�WH�aS�@j6*�Ѣ�2�.r������g0B�P���|/>d���?O�sj����E�]�Y1ss]�b�T�|��!�Cx����?��"�n�>���/��l6C�W��:�j�_6�G8�?��8q��uFY-rޚɌ��92��w��=�I��d�"�g��x֫�����"J6��_,���;ω�I"ކ�[�K�?��_��ѩ���iҖ��%\E�殾eL�� �h�����(ں!���ăcq4+�J�FC�>���ϑI�P4��e�笠]i������9���t-��~}߽ظv9�.�ÖM��M�gۈ'bbiE"�p��He�x~�N��v��`<U�o�c<��8��3���^�l�N�~�o�4l;�z�(&UT�"|nʊ�M�z9��Q{֮Y-I�~g�$�c�Fg]t�y���b͍Sɳ�V3mB��!�W�	��M�~#�Z<Z��-���:3���E�J���	�˧��"�I��,M&�R�E�~̤F�jy/n���C4�?�b`tFxu���W�O'���;KSח
�sJs�_����Ά�usD>�jV����>��8z�l�Uף�����H'HH�f��GmY{\�k"B%=tuĚ� c��^�bIf;��&zUU
��"V����a���-�}dAd�,���ut��P"Z&4�d�pf;S�Y��ȵ��aR��?�G[;0�ck��	�S�M�B�+Ā���d�s�i�)�_u����}�\+xՅ��-��K��Ϧ�E��>�B>�d4,�C�hD
GV��PD%5-d����WLhZ;�8p��&&��K���,��;���F�m3�,G()�	��o���QA�cc����_��S[���@�A˹JA�#}&5&�/���R�B^���d�r��(�<	qo��R��Űg��8��h4(��l���]z����@2$V���c���bwJFt(u���je^�FPHZ�/))�uW4���Ư��H	��2�ͨ/���E3���i�QL����cy7����]�p������)�Ku�Z���O���"Ѥ�67h��#��8�C�t@�&�p��H�IH $�&I
�ㅁ�2w��P6�$ӷ�c@f89�Q%�q,_�TFԨ˾~�LNL��ƓO4�`)z���%��Ʂ5�9z������..gG��&�ZGE����q`e��K�ur��h�^!A�؇��o�	�*"z#���&9A]I^�0%l\҂���!�r�8 o#��x ��������
�9�ю���ٗ���ڃ��ێ��i�͵�i�q��o ���݆���j���.E�D��g>�+<��>��D_�Z���+��r� d'ga�*8��d�:tp/�y�ո��xz��~�7���� ���D��E��x��(�U�ǍZ���l���ȳ���)5���f��`��S�9�&��;|$���_ŴWϓFQ����1~(Ĭ���������Eh�VB4@8N� :�ίނָy᳷=�Ƕl� � αM��UB�A�Ӣ#��u.ϒK�F?ǹܨ�<��9?A��u�`�ǃ���1�%Ϛ�\x,<^u�� �V����ޚ�Λ)��(���s�S�����sP�*lp��ҳ3�o�D�X�E!=��z�_��+/F��i����g�a���&��b���^!����>�*0�Q����j	�B5/�OA�i�Q%� e_��6��eՀQep��$��d�=��
3d�Hg{��|(�5��;��m������o�(I��%����滻:��ךL8*�$:��$�B�����p�LD8b��!5;�(�qlp-���b _k ѹeÇ��)�#-0	x�!�C��O���=���~8�h��+w���'��T��:��j]�����Ը#�j�. �\��>��@����]���a�sݻQ)����G�x�tI����D+,+ �%�Valb
O?��T/�\�GG�1,���;Qڭ �9}JnG��&��'��	V{NP����	ѱ2���쏐!��TZ*�Ϗ�?�X$.3��!�ϥ�re>����u�������xj�3`���9�`nʼ�l���r�B�����	'm@*�X�
H
�d"��E%�-�9������j�1@s�kI$���SP�ެ^�Ft���Fd�������!���vczr
�d�x�d��rM��<~�
��%)Ef�nO�?�TfB.R�T�8
H6w�X�w�]������12���r,��*B�|?njܸ�����	��*v�8��%��u��!�w�wp��pډ+���¢w2<n4 S�q�ů���,�۶�_���W�v�8��ۂ����ꦅk��Z�|�R��xj�s�L���Q����H�0�����c+gr�����]r�x������ox?��"�;������?���LMga�ыbXs�MXd���Ɨ�RU�*���̙Wޟ�    IDATI���V�^/�;v�:��`���GdԺ�D0wB0'�:?�Z�y�%�΅#��0Dp(Mn�߃@�D0��h����7�Mox^�}߹�7��PNbH��hy�k�<����)��&��mv<?y�79'G�C���I��������Ww@�kI�0��L��f`��c>3O0�!��E�	5�H(�w�0h���ͤQ��dȃu�1��4n���X�Mt�ՃO 1@ο��O<�g�ۃ\��5'LB�d����eA�̔L~?���rL�I���EP�U�g%oz|�>9�\�>_�!hX�j��q����
�"����kv	a���� �/�Ɵ����L�'��{�mE{,�V��Gd���s�Q;�KY �:�K�� ���T�'�}�yz���#����9
����X;�4梔�7 _��2�1��������yos��|�{����;?�/bQ�܀�fK@7}	�"^I"I�@1�A(��]+K�K�\-q��)]��%�� W���ē�!h)H|dd�!��V�?t�}�Q=&A�Vk W� � %Q��!M������I��O/TW@wU鲐�3@`�K���y$ے�PN�̱����i��v�i�Z�#3K�qK>��5#�e��p������ؼ������022�H�=D�+�j�]�Z�	�ƙ-��RJ˶��I�Lg#��s����<��c���jF�BGI��Z�����>tkKB��S���۰a�����#	ه0<� �mg�;kA�R�'B�<hE�
D%+(cDf��*�+�[*yQ-t�NM�ȅ�T)D��ή.i-�0E M�kJ�Aw��޹h(p��Qº�\y٫�����M�`Ws�=:�	[�<"� �|�>t-_��T�w�ǋ��7|
�>�4��v ���hA��(�	�7�"[,�2))�d�U˃6�&l�b�BJ��j�L���i'��b!�����}�d�zJ��_��#�}�h/ҳ���M�@&������dNU�^�r*Tu�й1/��ͱ���pyE��7]��sW�rO����p�Q-B���3��乤3���'Ǖ�5�ֶ��ǐl����\'������%�&��I����ה��U�7G(�9)����	׹�����&L|�lhޔA�[���6#I��S�kֺ{:@��ȍa@%І
�E�AJYu�ꉣ^��5�z'.��\:t��D��}��>�D�N�UP�� s]^>�4��%�f8������,�јU#�#��^Ip��r�Y,�**��`��V_�B�dH_!�������Q|�k�c������H��%�BHea�J�@�;
��'����A�8��՞���L��Դ�A�5��N�����n��{ѳr-�&a��̀�slo�#��Y����{���S�?�/=�B'q25�annjE�\m-!9�(��Ge|����\
��Y�g�q���X�ƢqQ �8����ȋr�wpp�/(A�cټ!2֠�\�@����>?�v�g�����LV5i����g3R͋��L*-�4��9rza��(������)��L��e�nblR���c�d�e&i���`\S�f��y�eRf�I�ы9��/=�p$.����k��/�0Ûe6)�����\#��0RXE*�xK�-	ޱ�QlذQ��d��ߧƩ�Xp�T��6q*"���^���f���Ju���K64B���`zT%�����0̙<4�JDkIq�)8�@F��E�=�<8>5��lZF`$�	;�14i�W4D�)����u��,�����q`�n����� Z��)cljR����Ä�
Ἃ_��v���,7�vJ�k�
��R�J�L���}�S~��&���4�� ��<��%k$���6!���9l8q5�;�L:| /�܋ٙ<F�gQ)Ta�/�h��P4$��6��?�`eN$T��9��c7�.��<�P�w���)�.I�4��������E����ދ�,o�O$5��I����� �B��D<��A���1_ .SLf)H�$O�|���=u�M?���zLO!^���x���"9/�[�eO�mT�t�	\O�f^�TZ�e�T����~˹��\�.e�㛣r�>�ڿt@7��	�2Ӝ6�Q-�Df�S+�3��dK'���m͍��;���T^\}>N(G�HD��ن�d?qHn�A
�}p�B~�r_,�
��uU����S&����⚯TD��h�gg�a�R��?�+��>�#/�Fjb��2Q���:�|&�B��T��c��tK�lb���صc�� Z�*g6���[��w�2�+6���!_3p����s/��hg<�4$��F?�W�����W���q��~�eۧ�eoo�JI�"���TI�����X"(Z̦��q���ى�Z�&ջ�c����x�8Y���v�UrQ�m��-��eQȗ�5�8�W��ȕ��<Ǥ3���e�fq���`�I�R�.p.y6�S�5^�Y�����i��G.3+=��+�"1N�qt�"ҷ�T�V��^�C�7lP�}�:���SA�Z���K���]j���$!N@'dO��V��j�=��K%���^]��T��GG���'�~�أJ�i
c�5���/��z��V��9�[�eM�_z�$J4�k4��*�vz��+��h~̺��̝3�c��͖�Ix�U ��}}D���@z&�$���r��dBP ��2b�:�4�3�����V�$Ԅ�{0��B��92w��<��,3�
f
6��<��oācS0�	8��9����7d��y����Sz��,��j�u�u(~�(RE���6������E��HX���3�g����]��AWDP��2�+�����Н��#��e �I�[��%�8�s�?���!f�y��0�]͐q(��E��yt����d18>"R����Ƒ�hW�Ω��S�B7[9�J9���i��$���m'X�xeO���&T0WI��B<J�mQv���_/ii���
�;}Mej߹n��8}�Φ8��/}��ʅ���x��0G%ޕ�,�v�:�����}v2E��,|�#�p��?�t��I�0E2a;	��(��m�h�d�L�E&�X�/�B"_,����P���x""W)�T(
��p*t����C{��nF[��o��elX��~���?r��=29�}�~d,`ۏו{��
P\���i�[J;r�����)yC9Gd��!f ɎE8pd�@�\��>tE��`k7j>�h�c#�l4�ߺ�?t�O�jfo���{��ɩQ	"��m��$مf$K�@�11z�3X��C~�_�l	�y5?�M>���$�pL qn��r�GhE�����T�čN������s��Rي��^x���HFu�4h����-K�� �1�"� ���'���jE�eh���]X*��\��qA��-�Ϥ�
X�uo�1%!�i���P��ˬ7f�Z����ב<&jS���l!:ϝ��c��v��J�=6>���qtuvKR%�q����a,_�5V�P.u����Z;�05�������M���%��$�\��u�Vw#�/����|YF�m�_���i2�"�B�orrZ�Bx������ڱ^���吷�*�ItƣHZ!�*a$A��F"���=(�3>"&\�ӂ���ImI4�����;N��/����	7)�Kn���z�BbU�M��k4����<ޡ�AĒ�6b���O67+h	7.�6�7������ϙt
�dR�@��3*�mڐjU~'b���:���ϵ7������&�����47�/��_
	S_���H�3����Z�G��O���t���C���>?�+�DK�RA�1�J�^%�T�ˉ�3g�|o�9��T��m�$��n����
�e	�*���,������q�c��s];w����ڪQqFh������A������-eaԲ�\WQ����Վ��Cb&n�FKK��~�mC
"U�5�@zKDQ,�P��aӳC�^qB$�_��׃�~ZW�Ж�\!S,O?��sa�G���nr]��C&J�4L;�O�����w��O��]�f�H&b��Az�ƍ��?,�c��>l߾]� �F�+�9������wxh�Q!`��Ղ:r$.�V�b;������-m&�0S���/E��Q�J#��ۧ�����W���Ѱ�㞷�~��ϔj��:z������S�J���C%[C�h���G\��86|H��HVI#V%���%�z�G6C����EX�yqC��*o��J����1�[�M���*iGw��	q���p��^��SLa&&�eSi�h�M���X(����abdѠ%���(��s�AB�R��kq`R���A��,x��A�%���D��F>aVf��.�##ajTO���[e�����E@�^L!�-%+�k)b5e����q��u�g���^��.ے,7�6%�z�	!��!BM�	�!$�f&!bB7� �c0n�n��w�������Ȳ�03y뽵�e[��{���Ww�6{C]�
�$o�����O��t<�jj��&`�kUު�v�$��uF��jA0�/� C4�If�0���fG*Wc�^�1,&Ȋ��~���''��C����`������.��`�XU)f��sb���� �D��fˌFʓ�����iE����ذ$Xj���D��No#ƣ�M��[�D��$�	���og2I.�	��lJ���v�	����� �ѐ�q�+&x�u4�B(¯Ջ�5���x\.DCqXE�7�E���qJD�-�cX�f�%tu�w�U�V	}�D[M���yXK�=K���]���'M�gz����5`W'�
�١ڛ�h�F�b\pD�1*����"��l����t�@/j��
���N����@5����w��Y���Y,�+|��m���2�����	�����&����bf�n���'���ּQ�_�jq$�fU����5��i�t�E��.]$�qK�J��!	8��Kd�)�lu�鮁�߄tJ��]W�I�	��&���N��N�X*�x��$O{�Βz�G.���5D�N4��@ۜ�`�V�bI��lF��,�=�*(��F:>���,�h���o�o�#��`3��b�<���Dz���^·��m\z�%ذa�`+(z����?5~g��,����ِUD ����._�~��E<�3���^����x4��:�#���sԢdR	��j�΄��]?����)gܕS�	��Ptr�j1�I�7����=�j�a��>&�[/��l���	<���i
�SU>^v$�Oe�.|TQW��`J�Y!�w�LV�<t�xT�T{ ��D�ϫ !A�R�ۥВ� ���Ĥ��B�	�d�b_>�l�q��Xrߟ�c�z�(�&pY-Ĩ	ԋj���!dE̝7�rE�јз8N��^a�D���v���ѐ$B�����a����R9�@J���S�֤h{��I�z����j�d�}��K�����-v%=j��h�s�<)�x/�s���IT�����KY��ě���U���>��7
�O��r9�S	�
4�H�Do0!�L#g�huJ!AQ�h�8���T�>.k�"waf�n7��� 爻i�3���X�`�>�T���attFC]�����:�--�ƭ[�,bf[;�7ry&�)4��Ŏ��{���F����X!�ՎR�;B�l�cxpD�Q�:,hC(8�pd��yl۶;w�cb2�4��u��SU�׏�6������\��Τ� <��;;��L�&0�۫��d�]|*4h�H�b+�	]KBZq;5�-I��R�+�"y�(^��t�G&:pQ���K=�"��������g9�N�q�L�C愄�,�`�Ӡ�����<�JJ4��:"�$5ʜ�����)��t��H�:������<>U%�sz�g�B�'�%���������>�H���u����I�ڸzB�*��&j�D�t��ʏ��d*�t&����"��m���A*�G�@�e����g�On{!�@ht5.�N��q�nG�,�TR��e�P��,O�p�y�V'J&�Pkm��&�T>W  ��x"�Tt�\��=�������:�ɴ�6\x�IB���q�W�<�ڵk�x�}�����n�.'�JP�XJ����ܝz꩒���~w�m��O��7/\x��`�8�h휏-�=�xH�m��)��<��J�J��û���Ɗ7���E�Kr��`K�+�(&ݒ	�H�Z��u+��tiY�l�4`�!O�Q�͙����P��|E��Y�M
�Q�U�7��!MH�/¢��@-�C)�ꞯQ�Wr��Zr��q�]=8bP�����/����D"��'�o|��HF&���\
ۻ6�m֣�jC&�D,�����S��т��Qĳ9,>�3�����;{P2X`"e����DN����\�c�s��?�1�{z�Zݺ�K����s�kCmm���=c��Vh�p0"	�� ����W_-��e˖axpP�y���L@:;;�����)������=�%�M���yW^�2"�T�}NV�Y���vH!��>[
���~�j���ٕW�opKz3fcێ�vٛsZ2>>*�����.r��pD@f� N8�hR)l\��Z$�1C��FیF��˟af����w;��"J�8vnZ��'��}^���u�\��%<��K���g}ɔo�؈��{00�+P�]�X,��"���L��2j��M�`5۰�^s`��c�:\v��q�g����v��x��Q��@�b%,��q3�2��4fI�XQFE��0���E�1y�����{M���$*�:܅��r�V�B�������.m�>]�mW�����`Ю��V�Yv�6|�*~
9��I�	�L&?�R�6�?B�!�"�)���a���	j��M,�t��.4�
�|��A���(�MFB���"����/-�X�.�2l�������{`v��G�������&	�� PqOh������ǰ��a��kO��.@��pJ�	���h�r�yuX��'�`����ņ��1<�SVT�d
���
�x_;��.�.l���+�A���s��Jő��+����\>	��麫����k�.�+/<��͛E�9G݁R�￟ġ'�z>���n�E�x�g��s��3B�;e�)� �r�~��_�������}A�m[�a����˯��g�C��yp0#Q�A��V�mYs}���;<�Un)�\m�xȗa1m^�dhL���*���պ��`#A�����n��N9��J�`U�D��hi^h/�F�b1ZQ��p��RmV���a��Z�$�D�v93Qю_ϛ͛�џ�(��銦v����I���:m˾䎓����F��8.������n�rtoew^���~�y�4�̨��#�/b,�̹���>��(�t��E�A�d����|�p��|��a� ���M�p����G:�U+Wb���dk�iFm�N����ME�YF�4��PO�$��T� 3D���_�!����^D�Ay�۷v��$茒��Z��	'� Ҥ윹���¶���E#q̝;_<�<t�^���ÃK��'u��並�c���ґ�!ݸy�Ο/ԯ��a�6w �,���E�*�͊;_;tj3��A��!I���G9�F���8��c��$�\���fQ.\�p>����S9C����/F:<�������劼O�Ǉ�?��ߵ�֮G,��W��M�
f<��[X���݂�� w�E�q�˳l4�P*r��Z�w�f. ���;~�DBa6lچ����"��9�1W9�z���N_�z��D���%J�*��hIѕL&Il��%�\(}42�q��mO����t���s�>=�(ʴD�������jW�# -���b�
���%���)����*����z�YVl\�qm��Q��=i�f��Y��(Z*���nJ��?Y˴D^�5����������AL�h��)�A$���(���_���ׄ��I�&���t�:��R�T��U�?�h��*Q.�}�G�-(&�B2d�ػ�	�w���w�����02    IDAT��7ȹ��<�\}n֯߄Ɩp��X�y ϼ�%�:j���0���S0:\�)/��c���K1oF ��<�֯�sO>-t�D$*q���E�s�w.�X~&�]��<�tiU|F�2�~���%2y��������_v�E��ٍ���8��sp�a���jP7c&ƣI���k�CW�
���.�����3�xo�o�p�'�Y#�>�PdR:CA'�|�]�=<h��	��w1�k�L�D��n��7�I��ո]��B�}�lNLU(/�.'��f2u�9��Eu⒀MV�N֒� ū�~14(��_�І�^��X"�~�^/��JqL�5�� �;������זaǖupS�xr��:�^�sYd���z��g�9�7lD�d����M�57�+_��5	!ɀXkJ+��V��u���o�+�3^x���G���+�s�E:gϕ}"������{�v�J,�7_:kʮ��b���������'������n��H���7+���`o,Y�~=/^�/����2`�B�b��wW`��nI�g�q�{�4G���6`t�_(�D���b$����M�VV�˗/��>�E��q�����`g��E �+ad�2�̘5S%�� �L����;�B�C���#��ـ˷aɒ�����ŕ���[�6�XIc�� �vlF��`��`�_��,z��~��������q\��kQ�Xq�/�ƫo�G��C,_BKG�"��Q��O�N����-�I٫`FK3z�s8�����N�����CCaĒ��1��T�>�.����x�*yA�<R�!%��_���9�Ó���)�I����P��^0$SNj]�]:U�R�Y-�wO�'�=��t��+�p7^L'a��"���"畆!,��<�F5m�z�y9�L"O˞�S z۳�b1C��ádS��M¥�~�{1y�&��I�D�E����(��͜�q�D�Eu?49�{���y���X�.+�O��f:�M�������z�{��ZR���b�L��.0%��`n�EueQh�%�@&�}�᢯����`nG�(J�@'G>�b	�k�N|�~'���p�w����~XZf��)Q1��6]%�{�:-.�Dl�˞}���m� �>��_�Z8\vwwW�mF1��D�ȹ��#�q���<�m�q�q��\���N�׋��?N�gG�l4���K/�h(�dA�}���4��B��w��8���u�����𙯮����hV�?�@x�xH�4�h���XFCV3`c5���n3KW����	V�N(�!;Z��M=l���5�!<j����"�_����L&��~ٷ���n��P�4� 0�v��qGL�2�0`���?3p�c��ˋ�kE,�����S	��69�O�����7]��^y��8~'�}�u���d5#ϑ�ɆX���9�1�����`"�ı'������w(T������HR�I�#;�L��������D(8�|:��^}EW�z��с��N�&,XD��h���k?��t����h���[n����<p?6oވ��m�45�k�����El\�3���!y����_�o���̝'כ{�D2�W_}#����K��#��x����\(�S�u̞��.�הּ�(FF����
W���>��9���%�7�㵷Wc0C� �L�dM��V��.ǘ�4s2a5arx7���1on-6`�q���_�s�L�p���Nd�a�j*i��<l}��*�AĨ��_����a�Î���ql�ُ�����_:Mm���G�ʛ�l����-�0<1�	��ѩ-L��a(�i�	����k�sO�(aDc)����z5NI����t��R"�IR��A[���VC�H��c6KG�&"�P�1��k&$�TqǮ�Ego��	}*iL%��9OO��%O���4��v#
!��^�kYuy�h�1C��T6�'3�.�u	v1�	���$3��Ci������,��L|�nS���M�qK4M��4QG�W!��k���)k��oχ|IM\��+A�_M��iӓ���=)�mH�j�R�i�����!&V4���ԋB5�N�d��(N9������0���bݚ�2-�8���E����͗�ѹ/V�݆m�A��ڇ�Ӈ<�7����ĥ\���GN��$�C���G�ϊ�����yo���RdK�|�f�[,"�E�&',,�?��_�LT�:�����5���rME�.��흈Dc��3�W�9�,D�T�d<����Ӊr���u�<v��+�ݖ�8;�<�Z�I� ����ND��+fQ+*��ړ��lD]��:9qۡ���	�<v�Sv�D s �L�f�d0'
������s�N䫗�:������5��@&����H���:1-�$�B��A^k�,t)�O�{rb���Ϥ�5�{�p�4��丘	��Q�/����-X�v#y�Y��E{s,^�LvĲ9��D���x�&�p�`���%�x�Wa0ڐH34bd,�@��8*�4�j\��O�E]���X��=DCA���xƌYR�8���N�l���\̯��`wz�����ߵ}~�Q�ܹ/���^�W]y%?�p˱���c��k�n���6l����ǎ�^C1��OH}�w.��9}�#شn=��f�����Z�l�(\Nv�6�Y�^{uV�Z�c�;u-�����a�����k�`��~�j�14���:s��j�Bj�/��TD>����m8��������O"G,:��.�6?�3X��-��AG{3
� �֮�!�:�0S��T��'��X��[��;{�/}���c	����1{���X��S�+8�+����ēK�E�*T��#�=/t��G#m	��� B�k:CJ��^Ą��ұȥ���82W�:��j9�v�b�j����^���U��$p"�iФw�{�R�S 6�O.@PMȤ������N%���	G���� �=!���\>#����5�>H����(���������j�ȸ�bG"�T-�Gz&��G��Q}1��R������2�$r�t4�!����@2I���h�����q���o&�=h�(1W߇6Q�5vP�p���7���"�!;r��8%\������k6i�D�T�vn��B��9��	����A�GI�,V#^z��z�as5�?<��=�2ʵ�(r�Z(
x�D�P�̸
a�u��F�������X��K����BB�夔�<�7@�)�mpG�u)�2ݨd)I�l!b�
y��۠���&͍`�
\�E��ގ9�J�P4۠�٥C�yIU��7K��i��%���b�o���x,�J���"������>��R	�P�P�s�+_>5^;m9�Z�[6����&Ó2f�q/���N%���ǨF��3g��DX�i;���F��K�U���MVZ�M��+��\NF�<��͗�*��/`}E���0��߲Ï'��H���>�\y�Eذ~-vtm��b���?�Es;ᰑڥ��Ct7*�e�|̱�b��yX�r���cpy(�͘�[lS�~'=׷�1P�k�):`r�V���c#���⅋0o�\E'�N:���c�v9�s�t��"б����sG��^Z����W_[�ǅY3g��o_��;n�K�s�Ʉ��V`|tw�u���B�d�:��������d�q�%���߾ �7mG_�N�������ܯ�ԄF.�xL�$�L������<��
:l�:�s���k�*���vK�|8#����$t�g��5��̀��wO�M&��~W]v	<^[��xn�:��o[t�^{�M1����g�����U��߿�W����0
�Y���Y���]zD�P�6m
�w�݅��Q�:��.�2Y�d��^�����<��ƙ�WAm����^�1��)(�p6�Q�ߚ�V�"��.'T��Yf�F<�8x���D���s�	��h���3���J����m_��~�nÇF��q�|�i��u�;l�{�2� Z�A�gT���q�����/�E��Lz��� L��!�4��"
>�v�t�2RW6"�[B���S�_CلB&�l2���z�~���w�^x衇�a�v�RF�L��5A�qs��~a��T��������^���j�bkZB�)�l�	�+K/���I:d�a$�#8꠽�n�ho
� ^�P��
(���Q45�a<Ļ+7`�^b$X���=C]Jz#�Œ�Z���X��(���0!>9G%�cZ�_��j���?㡿-A=Ņ�a���rE���.|;l8���8^��кsyo�����W�t�~�Ͱ b~������@�PB^gB�lF,W���Ҹ�� ͧ����O���������PL�P�gP.�Q1���*�\�����m�!�
��·믿V�r���c�T"-7��d�6��169&;V�����ŋ/;lqp�!P߀��L�bx��G�j�&�N�@�O�BF�G�ɧ$��ޥ�dLμ��S�y���J%u����D��R��ay�L�v;]�x(-��L���_,	k�uh���`_?��[DI,��at,(��s��x��;%��Uk�kB�hG(����E�Aҏ�����|�\���xz�cx�����A��Yhmn����Z7��`P�o�K=��3`w�����cǎp��.�o���@&'Feձ��(�e�|�]?ȱ�+I���>_ .��Lo.G~ց��_��&8lV���)�s�� :fw�}v�$�`(��~�u��{G^��sro?�hl�9��X��o���,#Jq6�u��b�	GCQ���/WP���� j<^���L�P��F]��h��p<��!&B#شy-"��t���<^_�26lZ/*tF���q6�8��شa����|s�ar��hm���(���q+\n3����u;�_���������}��Z_��HN���X�PC���)1�a�Z2*���IXbFĂ�^x=��016.��?:
��j0$kE�`��y��g�KM��_�2'���J`�CW&��� 8�7���U w4�o�׵Ⱦ�@J��<EOH���h����Z�.������,WE�ST�#�c�沲�^�^�vK�ӵЙ�(����w�J>�����|�d4Գ�n��OX�j̶a�Ʋ� �ŀ\�s�=����?}ǭ�jԇ֙k���:�):b��ѷ��v{�=���t�ܔ�f�}r����M@	Yt�&�A�L,S%���Z��߀�D��=�P(�y���%�9��`F�,�^�	�Wm��D}I$�6��(w��C���f1-Z�6�ؑ�.�����S���'��c6}�m,��΢h�Z,�Y0hU~�Sb:Or�J
ig�{.X�8�I�1o�<446cݦ���H��0��H����oAIg6	�[�ʴ�pl��}��y�7Vn��gg<���B iv�q��*[G@_,:�=4����~۶��ͤ�X�$�Lxደو"�dk8�����Ft2$	��/Ip�M�����m�d>>��'�,b� �

�Zf����.7��^�����&���Ƃ�����$�qLg2 �
���Mv���Љ�l��i������ ��BƠm�[dDĠ�qy�3e�/�i�l�C���C26��D�.[��8m��I��T"���f4��_>g�z�oلg�Y�\�\��۪Կ�tx�y��e�h�hᖷ�~G����A:��~�+X�vV,[t��I����|l�fϞ-v�,�Y看+V��w�Pm�X���j�T��^��|�$�G��c�!�"/��ڀ��X uo�9�^��٣�A��yx��wM���c`�����煶�:S�Ո���FqX̂%�x��2h��h4�����Մ���\o/9ͦ
��	��,�7�;�cdl��M0K�M!��JGI�fN�j�Q�4C@Yc�a}�����E_��K���xF�]��啨�f䮐�I�)s�bI'��g��Uep��}��"�kz�=Ȗ��e��3q{��s0��\2P��3K ��g�ə�<V�dom���/G��<��t�S��*Aj#tM����[�S S%̟W,䠓�75蝢!ο+抂�)pM�"��%���+����-ʺ�#xN й������ԮoC�f�.E��ҩEA�=r�,ЗL(3���8��q��G����n�q	�_�݈$s��Й�Y���>�3*�Х ���5�=#��8����?I蒬����U��V�U�yvK�:!RJ�ى�;��_��m��b�#0sF;��G��g����+Q�87����?B��F������8f/������ۆtt3�݈��a�k3�8�X��ؼ���*�x�Q��0f	X�H:�Nb,φL��#eS|�Ͳ�*��(����3]�`�I��:Dֻ��#��z�jj1:��[g�U�6������%��ݹ�w��-_qu�n#h����K�y��ႾP��ͨ��fľ;�+/��O,A.��L:�o��L�"<���>Dbaٕ�k|r�M|u���M��Z�#KaѾ��e˱�Օ�kn��p��\^��?���X|@�1���=^{}9�M�d� �� ��Ռ�V�>�)J!V$�Л]����E܄��F-vlL�W�֑�V���3 ��U��9bd�g ��T� ����Њ���p@�o1f�jE�ߋ���`tdH��\)pr@}{���Zɭnnn�#��I�*(qRT����E
���@��a�&%TA�r��������Y8�k�\O�"��	v�abf��`|d۶mC,����١V	
L�p �;�Dtm�A���uuc�pA1�H144:$���&t/r�2z{�D����&��Y��)x��I%c�;�3m1���p؅IA�v�� ���o^��hE
^h2�Lvl�B�����4!�L��?�X��l1�`Goo/���_�\�35Z��5���Z��''¨�oT�EUqڣҗ��1))�s��P��,yk|�t%�Xpdn�O����HM���il1��`�;Q[G������gd�+�`{8���:��万+���?*���� ���hxS�����{�3 ��B헲RZ��N=�����D�[|���b)��H�(��F��P���1�؀�*�t|�ɷ&(�b��e����s�Y��Z��^}�HvO�񤨠��.���]����R���0���3~��۞I[��4�%�)-��ޕ��Ǉ� ��i/^ۡ��T�~�װ��M�t�$(�d���� ���]�m���i�y��li��Ą4_l|��9���2���V��B(����E�&+����F�� ˩M8AC���A���ފ#�g�y
2�0b���N9�|���L0>��"Q�,dWUA�J�@��7��j3&�'���sKq"Ơ�s��Ֆ�]��<'��{<��G�`��]�Ѧ��6�/ؕw.9�zo��ܝ�D�b��xB�Ռ�� L:J鬸����K�����_;cC;���P��d�)�.���#�I�󒄘0��g�㎑��b���_�!��y����BEg��w�㍷֡e�|ēe���Y��:�����3�O�>���w؝^X�iW�f���c�I|����<�st~cr��E���&�$	���A(GT�����OFK%&B�h��'�H��jR��e
�Z1��,G��f������L"
��}%�\"�x"�@�_I�r�Ja�B�A����6���8�f����$�I	�U�qA����D�3��p���/]��J�, �,��c�8:2���!474��� B&�ư}�qs�5g�pMFâ1O5�d���/Y��; ��W}#��L����0:2��
r��0�?�\��l:%��r)��<Fޣ��Ao(����X�K4�99�DS�b`h@����]��-��bN%NTD��b���Jaw{E`�� ���x�#ﴰ8�㾚'8�\T�h��J���"	��Z�`p�D^S�O:�i��?AmM���b�(���B�Ҟ����u�=�>�cId
Eq��p'BN���(�~�{hҭS��)�\u��q<�=�t�e �L��A���D&mA�Wg��    IDAT*S�^䕳cr�첂�'��a����pF��|�6�mQJ�y�Q��lV4@"��~�{b>���H�z�.����/�L���H��G@�é⊊rˏ�&D�W5�~������ZO����L�5}�D����Um_-�k�4�����������i��3����\N�瞌�W㥧a�%ׂ��<��?��:a��]����	����T:�I%j�a�9$��p�\΢�n������ࢯ~�x~)6� (@׿_��Hqf�A���x�	���<_u��ڦY��Y�$W�!���+",�N�]��c�cR-[�H�D�9-`��:�O(���:���L�9L�t�BF�h>�2�(f���� *r��y�b|�K���4 ��LN�UT�\�x��E���G}$����Յb�:jke\�Gѵm'�� �}o#^z�=�ۑ+�`q��;�q∣��瞃��w�޿< �lR^�����f�T��sy��V%��8�ȡ%��c$��M�e�I�+�5����@܅2��fU4p$<]�v�AU#Jm��1#wE�)���|�>7b��b S�$d�Y��)�AF�C&�E2���b���t&�5�+;x{�.�=�`kX\E����k@�v��<5`"�/d&c�:�.slL%�Y�3h���[#��`�L0�[�Q�Ҁd.���q��8��d
��\0Z]p��spTvY����624�r�  ;j��˝Eܜk���8���Bu�@I����;�� _7A��X�s;E�:����ͥ��o��0��T�Yo��bs�m�\�#�����d��zNm�JJ�òw�)�R���0L67��d9��������=�-��%<��@g=(my��2`���8K%��$��$���$8��
M�`���,��p8��'��+钨�v�*�j�����Z��aMv!,~�%{���p�^��+��(���	�ȸf��b�R�fa���DV;,.|6�Ԡt/qL$\�I� ���^ N��]N�x-��s���yY���!�V�,���mvd��O��-pɬ1QhE���غ*m���D�����1���?)�O�>{v�R~�`��i:{�A�?k�lb�Ǖ��i�-4��!����^@qT&�303�t�}�QHN`ś/��JL�=cb彌����X��`dRL��m�����ZB'��C#l��YavY16:�|$��.8�>^y�qtm� v�Q$��t&��Juu��4=�L��T�T�[����ؽ���)8:�D��sJ!���ONIˤs�M��4 k2a���Z�,>I�<K�΄~��'���w[�y��3	��^��$�o��F���0�&��3���%] })�\&$#z���wA*j�����I�s�l46�
���XI� 1p�yh�t�!t�ƪ5��� �*(.C�6���|?e>��9n�Moh�-qI�Ug(њ�,%9�}ŋ�0�3�U(�A�H2!��/8
��I���`N��諻�]cu�U}��D29�e��ʝ���t�9ᆢ�q�oHP�NI��Ɋ�"~�\N)��h�]�ۺ\����	�H`�q�L��z0��-D��+x��8^�.]�&����^��˼?���Y��f�k	�]���{g }���<�Ѥ 9�ә��zkQ6Y�%�Nj��8e^+%����j5�(��w�(:������,�������b�2�ޏr>#R�"�k2��N���x�n�$v�1����i���;L
�$3Y2]��om�&�����n��v2�������@-L�2ҙ�P'�[10<!�?��<LV��`��L��̥{���3gc�ʄ.v��X'��
�#c��]��+���:;���o����~<����B��G,�Fm���Ϗ�@Q5Ak	]�x�J^{&��	}�.V�l%7e@%�2���Y2Ȳ8Sןg�*�y��9���IĒ(��0�lS4W�{�b1�.��u�C)���M�=�t���Ʊ �� X��:�EX�)�򥲈߰X���1	]K���.׹��������0ӯ���]B
?�uמ	]� ޝk9Ĥ�y���|*�r:�C��Y���X��0t�!��R�b��4F����0<G��N�
z�Lf�V0p�G��N�G4����:p_|#<������ނ��L���S��,��N��c��ٌp������f���vN�aF���*,�NJ�9�Ķ`�*�]�@{;6���h���i���X��L�W��c'����w��sA<�ri��dS��ɉ���I��%�an�`v[���
�^�&v>{t���<)޹s�K'<>:,8���B6��_��ރ��6ʘ�u˙d�^�eؑɑ�:��:="�iw�d ɑ U_ev�)��؉�ʂd� ܫ3@s$���.��#�M/��p.{>%Ԥ�ţr�Ű�f�q,G��"-[E��z������>�Bfұ����3�M��|2`Wc��u8X�b�	d�i���5�U�*yx����Qȴ������ɘ�c)Jn��A'�Kܫ�e�Z~�h0	p�#g��m��J77����*(k����f����-�Ŭ��T6���v���Q[�$�t��f��;k�ĳ�c[� |��(��"Tɕ	E�\&P_���f�`br��pZI�)�F�I������;_:�PQ]~w����8��f�2�X�hm6��)@$�eyd`0��j�֮��C�/Eӌ6Lv�z۝p9����&
�,��kq������f!��cU��\0ځ_������[�@}��FeLL�"C��C���6�'D,̨ ǂ����Mj��]'u���/`N�l�n���⮻����x�x��W���[\��[fBo� ���A%t՝Wy�Ue9R��Ѵ@�9�M���6Eg�
>��y� �JY��h.hF�ϯ�rŢ��f�BM�H�+��;�^D��ϥ���ұsbB���\���􎯔%1��aqM�z>��G.�ݫ�s�O�N�y�t�L�j�>m����tG������CM��	���t�s�w����lL����0q *����X��IP��E�k��$t�Q�Y���Yu��W�s�K92�Z��cx,.x4��9�~ۺGP4�`�yQ&��nS�-ņ��k�B_@,����.][W�����������N��'��{�b`�̰��G.��ZQ�ܰxg�gQ�F���z��-�v�-F���L�`���h_�;FG�5�`q7ݘ	��m����������ާ?���۳E���h
�|�b��L����i���LKT�̊i����uW��7��� �e
a$�Pp�{�ٟá�*^�8�N$�X��;x���W��(U���t��� ��	��6l����q�PHu�3TU�h�����0���"�׭%2�X��"�Ȥ,���$����S0��� 7)���1��+Nj��a7+�Ʈ}��NVt�<Kg���i� ���<��8\NL�n��O�Z0ػ�D�-��|�hX�/>��r�S� D/�;"��S����edk�I@䳌�}-�ǂҗ�%J&D!����)^?�����ɵ�׊5)���˗˲Z�D�3!P� ��@}+�n+�_������� 2�������~(Ah��5�*�&�ʆR� ��#b3v;=p�U�s��G�zf4����Ҥ���VA�o��%����W�Kss#��$���t����Ҍ�_�u��a�6�� \|�0�\�GSbS�e�E}�[�ag�L|��+0wA��1<���y갽g������L��^�` ��#�	%�A��|�{��RW#o�k�E��<mټw�y�(8�q�(���!lܰ&�o���7�?SJ�8g�ڛOS1�5j���ϒ:;x�q>��Ő� C�D&_�.�K�t�'Y%��Eɚ�P@M}������n�V�*�q���r9�f��b��?�4��|i٪q�EE��>�v��<�W4b�"$�`O4Z��u�ڸ}�E�n����4��Y4MO���J���xr2l�U���
��؝���ت�����C%�@G�����5{���0���9�~�n��q�	��������N���N����uJ;�XB*�/~r���V���>��6��q Nɺ���:�T2�R|6�A
1�!9׊L�l���Ȏ�.�<_u��|��KVL�3�a֙ $a�um�Jđ�a�׊��Oe����9j���3%��H4]>�J��ۀ��~�Y�rx�N��j|�3[����p�M?���vXL4bQ
@��	�:�c��1[�7����a�-"<2>!���01����؊��q��~�ֵcl2*".�t��)�YjQ���Œg����FB���*77�������"<�fD�I�$����N���I�AD.�̄�+�$��W��2D��73p��LL�90Hǐ���������+/��o,��@?X��3g��g'���PP���`�48<9�E��u"G޼�"��HH��9�͒е���F��V2��~)�g�r��9�� ����c����Y��*�Ι�QL=��al�ԅ�@lv/�Zg��/���p
7���X��JDbY��[�޶H
���V�b3��օ��I�#zdR:�)�X��f) ��-��#C[������|K��&,F�/�'��o����V�y��r}.��$1ܢ��ՎP8&r�?ش�rF�#��1Œ�IP��f۶n�}�y�����|��ˑ����a��~X}�`r$���]�D:�KO����S� �GdO� %]G�� �Up�O��0ib�"��g/��7n�>��S�Coo7V�\�H")y,Z�(EAZ�j	��Q����q�ũ�#��8>�aN�T�㲙 pʂ8�G1K���L�x~X<2�9�t�S &t���zp*�s�����H�y�+rF;U^'�����_�I�{6B��J&	^7U�VP(Wײ��2a>�h�6�u��d_-	�Ak���?�����v�h����U<��Sœɨ�g�F !^�f}��_?�4��y4�y���Bp:XPD��j��'�z&v���Wׂlɀ��.	�@�ci�,�YPw�Y\s�Ř�Z�M．���6��I�@@�g�y�<�;{����F�x�3���ʟyF���Mܱ�6�����x}�h��*��m;഻�� �.Էw`0CJg��Y�U%�Oe�~����jK��ْcQ4�G>��M�#��t�i��e �\r;�umĬ�������O>��"�]c������@D��-�B1�����q��6̙3Wn*�䂴���+`�R��<�Y��2��i����%`���O�d��4�7���e!XLF�3)y��6���R������;=u�ƒ�U�~��jv�}1��u��UvI���Y�������Z��D@;m��jdB.���#�Q���p�'�s�;����6���O@��*���6�� Mu���"�yEO2��*H	0_%&vYL�t���U{'a����@�쬢K�3�ޛ������秷tE���f,�g�T����ϧJ�`l���zT������w���>�W�kj����:O>�"n��n8�8�Г�n�&���˟�u�	��<��Q���Lcfk*�0"�>�q�MX��-�n]�{n�~�}��xǪ~����蜍��Q<���w�/n����dp��	��I�������de�_��o`��{�A��-@h2�D"���ň�[���\�SO:Bt�׮Z���0�fv^zk%�Z;1!U�&8�g�Tx/� �b��D4&����qNi�JWj�]�I�Q�0'��]?���Aq/dAK���hnaq��zjj�Ū�~�����E>���i{Ҳ>.�����y>�;�z�ʄZ
��xt�?3��������n���,������4��έ��� ���\rD�sɠ-�f�EV>l ��&���SbF���ȃ�]6�;I����"��=���$=�����{��(|��>�,����8y�{��}\B׾�(��J����&a��6S�O��R+dR���Ch����O>t/�6~�"���LD�O(���^g��8%[=(�0X=�[�Э�УL��[�t�`#3j���Ytx��G��cK�͆�uob4�Z�<�p���l_���v<��SrV�l�"TU2:�^Y�ʦ�Hz5~o�ц����ǋ/���_�97o���PA_~�%LDbH�9���t&�����Y~*��y�ȷ���C��XK�dW^�%�uZa0�0<8���DI�_���.�Ϫ�׾�9lٴRn��~i�����0b�8���:���"��!�ݽ�^(�K�,F��N&�1���:�^'hl鄞Jk�pf��3���O��t 	��턎��LB�P4`I�T�|	�p�nL6':�h8�5�闿pG��C44H b�#}B�54!��h�JB�����6H`��TBW�4������ �t����J��8�³K1��_9�<���+���=�O?t�$KypEfJ-q���E��ªY�^���~Iq:��?4�V�Jpe�P�z�QONx�UbW��Լg���ɉ��?K��UvX���Hu����8�ē�o}�.}���g,\x^}�-|���q��
�Tğ��nl�ЇD�X�,|b�!��?�p�f�؄;n��N����7�2�ǂ{K��ēK���{���/Gs�u��ٹ��m�3Ͽ":�:�>�'�v
���yޟ��&x<�@� (�r1������H�S��݁�@�n?|3���r�x�p�4K�nvxP��Ne$q�k���5%�4��LU�#5W32�6��V�	�@�\�/�ƌ(�F^�\��y��6��R�@�0ihv-�H"����3�|��8�?Es$U�ML,t�Ҧ�e�����^���4�'�1��#q8�>|o�ا$<|a�TTB�-+��gjpdX��Y �2I�j�2u�ב�X��8y�	c�\M�suT�;z_=h����}᧧����I	]���v���s�4u����V��o�5��&52Xi�`�\.g��<\6;"�}8�E�u�p�]���ε$-��2���J����䄪�%�0;��FP��j�<���@�\���h�n����އ��|	��.d2!)�Rq��[q��J�ͳ���\~�l�2�y��ַ�%y��F@|M<Cb'�+Kޠ�#	�J�g7� �򚕫q�q'�k_�*�����4e��RE�:�F�kʎ�S�C����{}���c�x"�b�;��p~Y�Q=�^���D��FFz�u[�٣@�E!K�CDE����B��K�Q4w�8�v�}n���)76~�B�4�y�}�Ѝ:?�z��b�f&+�
��N���mF
�!�r(��b�*b�|�e�����W�_M����1w��8~s��ᩩmnr�n��-����N�~�&�tWR��˓ƢF������J�F�g�����������ߌSO=�w�xϝx����s���	�4�A��9=���Ϫ��1_�*(y�yg�n}���-yk��g�8���[g�.��&ׅ��l�UEix�<P��)7%��(�v8�1{I�09��?u�%Qu�I��_lU�wΑ)̦�[p�a�ŵ?�O<�w�q�(L�y�8���)ُh��K����C�L��,ف_�|"c�X��K��o���p]���Ux��ELb��ƲW_GSS�����6�����SO>��{�y:��F,�1'�E]Jz\z��Q.�f���9�q�ϮǓK�.�7\�C��c��xo�:\��hn�^���6�(�P���Z��̈́ĝ(�9vVj��F�*�IQ��n'Ȍ�U,�W&���~se�,�	�#ȫ"#h�81)��pF�hf-�eu�9(���^B/��H�	]NՕ��c�
A�1)m��癣l0�?��9N
� ��t]�,�!�C� ��������T��يͮ�5'F�%���vUEs��d"%
qZ����a\3���%k�0���ch�S��������ߥ-L���IB�_N'H��?��l&�R&�sO:�N�[o�Q_�����å    IDATE�!�:q�cq���FY�\��;t�6t6�V�}�]K�:j�Gq�����T�s݇+�B���h����XT��O:�$��i��d��Y�F�N:�D\u�U�����$��ڑ`@}E���;Q�>�F���}��'Qxޜ����w���M�sd�^��P1�`����R���K�>���Ȕ]��b�Id�8@lhhX:�Y�R�������>����DRr�E�Ո�����a&����k�COO�\Lp;��cg�t���AMm��#��:%_K���]f�,�bF�dneG^��:)DM�*C�DR8����q���6
��]׀��I���W�3Y��2����A_�����!�H�Z@�0��P�\%�� ��	�=ұI�r����Y���%F�Ɖ�\�,}�Q�Y����Cǜ9رa����x�Υt�Ii�j;t	�DnV5���&V�� ��r�S�H�H��IC��N����xj "-�PV��f�(7�x���̙|_��0�� 
;��wl�{;k�,�D�Zq�q'�؟�txl�:�Ưn�߿�N���[�ij�gO<�}$�|�ؾ}۷�����s�+؂[n�)�c�X�拸��kp�g"�̡�{n��6������hl��nrȡ����d��V~��x��������[�\�����眍�}�͸�����.Ǜo-����G�;�y�I�Q���W��3�B��_z~z��ڶ ���hj��\و`���Bd�:T����.�g�tz�YM���2�2I U����7o�LC��g7NWA@�)E0����.�v�����KWY�ڜ���	���J����T��qI�
q�	�3�۳d����� ߙP4)٪��I���+@*?4l�[�9���"��k��)�L������\S&�J���.����9&�u��j7��)-��Zaz�eA]�%�g�矴�>��Ȥ�	�5�f�&d�S���d���&e�(@GfRظ"1�QIGpȢN��Y<p׭h�� S2���U���w���ъ|ńB�,�2:��r�b���gP*��K�J�a����~��31t�^�'�������Q�+
�N����׿�U��"��k�����=��*ϭ�=�7��dI�a:�tL!	�JH����4�1��:SC	���{�Er�eu�����~�Y6��{�����22�F������ܬ��A9?���nXmfQ�;x'�)���L�s�?O�}w/;�p\��+�#��c��h���ndu�B�����ʪ����/|�����`CӬh�6�7��N���[Z��0�$#�r�8lVβ�0h�7��8i8Ty���*��PT�U4xY��l��b�$x�])�ȤR�l^|��bX-2�C$��	ǉ&D!��0����<��iQ-*�A<���i��ĨZޢq���1�f ��z
�?�4|�٧bjKѽ�r�Zx�%rp�M��*��,@#U'[к��G�(��ο�Cw>�A�z�a�\�ol\�3g>��M�E}�#'C��c���ٰ%�E�_��p�2v�sԄ��PI ��a\�;VG�B*�(�1��$;G$z&�S�A��Q�k����>��H
�.g�	�I��T ����|�y�b����#���UOo ��n��>TՍ�U�܌��,^��n3`w�G:���`E:�ِB �3��7�@�͸隫0f�H��t�>����PR\�X<��Fc��8���p�W �˘�a�f����'�X�d9�:�(�����ɐ��<�?:/����s漈{�K�.����;�xS����F���g���PO>�2L�"�c(��F$�����T-o��$S����U�G��T`�Rt�T�8<⸖H(,���UZ��\j�o�XQ�h8�I
����Ĥ����?�3%M)@*��?K��"��|(@1u� �d5Ģ%� �q�7���MƌX'}�r��:�;�������ۥ�'���ӫ�֤�b�K�#�!�N��Wl�D+�7E�Ϸ�I9��|��L��=��B�	O������^Þ��i�zN����)�����.3�,2!?�N9� h����F��(�T��0��|'��bUc�#�?Z`� �C�%t:��I�arXм{���ʝ&t�؂'��Dz^���RQu
x�Z�a'��g�}&+Z^sq�:��riy��P ,l�M�7c@m��L�fN8�L�|��˵غ}'�5H?`6#�!ʽH:���Ȅ���˧,\�sV4��$�K&��G�[�@p�Ʉn�$�� ��r� ,�$&�����I�VXD"#��N��@�Q��0~�D��;vl��'OS�ݭ��x�Rh�&,Y�����"?����iA ��Y��!���I q�^�Xmz�N�������E,ɽ�ټY���R�,VDc	t��ňc��(��D$�$s�G��L.�<_V�)r@h�>z�F�+	=�l<������0a�`�|ݕ����0��)ؾmF��d<��[�e�a�����Ұ�ҕ�P�����pT��v��n�T�'L�](H���S��(�*�[D���2Q�*�tE������8����޳|o���XNA޿��k"�J	�5��b��7n�����[,_�o��)�}�m|��q �}a$���	��Z�_���1�{�q�"4n\�{�vJ�lذ�}� d+*���b̸Iظi�$�믿�"�vm������+�fC ��Q;����+4�4��v z�A�9J$���[q�C���O�Ηs�7jİ(�U"^y�{����P7�[��z�J��r
�@-�
UN	����~�(:����ʪ>FӒ���И����$�c�]9')"\�kC���ɹ(�[?>u���w��g����gO\�:�VJ&�"e�����O�!� �$����Y�}���Ʌ�l�B���F��� �)�, N�С̰`�!=K�C��T��eW̃$���F��F�IYW�]�HS\��"��=�p� �c�ZeU�`�ҡ���ۥ�-����,g$B?Sw�{k��	]���EH�S�г)D:Z�v��C�S�O�{�TX��X2��N���S�`$�`,#�����݋�ь����
�	dS9���,�Qd�1L��F<f(�{�yԯ]���7"�M��t�ue�PE���y}D�`��3��BU�Aq,�|�6�Q�=�J�΀Au��e����o�s�����L�,������p���5͌���$�ɔ��Ѡ���B�N:�ΐF>A"�M���1�0��=��| b�w�X�t��F���
�����.��d�"\z��X�a�p�?��+lݲKoB(�μ����Ѹ�\Æ���.��j�Q���fZ���N4���M�(xCs@k�Ac���I"����BiY�K+�����,:��@���f���X<��ZI�
��G�88x��=x���X���ؼv�P�����gQI����oi@<AuU��*��I�R�
Wv��9S�C�߰+�T��σ���	;��TA>V����A6��>���S�D&��g��>3�Q� ����C+݋���g)�_%�����`�֭xg�;�N��m��`���F���8d�t�	���{�1� �4"A�2�#���a��`3���Ҁ'gߏ��6`�%x扙H'���ӏ�g/Z�cF�CՀAp��������w߽���[�w���*7mڄ!����m���p��w���b�ɧ�S��~���[���X�v�M{��N���?;�p��pv�j�Z%q���+��}����R�)Œ��E
��}.e\�0���a��
���n�H��c��Qr���;�3�@��V@�����Jc}��_W�?a�p���	��)eG��5����γF�Z�2#igј$B�dQp���Z]Gլp�9%�c=��_�{<
O]��o�p�$5Aw
罐5��j<�� <j�¸�|��'��5����fB'�`ߏ�
��I�"��	�  z�;�Wex-�q�'#0�C@��U��̎�^y*��F�p�%1�\2�ēYDi?ju+6Б�/r:�$t���r)�<U(�R ��C}~|�]�-�������r�
dJ,�)c�8^7�d��8�N��
�f�޺Iku)�~2FS�4��%JF�{�"m��B7)�zL��������x�1�7�bB���b<����NLVP9�T~"W:�&	��4����;���rn��fQ�b�ew9q����7�X����f >��C�����S���ckK;&;��v~��+a�zE�4a̸��񆫠פ�f�2�o�"T���f,Z���9�gg@���n?���њUk��+Ge�@I�&x�Q�t�X\�\�*�*#&P���r)LC�c��:j��{��p�o~���<��G6���,476`�����DK�nt�u���L�3���F��
PJ�q_Ȁ�
���v��xJ9ǝ9�4y�#�5�	����,��LJ�ħ�(�6�[��@��5+Jcґp��D:3v�*mF��s2����˦��|��uX�~�HA^q�X�t���q�'aws>���ڰ	Ͽ�6n��ؼ���΢DS�7GE�\��ä�v�c��м}#�-��?|?�7c���X��{0N�p�Labɼ�ԙ4zx�����X�r��v	����/�&1�ǎ��Ukp܉��+����f��&M㪿\�����j&�1�X���VD8=%���c�,��V�����l"	���f���u%����"{t� ��FS���E����>�N� ���d�� G�ڔr�جFʪ�ؾF�}{�����6��بY�=
>��x� ��uJFвS#�[r�)-�:�;�OvT�P��XD�.�K�{�y�y����	'�v	���p�`A8�O-j�J�@OJ~����f�)S_2�=YV�+�:�wM��?ա﷽.�ׄ��ޝ������Q�iM!׵С~��
�B��8��I��ɤ�=m:ԋdO��0g�|��Mx��`�����b�XG�2���Hg�6Bq&w-lE��FU%��D��[\!�8��
�9�6ƜG��Ȧ��ߋ��fp-ǂ�Όja&�e���<?��$�k.�i�����E9��˄��B,ϸ1����Ԋ,U0�:����{�l����ew��>Xv�����������#a��.UZ[K�t����O�r��� ��9lvo_����g��DXA���ګbi:u�T{�qr`8Vf�6s�L�<�$�W��9ϋ]( �ގ�˷��O�d)C"����8q�!0s��% k�zP�裎�W����{�$ �Z&"��I�^F��Hv�%�e��5�l(0�>=gsZt��.h�302�$�CJ�t���8k���	�aw��F)�q�՗��q�q˵W��{n���r4�܆C9+W-���9|b�%�B��M.$ ��dʝ:�us/��ݬ҉3X��4�	L�7��;\�[c0��O�2��@��yc��( ݥWǉ�v� 2F����\�8po[P��V�!�� LF_͟�-[����캤��8����9sp����/�����ӹP\Q-V��|J��<�v�Q����(V/�M�kp�5Wb���Jw�K �jf��n����0d�0�x�����ь���r]�Hc��Ո��8�Wg��S�._7�����ow��/>�G���{�K��.���0Z�r���|A3="�q�sHSc��O(�j�A�UUם�qJ�j��塑��N���*؝N��pz�k�6�<e������uW�n�U�ɠ��E�k��]Y�y!�+I��8$CqN`�"e�&���>��?�EwA�+B.�'jW�T��� �,:e�K�Get�c &C$�S�+#v�\)�c)���>Y�R���g�W��` ���c�^�o�Ix쉸���M0�w:]��K���X��טۅ��Z� �j�V�S�?r���cO�W~�b�oBW���!��y�HB�_@��3N��'t+� �\��C��q����F��m�Y��M�d�D�E����A�����}:��VO)2Z �9JBϤr�(z^�E:�ˠ�.D6���;o�ı#q߽���ݎ�˗���V���~�1����x�T�'Ϻ��ld8����;�\#'��"�[��7E(����N���ɣ7Qx��_��}�G+�_���H�6�R8~q��0���ީ�4D�&��S+;�\�NCc������gp�K�Wv,��}W\�HCغu3Ǝ�%KK��z��(�����T���nx��X�h5�vwCk�����v�S�������x�6�Æp���O>�c�>*�h���!�	����/�]˫ �Bg��j/�&Z*~��(�@P��Q_5�JF���d �X�E��t��A"�A�d�(/=7s:���[X�x�x�A4l݈�&(T�U+���;L|,�b����@ C��$Pq�.t蹬�$� 92�z�����{E��T���#���U�Y��E%�[�׍�E>�χ���n�R�HԸWǯన1ed�uK^}�5����~'@�ꚁ�;������«��ˮB��8PT<@l��s&R⌗M��QZ��]wߊ��[���1}�]p�m������+G�,tv4����߃���7� T'�NQ���U��)AiE�-[.���<�w��|ƌ�0���q͵wbs�N��Λ�ӕw`S�nQ	.��W
�A�NX�[Z�Wv��K�����9��{�u�V%�r�NN�Ɉ!Æ�Ǣ� 8&5-�ד�� ��+���|D�&(�+ᇝ���-��v檊��ű�Q���[�A'�nZ���*�p=5�+>����)����X
�V�+�z��|G8��K9{te�dq�$� (}�LD��R�G4m�iNu�ʎ��	L����y�{��fE���Rjx�a�`6��r�[Z��n�L��J�'Kb�ZE3��&[����J�ƕS�^�{�[Sz"�Ȩ����v��������Z������5I(\u�>�Ϗ	��c6/�2-ҡn�|m8������W��օޮF�m&I�,�ISf����セ�3�|/��."i��5 ���F�]�����VH\�5!x:�mԢa�BL1�|�m(7��_w�MP�j�V�1��������Iy�$?��F�Y ���H&�����iws�<4V�y=Ry-�k!�7@o��ry�|����v=�X�vG��RT�\V',�Z;� �	�AMZ��Tv}�'��\�H7�K��<w������x�U��⋅�T[S���&<��s���SN�v4�BEU�.Z�h0�[��a��uV�T�JB��^S��.��-;PTd����G*Ƕmې�E�j�H������1 ��{�@$r�/�P�)�0�K��f��%`򦯮��/"�we`#����2"ء�)NC^c>�r������w4lZ�;o�Aϸ����ö�-b,"d7ٻ��I�߯$��1�nTzb����8&W�%�l+�����g �3P�-��JB�&���`U�5��:�C��	_7����^N�f�x���[�yoSя�e�5��?�+����ز�^��u��EK��s/a�1'��#�ß�|�hh�V�E��'��Yt�H$ø������O���\��"�8�Q��,d�;&����:j�B� �#v� �A:���_t)�9�(̞='M=Y�ml�ŗ^��/�S�9	��64����(�q�x,S'�U�^1�����_��_���V��:�D^�Y�`�y��1h�`B���2y�Do��Ɉ>��1%E Խ?���фN>�R쥸�`w���N+4�$�fE`��(t���q�׋5.��P�����!�J�ȈdA�
��U<���;6�)p[�Hc��G�<�W#��0��8�F&<u�M&v�{�h���b���X��/
g�=J+��ETQ�ť%�~7�5�׹
b7��O̐� R�"�L��$q�ŒS�=ԉQ(<����c��I{�d��1}�+�QJ�Wy�������.�Jȳ�    IDATC�	�%�ǚw��#&��'���o>ƦˡqG	�F��[h�RD��U���շރ�U
�ŋ��,��jCO JCI�K++��ݝ��)C��VM
<�7�<q,��o�+�Α3����ןqFŒ�Q��P��֙�>V�'���%��9�~�TP��,�h�?�d^� A�;��<,�r�����_�RܴW��t���bi�5�˘�t1��	��}<���X28�ȱ0�c����ePWmm-��r4�O�>�{�1�88㎘ 9@ƿ �X�e�9f,�����Ԃo���77�qW'*�F��v�;;���ø�Cp����a��C��ۃ�O�Bg[+�|����Î7�L����J1��W����Ѵ��)���a0Z�3��F�c�Y��]X�Kb�rX3�jw^h���Y-t�JF<t�-x������W^��'���7��� ����J"TsNI�;IB�*�V���ⷮ&t��9Q�\��E���y�LŮ�� ;t��(EC���-����^��ڹ�`��]ho[Pv�|���lll��| ����o����<z��ٰO>=�����GMŭ�O��<����*�i�:�H�c��h���cqۭ���I���edOk��A5.��rټ����NY[P��m��\��P/ZZ����f3���P_�Æ��%K�h�"l�фÏ<���_���ذ�:��(��]��5Ԭ�b���!-��Ի8�8�HIh[q�Wc��r�X����]�z�����������E��G�w$IU���a��1�%�(Ԭ}��Q�2i)<G���$I)HI_d�"?<��붉v�� �sϠ��a�k���d,O�\����쐙���[R���n�uz���������+��g�Ihy<ϫr��r���<'MfE�FG����	-%�SI��:������1��q=_#�����ԙ�Y��4I��J<�P�>���)j�|��:G,:]���ٵ�Y���O���{��Q�\���w�?����(��Մ��C���0��CO{ݽ��$���k������n��:e%��>k��2���f�VD�@8���^����+L��0�Y��W. �s���N3B�fL9p,����_~�-���`�B���R����U靼�*�F�y
�"'8��(ar}��#9�ģXL4�Ӟ��B{ 
��D0 FW2;�V�ĩ_�9����hm�X�2�7�D:���.�Ig��.�FM�\y-+�,2Q,��/�Ô�I��)'#�}���0�?�<���z,X�@r �Y#F������a���h��Ɉ���-�b��u�Dr0��Ej�⥼�%vF�^&�-��p�����-ͻ��*K$K%P����֮ЃH�!��dA&OW�*+�7�a�����[k2 f'k��\E�2�3P��U_٫�Rst��B���&��Y���gA��W��B��ލSO>�7mBkk\D�s"�K@�t,Žya��(\�4v�J�Pw�LȬne����Y�r��v9���J�(�D0��]�l��yy�7�8�q�nTl��Z����\'�U����-+&�[n���o���A]�4����Y�`��	5�`�q�C���`�z`�;do,�I���� ���ѣ�	��j2����|Vƹ��S�%Jmp�;kPSS#_���� �I9����|��g��_�Đ��p�7��O@}�6lܲ���\v�������nO��ƙ�5�*atV�F�w�ݑ�p6t�p�ᗕ{1��?�ן�˥���s��~Z�Z�����&�Q&t���e1x�pIJ�v톕4MNl�Bu������!����`��� ��߉����qh�����"�V����W�-��� $R�V#ht
��V���dS�iQ3b�$wZ�
��Fm� w�:��$�ΟI���g�g@F�y�Z[e�n1`�k��X���X!�'�5}ԹF���ѢC<�+�1��)���؈\V+�Oy����r�дHQ��@�����H�{v�ʵT������&a��RU��^�!�F�*��@��h�`bm�0y�0<�Ƚ���),���6)X��9��nz��p�`Ԅ�«o`����S0�K�Ә�י$�����:�U�����i3��8�7'��a�H���Y���	�¢Q֋�j��T4�ׄ�}Q�w��is-�ű
z��ڱCO'��h����� ���VT_ ��X�}�/2�O�x�IK�4>�uLO8!	��OL褅1�sƄ��F�q��6�����fH ���Icq����͸h�b�SvȡX�x1"���l& �O��o�eW\�p$w��|�1�._���Vt��P\9�x=��$�J�[�K&����->|;� �3	�\�Ṯy`�I$92���ppLW5�Z	�z��#h��.C"I'&r����jZǛ��21�ݢ؃lyp)��F��	r=5����x��ixm�l4n[�k��=��;z���� ��IX8�"�T�T[%8	��aW�����d��U+�*OS�q����[�p�wv@�=�ɍ�P�R.t����t��z�`�����S��e|�!9Y��Ca�$1�����QYQ�K�x6�߈��P=P�|�q<�(p�\w�m0ۊMdž�����(�(�M��%)'�B��Q�$���bTA�GZ4"�*@'�N��z�]m�HǓp��^�{ 2������b��w�ŗ�������|���'��$�}�V{�b�c�f�Z���
�Y����J-)���].�|x�l��ˉ��!M�/��Sl2[Q7h�L�x�(y��F"�Rd�� 0S���P�?���"P:tz2��N�R	�Y�2vl�p褱��3���-�����TL �.�mmزi�$rJt�5J �ė�uFl���Å�-�{o�:�Hgm�ѶP�
#v���ΤΠNP�ҭ)�B���;/��#�2FlE��P��I8�MM�"D#J�1�d��4d���	��q�ѓ1f�X���[4lۉX<�H,�T<OY�$�X2+�9�V��x!��*���Cײ;���룖h�ʋ��?��߷kW�q�J<���xBO�z����ɓ0r`9��6L9�@d�q�74�{�xd�P"F?,Y��]�h��AG ���aH��4���W^oY�b%O
W_v~��3�I���x&�C�#��P�C�I&��T�����{��s4�H4&��X,���SC�Ho�"�%3Hk",�.� n�dGJg��V�U�{��'/Z�4#�(v�참��й��1�g"()��y�f{v�eI��c&��k@8Ё|.��ÇJ� ���`.��Z�`PeeL�:��4*���V�Ub�w���BF�F��DiѐQ�~ăa؍f������T��:}V��T���+�:���*�	�w��£�$&r��R�;�#|�`��z#��%Ei�:�ac��i
��j�*�2$���׈�6�&t�N�x������~�r\��K����F��n0�Nt0�`�ٿڌ ��n\�hA;[n��F垫8��Ϗ���V�0�"��?�V�j� *^`���U:��@H��7�'�p��ظy^}�uz�d	��wPv����v�YO��3�ĤC'�ڛ���@6���`yZ&uV�����!ЍZ�M�)�2ɨt�}�v;B��x �V�f@���Ɍ>��%�=.��vA����{n�i���?�g�����b\p�ɸ�o/����U�X����ܑW>K��* ���$R� 6oX�K/�4NT��/ۀ?���fy����:�tv�h����R
�H4.�n�9X(�p�����,�롗iGf,B�$��0b];q��!x��G�d�
,\��hD�Y�fąa�喫�~�N,Z��sV�Z%Zt�����W^Ǆ��]�W�|�7�c�ైg�P<���k,�#�.W���Ƚ*t����v���RVA�)0����H@�2h�s�1�q�'����>�4�QҞ �N�[y^�4	�@T{��C7����c������ �TN����42,)p$�{����^���3e�a��?q���2��xR1��a.4
}�z"�]̏#��5e�p����q��cԨRPJ�6�k�.�Z�F*E�X�j-|�8�kG�*+�Ήt8L�^�JK���(C����=c:�����7�����v�TV�*���$�,�x�2^���:�8|n�w%����I>��F#`�/.� ���."ݡ�%��{˱�݇��
���U(��H���<uن]��	��ѩ�2r7j��l���нEN�ضV8�L�-�-#T�^'Lf��s18�z�h�`0*����%�
�G4�}]�s�jk���aX�`=�5t �q��$ձ@C�d�.����F�3�D3�F��Ǟ��`1j�q�Eӽ��]�}��
c􄃑�1����28�eҡk�6��9y��$���cB�q�e�J�UA��bP���5)\�OEp��#�o�?�}W\z>r�*����f�R)�g�׋"�	�iY!S�S�)�r�.Q��y*ձrW$3��P�hU`��Y���n^�~��>����	�!GJ���rVw��#ϑ���%�C��B��$���f���v����A2��ĉ��rz�����Ͽ�_n�Q&0�<�w��eH�(�i���h~&tZ�R��;�%e�U��� |�-HD���{� ��OP�ܣ�Q]3@D��4���G,��nD{Gj��λn���Dö�mt��Q7x�>�O���f���}�I\�)=
,��B	+\vnv��D{�r9`!�7����8�tԄ.>7���RIFT4��Ģ�fA��?�7���^��C4��ФB��]���T���K��d�"|����p���ƬY3q��g��c�ŷ��/7N޺{|���K��y�`[c#�:�<v*���o݉�a���Bc�!�� ��ʵ!b�	���p*H=>;��S��"�9������H�H*��w��q�����-<����������E��~F2a�]8�ȃp�=����zrx��w�y�v�jnG*������ti�8�An}���9s���8{q��w����D���W��~�ǽJ�I�2��CȏX�Nq؁8�7�cݪ�X�l::[���Q^Y.�Y�|5z6�J4���=��[1�n8�M!� �p(*��[V*E*)k���<�jJ����7��?��:���&.y�HL��(�J�'�lo���~�:�Pv*,�����M�"R�酑L�s =�Ju�g5�;�୬E{w �W���2y�E����`ůohz0����G4m:�wB7tBia�N��ݻ6aܨZ\u�YX��h5!�G2��f0�e,GjGj��$p���[@=αpLP��5UrAJ=^��yl[�������	)��Jf��P]Z�ݎ��&�l&0e�[>�^_v#�I�x m6�p( �ଳ�����FiU:z#ذ��6�#���܁��tF��fHp���f��U�fTY�<�a!MɌ<5�ca9̿:i
���,���sq�y�C�ˊD(�C< �G"�"��&5ڕG����U�lJ��V �P�	]��V�r��+^���_W�y���Q�����.�B5jp������]A��g��՝&w�,I�g)L�DK[;>��c�"������}���rL=�d�r�3�Clkl�#3���<������nhw+	K��iZ�j��;�"D��TrX˼�>�6EN�h�s�$˂�tD�8�Wz�x,��و�?&�����Հ`����u�]�&���#؏�'�
���_w>$4�H��I2b�F.6;q�t���5���(ҙ��h�{�e��NC	��%T�`8,��G�=�ф�Æ"�J���遙��D
<j)���5�k'����	lcI�.�"��`���V�t�e�f�a�������ĸ��� o�� �Y��;z4V�Z)�~h���C0;<��'_�+6Ao� �Ѣ;QA��4\���":ä�j�S1���&�Ϟ��2ʮ�n5"���a���f�i��~��Z��λ�h�D<�������钦��4������Qc����s�n�^�Y�t����|,��K�T��Y�a��j����w������:�H�2)*`�C�U)k裿D�EQl3��c�B<ԋl��W	�W���1���)|;;z�ze4zđ���kQ2h��f���u"��xUT^*k9�v6��g�D�ׁ�x/>���ރ��WT	���
�g��ׯ__��Pd��M���lv***p��������N��U+��lش;����ц�:�n������_ �����fن�RZ�0&tv��ݤ5���C@&��"�k߁��Ÿ�oWc�ү���C�bq��=�^�F���r���d�9N��"��d5)\f[��a���j�zS;�:#��STR�!U�D�R�3�&�Q�f���F������Q+f-�`���8��0��#PVY��]��n�R|���0�9Ho�Fo�?���n�l�	(���M!�:��q5�}nss�{Y���@IH���k�A�ⱇ��7݈	�cܰAh߽�U��uX�p�p��ʧ2��_�$L���C����93 ʾ>�X�2!���jU-��Ѩ������~�y�e<ꯓ�T���	��￻ﻹ
�2I($p�ϛC�����¾_� ��O�t�X�l5֬[������G�������7�vn��n$r�y���D��SR.��'
/�h�ՀǏ��܂��.�	�T�`@8�tl
�"�Q6b8=>��C�^�	�m!I:��S������������?>�e�h���Ǟ®�nt�b�q��&@+'k���=�l���GI�"Kj�[���Nc�ŢLDv�M�J����Q��bE��A����c!ɏ��jYap��<���F�?�@��e���s�F���x�6"��p�7�����w��� l*�E�Iѹ��G�C[s�.�^ $W�:d��k�,�����;�{q�}�U����Y�]��Jr�9E�IF� "���R$?������
�=�XH�e��H��f;���8��3e�ܳϣ��]X4�-p�p��g�(&���y�eY���4��G��< x�ifRX���I:�}��}�~��}��������������QK���Pb��;��:�v�H��(��`��`�^�?=~�`.w�j
 ��F�6��p�at�z�a�K�deQTQ*kHz�s)�q�_p���x���ㅧf��؎x4"+#R��9�|���e?��x��'%�ӗ�v���8�U#kde�7x�0�wuJ2i�D�s�����o���~�%˖����&g)\�h�G��J[�E��$�oly(�q�G�'���6��]ԄnГ���ӢGs��{���+�l�g0����ys���c5���Z�f%��/�W
D��vqQ㎌��j>���o��דƺ��(<�ÅN��&�`q����$BQ?LV3�{����a��a#�ECa�����n�$�d:��"	"��z�`A��rZtt�*A,W|�i�J�q{���'�����p�������!�����c��n�ڨ��~ϭ����"�݋M��b�С�<���"���j��J9Ʀ`	�p���e@��-�}�J�7�
6��׬���ʸ^�jq��b�v?�)5�(	^ղK��#t�(��A�H��t>�~�bq�q�ۺe�ص<Tv[7�c��Ex�������=>��X@I�9�]9�*�A"^�p�fuR0d5)x�vX:���Sq��Ѩ�*Î��x����,q�>���]><���0� ̘1���]x長ŵ�q�L�~��7���f��}#���[�t��V����XNW�n/�:x%�z��X�aZ�v��+/B$��e+�sG3�i�(f3z��@�ہt&&R�,��z��ɗg�����G>������{�o��oB��@��ky)va#=4\YŃ�������O�⯿��a��������ł8����so1Ye� ������j\B(Ek{'j���BQ� <���08K`�)�4�3#�W�݂ �y�2��P/S�Q(`N�V%�-�B 0g�    IDAT��a��E{,#��Į8��j��m2n��������V@�v�	c�W�(�3YI�b�Fʝۉ���U1aE���Zj��{n�o��3��}?k��#_W�Ol\��+���L���81P*�E�f>�ڞh
�Py��S��Z�w6���4�� �Vɔ)(�˅[w�lu N�D� ��5����Ә����+@�lF:t��Q-�Ӂg�����ُ�����jV�y�:|(+���g��y���SN���^��?�\:m��O�6M
9����2i6�g�<EE()����]t��J�1z�,\�3����Z�E�5b0�s��И�<���[�%��g�NI�	�~cpzgK��{Մ��mw��c�}7b��O��ѷ�SƎ�	l4���cƌ��G-co�C�edr�\�l��?R�(����a��m����գv�$1�xK���QCjB�V
�H<*���h�D�XT�2`d�@_j��R��z8�^�Ef� �(M:l�A������Vd#�)����ل���=N<�h�X�s?��~I���h����ju�p`�C7㭗_BG�6s�a�noÒ�qȁ�e������X^O�ص{�54h2ʈOF�yH@W�ߪ�u��οM'��"@\�
X ��
rcnV����j#`b����ݺ���(���;��쐝fC�vl�ߊ���7�z�u�z~�9().D)��YX�q#����'L{���l�z�8~�dd��������>���*R�i� Ă��4��3��Ǣ�؍���ûo��^_��$������[\|�W��	����9Ee%���7Ћs/8�_p6:|�8��tte�j�z�	���3Y���9Y	0�gSw}��Z|��<\v�E8��c��c���xa�+�E4H'��50����;lH%Èƣ}	�d�HBW;�K�R�l��L#�=~�TBW
�~#z���5y�aT8L��Sp�I��d��8�7������%�PRQ!v�ޒb�o�*����H���/Z�r%G�^b���y�`踃���o!�7��*��]�Xր\a"$ӞB"���ߩrFpg�:�v��6��P( "ƽ��ې��
�bj�sЋ�rf��I�ȯ��q�Ap¤S��lWU_��t���+���AyA��_�"_��:;�~���T	���g:(rzQP?�QU7P�=+'D��)z���T�4Zй�U��N@,D}�zx���l�)W��
-�<t4�{z����&�f��Ӏ!��d�˼��h��A���=<C�<�3�|���()sJCG0c�ĉe�z��cҤI��`�LߏGyD���<w���?�n�$v��L�p ����^-���SN��9/��YO=����o9��Q�a����ew�{w�K77O��\C�$b��JB��{s�p�M:v�)�L�ikDu��^��oX�l��`'�����
b���*��0G&
������v�:�h�)#`�|��r;vm�ļoV c(��[#c�@0�2��f�I=S�?͑`Lv2�ψ8�&/���#rWHTV�r�����p��EP�v��M���,.-��ȫ�#Ԡ���#�`��f�	���h��_���+��V���'�1�@K��n�+&����rF������u����T��N~n���@K{�$�`8(����|�Z-�6�x�¨����ݶt c��L �����y-\���h�;k��U:��͉u$o�	���,�x�t�:P�uv���ӊ믿k֮Ǭ�ϊ_4���a#p�!�����׋��*���=^���p˞���#����Z��;1��S`�������:�����wBg3⌓O�'}>��V���>�ɨ���+������v�_���� ���JȮ��$��z\wݵ��HeS(-/�1�??��$�uC���$	�H��3^<A�� �v�-8rJ�;҂ԝ������)vc8N��
4�K�[�	���TYE��"����]&Y�@�����z*�H�'����W\p.<�(lY�F��5W_�q�ăBKk;l'���[�,��야���7�[rB2܁�QT�Ł�U��f�X����h������������+R�����~G���؅�fA��������,Ȱx'ؓ�)=�u�P@)x*�z�r)I��3���Y����&�	tB�bҦ1���dM+�3���W�)���?*{�����������������?	`�w�u�P�0����uuf>�3p�ic׮�v�m(r�"��z*��U��3����l�T�V<(���ҡgDT&������>F��%x�����X�EHKd��F�������i�L��ܹs�1o�kE���.r��*vtt��L,
uQb�����F+`r�Y\%z�h��]���t�La�;�Y��%���g�!�XJz�<t�C��Y�P��M�ǎͫ1rp^|�A8��ޱ��6{
��d���X���ܘ<N�$��IZ�TF�|-�{v�z�	`ۖf�q���a�T�[;X:�ʮ�"b� r��k�����C:���p����q�r����XJ
�Ȩ��6
�S ��4�n8I`��c���Bg.��T� B�(�~�Wj�Y�?���i�!'0L�R��P;�v-^x�Q�v��uW^�I�GጓNB,�GÖͲ���;�ѣF���#�-Hyx�����-�z������j��]�iT��f�x�	��u0 �.v2�fr�d�F6��	B�\����M�c����''|o�\��!�h�Q6l8\n7|�a|�`<E�6b��av�,_���3f?-��w݇h2���P��nԌ�Au�X�f�<�H�|rlV����[�a�z)��r�(�Q?\:����΁���=]��/O[C
�ͻ[�ZS\"��N�:��=��"��mTO�֨�p��PY'ԝd:'q�8�x��k$Q������N���o���>���[d�:Ģ3j��푎�-/���0����lÉ�`B��	HBW;��<�����F�lf��]Sy��iB*��Y�N�s��]���^���p����z�E���i�\�K ]Iv��B'E�ta��=(������8j"��d��BA5��������'q� (
�����u�Si�S�ns�?Ϭ�j���3˂�?#��e�R�i(`P���z�ڥ�
�A:x�hPFԒEҘ��IH�.}.��P�)����ρ�~.�N*��@i ��w>�մd��;syTe^;�W��NkA�����1�Y�>�"/*�{�}�/�9ݾB���"��KN'@s_���t�\a �\��R)�LF-��<u�=�tY�����ހ�e)g��:!������=A5w�6���.�%�s�xQD
��� L��B�+S��`���kVoGIu��4�	�a������zk�YK65=�3z��?6�7�ү?��١;��|MR]��o�*���>�r1�����lA*�׫D*���jt���r@�t`4�G�w׈?8w��D�H�Vo�cO��0l0U!g!�ǁQ��(r�**��_n��v"q؜n�"L'�����N��B%�M�G*���b��Ha�,i��i���8��6��[
���.���+��!+ً�#��nH�v����E<�����[�K������g��".���S�>��"F��&�D��7a�����VVY�)S&��^919�9ѥ��|-*��H- rB'�)_��B��/Jo��I�}w�jܡ3��߫�����G ��������_|�~�9�6��]]n��SG���o���V��_��G��z�.���:#���<(l{{+��N�������`�}����|u��2ͥPS�E�U�`O��|�ۚd���	G�m�~���GU� ��.��.4���ls�M�5��h,*�P4$�?��`@e� �F�#s��N|�:�F���0[��;��)��*�qC#���%r��!��B����?(B�^�.�O�.b6�Օ�����[M��2)Q����H�qǵ���3�����1���G��d*�`,"*�=��	�K�Q��OJ�}�x)��pH��ɞ�uZ��Gp�	����^EW$���) %��M�#��C ��ΫQ��--t6�N-��8�r�,�ʫ�w��?���[Di�{g�V
Te�t�ܗ+nr��[!G�2��I�|�^EjYgP��{�S��♾�c���u�?��?�����(�Ay]R���|��/�{�`��G��]�I-��=n�u�w��p��������a�WQ[3;v5#@�w��dY�^���Ly��TPx�Y�B-/	=�ՎN9	7^�������@G�%gTmTX:j�V��
��ج��� _U�����Z�P�rga)V��\.��H|�PH��X��8rא��.Rx�	���j�J�?��7����wݟ7�%�t"�ͮ(�5w��:z>D��	#���i���� �oC�ۂp�\[�tp���ޅ�N_�Iw�Gq�T_4�ol�%#.1Ie�˛�t�:��ѿ�лa+�E�dAŀ�Z[Q�����>��n�����DY�AL8�%���j%)��yɞ�m�N�9��F�+3�8u57�Ѝ��$����B(FgW�輓;o5t�H<,\a�ǋ�Z���EmNg0����-�P��Ø�b@����W������g�n�`Pm�$�"�C|�)J�	�f[�P��12��n�d��F�Z@(g	����C@e4��+�c�G�F~�_�1�8���M$�ͭ�q�:fW�X����gwğ��A��k��܇��u'���6 ����]o��.-^���_�ǯ��&�jiG	��f"	��Z�&�wn�y瞃�n�	������?��V�4�����s~�+L9d<F��w����" H1ra�ʕ�������o��b ��bx��lu�2��S���nx+i.�c�ַ�aEO��"/F���;���k�Fqi5�&'"ty������Bt�#��0	R�
�bb*���1X�s5���T��%	���J��Ց�ޡ�h���8�'
�t9AQ)�u)\�ۓ����O���>x��6;�J�,'!U��(�錦��I�Z,"�G��������p�QS1��7�O��ʃ��ۊ�3ZdW��Q�[DOI�����e"��!Q$�Г��$ Ws��K���V�>������g1ϯn]&�4�\u�^H�L�}Fe��獮��S.�p�%��m�_�,����(����G�t��T�|_Ǯ���%x����kt�N�j�!��*�]��aqke���ނ�;w������f���.�k*�1h��p��%��1�)t�)�*K��$7�݅b-p����&�٧ÿ|%�
�!���d���)1E�R]$��Mx?��R�P��p1v{�����pDi��6r2,,�'a)*E�l��NY�_����o/<{�����xZ�s�AtA""�~���k��f=���ǐ�"<��=hmX��k� �0�7�����,M�jѵs޻v��]�����	A�=�G�� ��^AQ�G%�G��5!�dA�(a����g�s�w����v�z�_����WSU�����}�z֚�����J��Z���`��,���L�:�b�����t*�G�x������U�G&���^l���IOx~�?������[>�/��Mԛ=�US9���ƺw� ;e���oܸ4�pΜ���.�C�.7�ڪ5�nl�tezz�T
�J�jI��j�ҁ@vtԒ�y�O�`k{�`KcAh�Q/o��y��/þq�m�8}�AT
�8z����HM�ZT�Q���T���#=�4tB�w���F��M�B�T<W	�3�##9�f�T�"�}��AT+�K�<ɗ�z=Ӧ�Qv���rc�L~0G�b�-�v����Y���U�v��eM��|�_�G��Gq��o���/��~��pumM��fr#�7;���2�\D��CP���c���̹KB����<��F�~�9O�3�x;��]���_�4��/�7�8&l����+��?|��/�7���x,V�;����G�ތR��f/���Y��x�t�d�Nm�ﰌ	cjnVY���&"�
k%����=RE�Qs �J�5p��O4��`rf�H����x��c1�?p [~lm{[NE%�hd0�Vm6�$�eQ�s��ȮB]�0b��k5�Oph*������]��uXZ��l��H�A�D��o�̷��½Kg.u2��[])�1�"���������V��)l�Z�ҩGM�����ឤ�p*[ľ0��(+Am}�wO|��{.~::m��_�J��3�;�E��۝��g�{D�;&8�_ݢ��]ߎ\��@���
�XR�����N���Ө� 
➮� 
���� `���	}D{Q����p��y,5:elV5Z� o�c��adb�p�P�nU��v�~@��V��@q@���=�c�n�����_����S��v��OިQ�~�_���yp}[ª&qO�^�߀�-m3G�ɤI|����Q۠�|u�ҩ()�M��v^����vU�^8&G3G �P�s]:�W��K?v���W{�#��mWkh�kȤ�����%(.���BX���N����Z�z54��h7$�ǰ�F���ǧe<.^���<9���U�T���_���)��9|����'��QF�B/�@R%�>��?�<��:�ƻ��A����b��D0�TFA�T�B�xPnI���Ҩ)͸��r�c/]��n���p:,��
Eq���gI�A-�.��C��sр4ٳլgH��JhL8� %hG#�^��3?�'�~�J��Ŀ|w}�"��$�K%�̷rbY�(P��c]c74U]����I��洦�{:%��[�c�;D���썂���w�E�	��-W�g�+�N�s܏��^p䇽ޕ�T�u<��Y��9���Ocvn��>����j_�&T���2��jd�9.���j
oa��̸Ҍn��Hg�
�n<�O{��<�����O|�T ��Q���*^������#R��ƷNcb�:��@4�hfLQ���&��*������;SNwu}I���"%;٠'��F���T�$9��M� �y���X{��#b�ϖ=zIy�#ط�:�*n�@�f)B��-D�	�8=��'�.i�ˮ��a�g8C�z!IJ�+�%���d��1���ó8:?��{�[��٘����'O�̹���[e,{�����[�m�:=<�q��(�G?�	,-.cvv�<@A�B��	T�lwE�����롓��e��B��y+��ɑ��ί���Z*�hzV�D��5�:	�l5�a��
L:m׳M��v$i�!�C	�<�}�~�Ǣ;�k���f�3�^����L�`����!N{��5_�]e
E������N��r8�shi�8��ʞ�s/�%��R).zhV�z�R#D��qO�f�Fť+�
�醃H����Q�&���19�����u��jauc�"+e��|I��q@�T���MoF,&�XIGכx�����5��o�� �SQ�p�r���sg��>Aq���/��=g^W륏pN��ޝz�TVZ�̬� c� B��nt�(o ��x�#�����h
A�
�����NW(D��i�8��LP�%�:ݮ�������ruA�(�u�q�oW02>�R��9q�:�u�mG�Z���C��i�-J�}�|�O#�IP��oؾ����B�pH�D9tf���?�lV�����,rqJ8&P*W��g��R�R3<U �������E��D������'>O�1;\8_��{���ֺhv)�b !cN��bڑJ$d�	.�XK��?��ƗH>��`v�,ZHxDE�ֿ��d�%:�=�ڐDi���L�X�Z`oS4�՚�	>3�+����o��1�B6;��W�������8O~jmGq����0aav��:K�;t�f�)��ҿs��D�Һ��Q40=�D<��'p���Q�u�=x������W�R��3�1=}�����6�)�/��V�gs�
��t�'���y�l,i,�Ql8zʐ�Ƽ���9�ڸX5'v�v    IDATE�,tdlT�DjUСSd�9�P8bcz�F7\�,\�З�6M���C��(F���¡�$�%���N��ubbB�Z��d��l��_���������p��>|�#����c����;~Ad|\^]��˗��������'�[��Z\����|��W�K��H�ǰI=����b#����Q0���>���p��;1��r'Q4�e�q4�
.���A�S��%9��ZSDһj����φ�X�I+̄�˖^�JP�޹��2q�=i�u<��?l�mxn���;�������*ā�V @㿚���uq\����D<>7��Zt��bZ4B`l�b�c����Ѫ�1?�G*�E����|�Z+���'�\�r^����%=?���,I��mτm>NS�����<��\9񳹽������E����~.^ƅ�WPkuN���I�P7�@xt}�1����d�c������vSr������0D���]��R���x��ѭmbs�2�:��������㘚���p&G�2�Qk���ʯ����s��9�|�A��Pa�G=./ⓟ��@L��1D�-D'�<��L�TSHk����DJ�P��D���sN*�	�@ύ�С3C_�|U:�]��,�6�6�"��Cg��1'2V�	�@F�aE�,�Rx�㬓�aM��z:t޿.AW��F,�n9q�>�8���`��#�&J�m-p��:�X�=G�Z@B^}�d�
���@r|f��Y�ne?���w��O����~��*���&{2oULX���ý�C�������^|�_���'瘔 |dG#�T�P�,r�F��
5j� �����g3 ���J'5Q�����
uЬn����ib��#�Q��3����QN�����I�{�Z4��F<=�S���2(�*�P jV�EϜ�w�䡦3�;�.�F���������GNC��SS0 !�*7��Ю���,����KۤO��|��$b�Cz�=��]��%׼���K����Jٝ��,l"ܮ��v�y�p��^lo�*�<{��.�L���o��&����4�@M^۾����_[�W�ՅU�K��&X�� =2����>���dP����CwY� S�A)�E��B�xR�R�a���mݺ��u��Tᏹ�D������oر�v��T7�P������-�V�{'0PB04���9v:`?��H�����?r�����U�hX�Z�%1�����	 �h��@H��Y�;u)�M�R84;����p��C�t�4N�z �\�HL"UY�PH���<m��$b!��5"�Rk�̞��b�D�u�%L��XВ�m,�h&�n"3p��m����P�&ӡ��8t3���R4B�VA����#�hU�ѪdL���i�pc}���QqAs��\(
lF6��Hi�8�H�S��*V��U�HZ�ёL���8����{��eF\k��!<�,K3�|g9��4_ʞIT8f#��#��ӡ�ѡ�����z2+��~g���Ҙ��F6�i�OM���Yy�FK�<��F���\�F��@T
�M��;{|Zb�l�s#��g�,_5�pDe&9zo��F0�-�_��ݼgDX�Ans� y�=xF������c���#��r�IJdv������;A^�j+k�TI<�B&�����M���ATJ[VBcO7�q�4�����t�0���a0�J&P�^C6��o��y�p���8�������S�����i~��D����>�)<��B�»>�,�S�{�`�DB�+��,���;t����auuQՎZ���SvIp�f�3���[%��Z��{I�����Z-k�N��#t�C:K��:I~�"Q��Pۛ<�������ŀ�r��D(�8˰�&b�:�.��Z�a��[�^���G?�`rzV��
��c��r��r�3�$mw����'P�6�]�b��|�#YE��9ts�ж6�1�q+%�vU*&P��ʔcAd�Z�)����a�474�-Nye��|�R�b�m�]�0�����Z{`����{�V��w"��	ٱ�>�6�����s�M��r� �Gի��W�<e<���%섶�10� ���]���^��5����eԶ7��~7����Ү�^0(����}�8��������:�BX&7�7|	��)��~��9�R`ˊ�O!����8$���BNS9�~3�{N-�n��8$j�F�Z�tNLKt�������ˣ]��Q)"��"�M�Y���/7?f�7HG��xH�gx��M�P�T
U������X��F�XE4�To�$���9�굦#y��)���1�|𴒗9���ۇz$`%w�H3ɔ�9�N��=��?Ec*�\*��+����BqL�%��;�T*7���mYO��F��\��I
���bcc�vsk��u��Q��cS�'�����uap�Z13����XT�a� )3�2�d@B#��A��uM+'�YV�N�"�H;�����8jR_NK�O��I.��b5=#��a�a�;_��42 F5k�w���ccmS�Yd�A<���Ə<�Y������y+*�ma |�����N�Û��V�I��u�Oz�� 35�������n�p"�
��2I��(�*�<�������C�nsW�6�*k���s�:�>?C�: �$i�w�t:r�����9+2�D`�Ɋ%c�Bc���_�>�z��=�J���NK�8��H��p����"̍���q���Yq�TȌL�С#"?�S��Z ��-�G��Y���]K`(�Ş}7��0p���.\Drr���[,����@�;t��ӡsF��6�G���l��S����F�MYZ�2s,���t>��S����O,Gn�,����=C�r�ow��K�����ݙ��G�س:��č��)�>�W�֡����Ua�C�߫��۟�:�2r��#H[��y}�G�G�4�Ϡ�A�ۣ��a_4A�m9����*���%D�"Qlm����8w�7�W	~�g��@�����:��3K��0ґ��O	jǈɬ�8'ڱ	�X	��U8b�H�TV�;\����ؚJ�P��S�6�h���Kgu����5�A��,2&�cTHk���,y����"�"z�&�R�/5F�ubu
+p�,�tEC!�U輘��C���$�..	G�e���cٕ���\d,��-Fe�ը7k�&T`� ���C'�v ��}4�x&���ulnn!�H#���܍�pr�yISe�8g�t����̀�p���N-�A���ܨݶe�l�v{
���X]^���M���������6������H�����}���,=}�"oGIg�h�t�|��ȱe���߻ѷ�p`>C�ȡ9�IT��uɌG����KC@�7*Kh��U���A[�h�[�3��X�܋~7�����8��I<���k���,���߂��i��U��{�{sGO����M��v����,֥����:zM7v��N�3��5��+���#:t��@@�q��@oEl>[���нC'`�ψ���F�C�C�=aP��+���$[u�U�/Ζ������a&XggL�B��h:��f�UC���X������?�Rt�e<��Illl���#x�ޏ�}��C?�_4o�5������q)^�wPY��������06=�p2�z7���^(:���}��ru��[Cc�sؼ׼�����{�xEݜ�"eX�|�?=#�����e՘��ٱg�s����)�o��t?�X<��-+qU��E0lcv��w���]��o��9"��z�܏R,j-8�Ob9�����/:G��j�+d��H"6�܏ƩNh���N������徶�2�����V}�e�a	3���T�;��\�(�I��c{��3b�bq�cIMg�>\���_~�=�__���v�Aޡ���Zj�N��3�����'�����j����8�&~j�|��G�+�QI���&gI�ʾ)��tm��Hh.�k��QN�,������s0��,�^\��;rn^:7���G����u�a(w�I���Hd��j�C��3ui�����D=yK��sf�ý�a"e���@�����U�R�c��k�E��ΦѬ���`q<jfvZ���"\�x��Hq�D8��^�� K��n$��pf�_q��.~/�X.[)Y�;��ms۬0#t+��9Mpn���a�D�G�_<��:v<��$�.h#!�v�����y������n��` �v�c)���hc�N��O�L���5�}����)�:s�./�ˠJ"7:�Z�ً�jU��JB�&�Π�;;�2�'��1s潣C��w2~���Xrg�Β/��όXa��,���<�*�CHf3Ʀ�sN���w������ͱk�ҡ��H���3�����(�]��d?�������;{N����4�v�7���E�m��đ�;|G�Ο��������+x���Fg�L��cam��I4Zyǡ[!y�:�ܕ��}�k��s㚳�����4�谺
�ͧ1� �&9�6�f~���T�2t��xڞRF��ߡ�p�C���:ײ����q�{���Ts���#��v;���Yua2���_��O>Pgu��C��{߲a
G
މ԰}D�VI@;��ʢ����h�����x>�=�7�K�����f�h@d	י����Qc�t'+�n�hǉE�mD�>m�j��I�q�:�_y���]�����Cokt��#9�j�)��~/�R�,�	���m�T�&�������Г��8�c��V4LIʶP���Jb�'I�fG�;}�ÂY�,Cٍ$]��n(MST2'晡���Ϟ脭�GYW��._(���cf��:y�G��'��g��v��1��OY�b��4�˨��g�L"
@8.�q$��1
)`�#(.z�$���~L�L��JoY]]Aqk[h��o���:us����~s�x��Q��u\�l}ģQ��y��.��G���� s� �5Ə��پ��Y��.�Ԫh5m�Nsﳧ�uC#3�?������͢VX�T.�fa����/~�^:���.*ҿ���j���^}^bd�`R�_����'҉ˋbHT+������C�����5[.2�bP��d����D�X�X���Ls�;�щqAw;t_r'3N�X��v������-�),�brm��;9��9trp'����1��]�T����8qp����4��?{�A���?�O��?�u����ɩ1��+�/�5�z����?�Ǎ7>�?x�W���V3nD��G�D�=�XBY�w�����7�}m/�g�ޡ*���������w�$��JՊ*(���"g
�9㜙R��U�s�W�;`����C��]Nv�����Lm����'�Ǿk|Ͼ���k#j�<��b5��k���=������0��g߾,/��y�j��7C*|�be$Ƙ��s��j��8��K���j �Lc���C)"�^q��X�H}]2@/�Ud?;Lx���!�tV�'q�/�Z�L�I
Ƭ��ʖ�IDU~�*3t��Ʈ3=�~�x�����w�[}m��:�ɱ��e�i=���M����e٫0sN�B���$4l� �mJBrƜ�Hca"u��V�*���´�o�4H��2T�����=шrAr��#���<j{'U����*���B��8]���iw����[�4rc���(�JB^�	�Sob��>�#	��`&	L��T&-����T�4���m�{caY���!>D�n��(x��9�|3��ir��QDK����MLO�+J�B��C�V�� %@9��P1Cak#9�ϡ�R7{i^��υ7�Ԗ6"J,Y;��q�	:Į{��Sȍ� ��2���eF;Ru����v۠�ͫSF4�)�*�^�@/��#�0^q�O�]ZG<���3'q��������z��8n��1X[�������M�'�q��b�1t�1\ZZC������RZu
�DD���z���W/�]����U���c�a9���O�pE���'����ǲGY���8���f-�,$�l�&�72Y�0��uO��*BCX(�i9�q�~o�̱���^2�L��B��ۋ�;��{��g8<�����=M�Y�Q���&���b}s�/_ć?�A���vB63�����1\Z��������Dfr��j�J5��l��gQ��R�Mɡ��Ή���,�k>��Q֦����	�0l�Թ�[��*E�$���k3�흱@o�.�I!����9�(�?�9Έ��k���/_�����L��e7	"SMs';�1]+�W�.h+|���^`W��wD�k���Y�P�d�mI�*w.;��t��~��%�`ϐ��* F !eI�T��yP����ǣn�����?��ū=�jg�IG;ZށM��ر�.��y
��qם	
��1�y�R*�s�gl|�����������|�����z���N@�[oȡ�(���;�"�=���h4������N���-
R\XafE�3��m��M��;ѳ�$�K�N�(K0vp6>@#�4�̜hd݆�#�M���-a'��>x��̟���HjY.Fr\�����V�BA@�0BH%�h���1���Y��ɐ���]��"��������		�Z睭����qdψ�2k+�����٣�K��(;H�AQ�ѲR16���+W/��yiJ�vZr��m�t KHfVπX�P@8��p�܁��H	�fe��X��ҝVI:�7����\�޺��f�ɃO��D�0�[�������JD�y,]a�F��3.o��v��2o:�ů��e�'C8~p�y���/��f����L���O�wމB��7����џx.�T��~|����G��"a�T�[)�é�P\��TU�,m�X�B�c��'����T�,���A��-���)[C}}s����Щ(��R[ ��0�#	n�"(��Hl0�E�$u<�й��<'���Yu!-�[X��!�n�[�B��������H��H'�S|����{��|��w�?�_��8�t��y�韾w�y�t�]���l�q�����w�#ʝ��{U)5z�&`�)З�����0x�z���]�j�~��1g�� ��c�I��HX�[��+�Z���'��|�lf8��cdՌ�C�+����R� zC��,�1�����:L�	b�U7��6 �qvt�C�q��y���W�������;t	ϙ�H��������ar@�T����g;�UW����Z��`���]�:��&�Lp/_į�6�'�}�D��u7��̒?��`O_�Q����=��+�d��*�Ρ��$G�����_������~���oӡ�����!��͍��{X�`�ܓ4�M$�DI{6%˾U�u���?���vV���^��8t.J��H!p:�$.Kh�lX1F����N��c�����;t+�������Ƣ8��&U�����P��4�+:g��	֛߿O���l
�t�.�w@"�7	aܼ��r����
��Aܨ���g�&�p2��:-$v6ǹxj����"����.��Z�,�ّ�Xe6fm9O^�jB�H���n�P@�"\�pF���s�>r���YBp#�R4LpX�@y�*\ϭ��U��0����Q��`��{�ʧ�g�uBf�L{-�]ǋ_�#x��'��O�{Ν~5]�^��#G����.��7�In�[H���]�<�b��@<�V7��#���
�V��(���i�6�]�0�Aǰ4�|�����֚U])n�ډ��U�`�N�N<)R����JE(l� �c�G�nG�'��g&��;_r�#1@�ϟ������w�$�a`?�VU�"��ƣo܋����G�_ř��Em���HA�ว>�������g?��p�whݖ+u�|�,�	�����?�K���3�Oc���X-هk��k�C�-ΖȎ��4����VR��3=$�I\[��ŁO],�������D�+`�����!�Q�J'W-#��J�"�G$�$B����OO�S������u�m�������k���
w���z�zV;�w�F��    IDAT�.�	�H�Z�/0Ti51v��v�}fc���xJ	�t'ȿ6<+ �>�x��!N�T�5?l��N��:�`�_�Ml��t�ՠ�i7v���?o?� .K�,aF8ZJQ*f�D�9��C���zŻ���{�.�V���/��P��;t�}����Ә�8�f�,��c��,�
�W���rԑu ���<La��n����Y6�%nf�h8t�wh���i�#48��h��EFCq����=e�K+hT�W�F� �K����L�X��`Vd�Y�x
�R��.[#k7�qE�Ź���4̐]�=(�_�=IeX�%j}rr�hDz����| �F�tJ#t�Xc�D#A�gW��(��Fa_Ic<���kND���^�2��m"��(hX�z��@r��hs�:�l$�c�������4��`pg�;fCt�T�J&�H�Ө��fb�LpC���s�E����Y��h�"�k��=4Zu$�a�6���g=����D�����g��2�\�{�㕯�5��7����W�A�C?�E:?+��F�$FCI��u4��HnLtiu	�0�5i]YJ�5שԑͩ��ufM���Jg�

�65e�R��=��`ԡ��y�TR�$�<lup��"E�Ö�A^�d�Dctj���Aއޡ/)����M@����]������Qڬ���F�	4�}�{q��C���+¨��U�|�}�~ի��]�|�e<��߇�����7_�F|�k�B(5���,Z������k�����9u�lLk������u{v�(��h���gj1q�"d��y)3`6nBy>��ջ�Va��?� ���5b����w�6^�؅��M�g���	��5���s����ʁK�v�����_��k׉��ۃ*�s���)&UY�F,�#���@��aq�����TU�$�ې�y|�O2E�M����g��$�� 9����^��PE���<��A���{AvY9t���ǯ�z�����9��[�NB�Lq�����D�A��C2��h��BW��0�*+*ǳ�a��;%e���8v��5�zT��� ?�R�4���]	[�%��
�Jh�md�l$��z�h]�$h�҂�����e�4��ӡ��G�1���N��o�pkk���8?��V���}�c8ޡ�Z��S���`.6�WOL�펀#�W.?u�Y[G����r�c�����Mp+
$�Y���H4��܈���%kd��\t��BΛ�:#l��6��B��$���)��h���	�4�C��������m `ee	�FMR��v �/-"�o;9��	OcQ$*�F0�E���gї������3��B&C,���>��gH��XX��J��mf�#�����ٟ�)�_��hr�^�d�	�U0�@��@|u�N�����\YP��l7�vTr���'��{�t�L���͐��X��CH�
���ɹ�����/gbټ��/(�L�l4}�߲VH<3���~I��)�F��P�O�� U�Tݴv�ٓ��RB�R@<��co�����a��|�˟�m�� ��<uZBKB�PQka��y\]�*���48� <s�p��K�/��<�-�"62���[��9P���5e�k%_e�&�U�0���^_�_2é������3bX�`�����+,�Wf5F�V���!� ��/� 	�U+Hg3:~������y����Ys��X�ݥy��f��=�UI�,-(������z���1������v������:,������b�/���=	��c���9Q�ׄ�ɍ��S����I��6���aŎ� �4���Vu>�c�y�й��V�ů��)�1h���J�UL��Z�2�@c�_��N��@��n����6��ʦ��t�d������ֺ�{�B��ZHe�h4�aY��K.l�=2S(Mc�z][Z�Nw;t��͞sHY �x�;��p@:I����#$(��>_(�~��q�'D9�6��+B�sY��� ��H���T,.f�H�Ξ��lj���8p����C����F��DO1�6��]��\%�nW:�t�s���3��|NƉ $��:K ��
 ����p+�K⾞���7��,�	�p.W�4�^�����o�;�%OhT���%�OED���/c�h<�:�ǒ�9%�jM�W����;�jD��C��F�PC�T�'K�9�E#���dy;���X��6�+��[ Das�*"�>ҩ���r����� �&&T�__�T�[X[s�]@";�XzD
k��H� ��N�9?;���itQ*U� г�F7h��JYř������Q�P�
�0�K%Q��)��9�F�)U(�	u����}=��%��m}�V�!���9�߲%��bȪYmf0���;9�~�!�  !lW���k����!,_:�#�g11�C��-r�Lv�Jӳ3��(�
�N^^^��c7�2w�؍X�(�g�/����	br�0�+5��Y����[���n�>�T;�^��֨e�lu9�����8ȃ&�� �/R&��)��1G+���ǂ�O�8�C�*R���'#C�i�s=��n��;�A|�4���`=��ϥ{B_*̧��S��}���n���;\T��ip^V�.�kּaE<'�1�K�3p-gI%>,���T�V126��^k7��~bE.��63~�Dª�������Rf�vF6e�_�1q9�Q�\����:m2�[$}�Ρ���Я��+/�������y:� �,�&3�rw�%w:�4�e���.���y<����������T���̭���.%��k^;ݔ���de���ȧXX&�hI2G	��i0����pVV091�����i��o�Dvd��PmVhH�� 6���|7AR�~[$:�cB�Ǣ=���'�?4�|�q��Ξ��h1���� BD��2��i�-�1|i7` 5n ��D
\Œ$Q��iJ�~��YDH�CTf�F��)Qn�//���*�g��u8����U<����vͺ�c��etl�O4̤።�ha��A#f�e.�j�x�	t�1�t2!�lL%�yQ-�tkx�+~������'�����Q��Q��Q)7�1`
�d3ds���Y�v!��9 �^�D�:v�.��=Y_]r�Kcj��=�ML������1I^���
?&~�j��^?� :X޶��X	V8�Z5��İ��",�)JA�'���w,���W�.��g�2�]�N���!�&�i���,I�,� ���q]��"�F��
��z�Թ�rSwە���8ǡz�m�����8�u:�~��7�C�QB�R����6��S{�&�}a�\
Kˋڧ=�9�ǰo��^��l~����latf�jݴ�w>;��g�
Jve�b�cO����8�>���^)Hlh���t��"�4�JJ�W���8�3>~ԓ��7tDq��j����!ft@�FK��� �X�ұ������yۈ�#��X��O'h���Z��)C�����u�������P�ٵc�|v��7K��j�~#�aPG "���~`��`"ߛ���
��'K'�h�T�jQxOMLK.U�t���
m��Gdi<������1�6lM�������cŒ�A����jď'���gt�x�W��3��U����.B��8�VWWus9%�ᮔ���06�Ư���@���m��o~N>x�����vT�i*���FV4:ol�˿<��a�8����ʑ�A"���Y���1Ұҡ�m�)�ZU�K�x����x��XY������"=���Q�(!�/.�:35-#��E�\��o����.�Q�:�_��?,�	����	�p��9LN�!Ƭ��79􀜥	�Yt�R>�4�Bcξ1#�RY`4q�G"cb��3@��d*�T����f�'�����O�p��R���&�lT����h�4KYF�a�U,OONM-o4�x:��	�_,Ir��]�]A!�p
�x\��7j[h6
���y*~�E��ѫ�������>�` ���m�Ci�����L �A#�����QB{1�fI��t~�~�A�Kkx�����X�Xŗ��%�>s�zc��a����Z�\_���#7(HZ�\C����$���d�3�u>Xu�3���I%�~5K�6ry�؍r�w4"��Z!t�M���!�J��siLNO�u�V�Ʊ�0ׯ�i�:����L�F<����:��:�9��G��P�`�~�I��A�q��r@���$��F��v����G��T�ۮ�	��1?>���Ƹ�m�T�2�[ő��F:t��:|�,, �̢�`}e���գ�*�dK�$�r0î���ֵ"\_ܘ*� b+�� N���>���ſ�(_$���G�Hj��ڽ�f�x��[����}��K�<��O�w?�ɸ�S�Ĺ��wO����I��@���+B�7¬e8���!l%�������N%wv�fW�6�l/k�$����|�ʜ�yԂlR�F�`��J���:�	��=�@����x�)nT��s���Q�C-�����3�ҝ���6��]@b�$O��?���`���(���1�df�t@�G�8:����_y�]��F��o�{R���D:��d&G�<�8��d��7p�cn�/����j��G>|/���!C�G�C�n�)�˺T'#��ކh�D�W/0��k- ���Ƥ`��qRi�E]F���D����IbСzP��$��^�����ш�'?u�W�C ��2�t4*�K�h68��Uk���s���8��������ɧ ��7�7��=���o��~r4�d.�H�FY:���4�;�L�{h�ے&\�tQ���"�I�Y.��py�F���Q-�c,�@asScyĢAT��hTʒ*���x�S��o��u��iسb�H�a��i�j����5��*c�i�<-�s��b����me��TSӳHR�Ԥ�
$�Ȍ"5���{�PR�L�N�^���������W��GƧ?�Y�j��ST��z�t��#c2D�r�J�t@Aε�+7���D��P����r���#�����w~ �y��Ui"?��P�&P�Xߔ-�C����'������x��Q�UNbS\�M�^�T�z=YY�.��vAkF(j7��RYJg���p8�b���1�VW֔���Oc���\<n@.�s9P��F�I��Wߣc�.Z�IB*�Q�D��jU�Z2��l�"�a'4�E&F@h��Fժ����C�'��"�����o�E�A!�6�ɘ�}gǂC�7�@5����Z*Ԇ4-���s�I\��Ø��(�笳��w��!U�c� h�/	糰���''���L���Ds�#��� ��Q#!��^����p�T�w�4R���*`����7ï���"�6��׿�M8y�%��qQ[<l!5G��#)�O�A?~e�C��V�����z�����)kM�P�A�����(�i5�XB�s��ن���$��lc9r:r5B66nƵ���q�O��Hp(���q�� �lu���M�$�����s<�5WVE��lc��
D��ӁU�J��x��d�H��Ɓ#�˞6Ŝ�	^Y5BՎ���bȩ�o��$3:�~�e����z�]/����߬��{h؂����#f�q.O��%ߤpK�l������O8������w����A*3�N��rs�*�Q;�9tƹ���M� nS	'�v��p��{��F����͡3S�j��a��-�5�a8�H�y.p�m�>e:�����s��	����?�E|��_C�F�Ʀo�\k�k"A���P�R*h��%����"��^�\<�_�ʃ�؝�Ǚ3W����o��� d�e�����<�Hy=�4�D��Q�[���(�I��om����~7�4��"]L�&��
�KhP��F���c���C'%�Q-�Y)GK'��X�=�I�04������D�i�e/6
cmcSN�iO&���'����-�t��ø���#��}�V����f+ !��:�;����������Y���8p�j[�j��$�o0� �|�z�D�;�6��>��[2^�(Юl����x�O<��E���~�^���"�cs'G��Y�v�d~ǎ���@���"7��4z\tZtL2vΨш������������˹t>ó�
3�\W~,�[�σ���HD���cf�c�ɴ�M� �r���]��?[��2o�l6t�t�|.:��9X:/���l}6⍟�<���N^}~b��H�5σχF���k�Le"�Ϡ��U��_t8���1gF��5�	��瑠#fK��2o�`�F ��$ێǂՠHH�IVQ(X��`P��fP���|���e�7V|��mU��ٌȔ��+�����\G	r1x=�.��t��Z[Z����R���Oi����ħ>y7���m^P�������ࣈDSU��\�蘭��{����[������(��ē�?�'��a�D���` K,I��)��X�`���U�V<�l7N�ͺ�7����Hyj�L�A��a/ %�n�qe�N� �b����H�`�UAU��G�!8��F&�R�>��\C~4zǙ�`OA�5l���<n(EP�u*���~?�w���K�vf�5t�ʚH��lˡ3��7$����t�@8�G��ūHf�Q���Ɓ@R@*u@��J��hH��e�TN�L���`P��ze`�.�����F]�4PD�"fZ~�E��F�0���	�C���	$�!uK�>�Ͷ1��*�񵺼�J� ��*g���X	i���#I\�zJ�2V �u�}�(T�����#2x,�R�ݰ6Fp R�``p9�\��bG
�c���;{�<��*F3cȧhV6�on���
P~s4���e0�K����?��7�����ѣ��&G�Fq��93�n��K�,���*:tf)T�c��$"��?y�)����O`nϼ��/.o�o��Q�:�y��Ez�����+W/b��C(TJHdrHgG�ੇ�er#j�P��e9��,��V�c%�AڹO6��C�0=�����$�A
�������l�k�9 D��m�np������F<LtG3��(՘u��ƚDvQ��X�eڑQ95�Կ��l���c�u���Ҳt0<3)j�=d����q|��N�N������i�	�c͕��P,��Ӱ�j]���ɾ�S���Ͽ�g�>{F���(��
`��h/h�©�����BF�A���)I�3x~���d@��1�;�8.�38S�j�~[g*��r�aF$ȉ������oasՊ}F�A6��S�S���-HYY^9T1p9
������=eV���p��/^[�^G��uW���=e+�mN��./"?��/��K��'>���_���4._a�G��7i�ޮ��7�B�uL�VO<�G錋�:h-�@O��^=����Ȏ�����ϝ�q0���]YZ��f;�NY��AV4�:.χA���L�	�~_��}UE�����6�Av�e�bxt
�:c�L��;﯂MW�,�6M�	|̩���1�5x�]��V]�Wg�i;<�ߟ���K��ޏg�{7�5�'E�8s��]��@�}뻿��{�.��މ�0F�"`O:�}��²I|j���A�:",�N��h���I��Ud).. {RF'��y�'Gj���?�P��5�&y���,�i!B�rfs��N<f�T���������n�,���8��JV�#k��9B�	�m��6RؑLVי�G��0#f�;39���q����e�\������d6���#��()���9*����{b���ˋKȥ�⏟�����&6ַ1��#�02�B���ᇟ�,�WA6��X:��&�g&�t���Ŀ����u�o���r�ܸ�\_���ЕU��9��ژJ�YU0���8�|�-���$f�����X\�Ɓ�Ɲ��&N�_A �@�~�d��8��	J�R�'���e�Ҭ�ם����ᥪ�ט�-��E�C�h�cv��N!��7߄�o�����g>�9��߾��(�g������ul��㦛n����&��ԑ�P)nH7����v@�    IDATAekq@�i2� x��'��:::���K45�''-�#xM�mD��F��D\A+�u����݂��q����fY�_U����A�OG�g��}iX#WN膙1������>���{	H� C�^�����ê��
��T��c�SA��LCW�\|K�X��c	
[ֺ"������-_` �̝�,�Y��2Qϭ.R��ew����k�sT�`D�Y9�>3���F��i�+Xq���6�
�Y�X���� ������r0d��m=7����Ѭ"�d֞i��:�S����!! ����I��m -@ҿ4�A����Mt��-�G  �J�$���Bì��U�+�.�+�����(�ط���Y�ZI��pU(�\�����m�E�INJ>�Ϥ�R�v߽�g2E�{DN��<��F�F���HZ&��g2�cŁ����9l��h�ī��Pd=aK���+�$�r�n��>�c0��"��6�%M3	��GP��~?�����K�9��f7>˒{�g:�#*[СK�K���I��A&I�@GM��v�f�sL�*�(��'@���q��j{���M7fG��զ���鶐�r��Ju͎9tF�~�+����9'��hhY��d"&b.4��P-�
(3�v�a��f:��A� W�抹���ݳ�c���T����v��N7��߂ѩ1�n���o!�`������;to,��V��Fr
+IWʌ�^kanf���1*u%�(o^�H*�~�$��T2�=3��x�Μ�_-�7����g~t=��"wf-/^'9�%Etx���AVk#�V����m|�3����x�R�l-đ�<�v($��g�n����z��~����6g$I��(*պ���?��"\i����a�*�"��5�*fk�n`z,/��T{�C�Ʀf���)m\θ77�G"��-7Ʒ��,�������,Q��ie�BQ����f>lA���ec�S%�4K�t�t�tD�Cp]13��#S������x�S����{�������ku1��ґ���4��GOc�yʽ�亥�T�ա�5����L'E���H��~�8��r�<<���_x�jј�V:�P��c��ŵ����D^D¦hTƓ{��b��5:c���г�5��?�s���#{�F��t&�Fr(d�f�Ɲ��y�N��������P����M�3w�xY&�ؕk�N\ ���z�4IزI"y�1N���P�}#��5)�M�oT����}��XV����
rĴ��6�?����`p/r}�9�	�	�#v����6�E��-h_k��4
x]
H�\��P�pt�_����U�vf�S�'>�����x|�Љ���9��歖)k��
+����F�Y�	�,-�YǂL&�%�j%�jɻ_f�bf�>���ɉ�#&gHH���h��s��y{�Š�1�iA��(cq���N>�b������O�{~�7���RO����Y[X"�'K{�6�2\���ED��Q�A��YN3P�Z$1F��TDC�Q�mayeA�x#�IT�e�HTh"� "��fۀ>�ye�-�6=#Q�4��!��y�JDc�s�Zht�ʄ�	�Cύ�w�[2��d�L�FXFӁ/h��
�2#����%҈��hD�ݲ|h]��1��ǵ����2VWV$C0�޽{����J�*�NF�p��x��t�����!�o 	�^)li��S�6kX_[�A��&�����
���}�l�СC�����2�*�:��Y���a<p�{��?�r'�Y�5qaa����Ma��E<=�>��������5T�e!�X!�B,np9��0S)�9��!̀h�0jTό�TGxA0:H�O_�@:�,�֌O͠\oav�i`Ӡ�*E���<[����o0�]+(Ü�߃K��Cn-�lnn�P������L���rt�r|�l���7j2X����
��J����S�N���L����t4,�K����y����?ao�t���9�~zļ/�������O�&'.�1^3(��v%g���^�����J�絝s�=k�#βԲ����q2�1�m�u��' c�d����J�l�I�̕�`ӯ���v���'�MVA,;m�I
�I�[7�!�Y'�ʙi2D!1AM�(�LR,	q��X�JU�6��t궎я�Y'�>�ӈD9?E�����	��+" �"'}%.��H1����S���N{ů=���6)���ET4�e�)�k?���������g��H �q��J"ۤ�>����5�@�*���~����)�pRI�:
Z��qN���5Ե�hPʗ�F�x�3����"�7���z膢h�60�FwĮ�dk���ޡ[��KW�/ �2i�}^�:���/���ګ���t�d�Kui�FDe�z�*���r,37F���i����,Z�rA�;>�W��7�'�+)ժȤ���tJɧ06�r�Z�d�h�NQ�c�Is�ѡsp4��%q!x.pC�w����c��ca��2pISV�ȍ�q|�4�5P?#~"����C�]�ͧ�C��d���.&f�"�����"&f�hv���Zʮ�2�Iұ�������{����ss�2��Z��S��ۏ@��^��#'�/�1�K$��sI�z�>왙R�J�����͚I����oq^����Q�:�k`���:n�a��9h:�����|&n��(���ON+�������F_��9lT�hv�$�B�@ґ����F��Qb�@�9jA�G�*v��e��3	�����N������������
�-,� �Ψ|ǌbuy�`#����O��s������X �&I`8aQF����z�!fA��H�1` �R���-�R��q�^����}&�K����\����%
\��Y�v�B:���;t>K��q2�f��ߥ��A՗aeQ�,&ty�J�^^t}��<�[dU�/^�����%Z��X}٘��ǀ��~�#�eʋ܇<^6m�BVט}ҹP�p�Z�M������-G�����������T�Α"�,/k?+�i��"+c�:���#�s��!������-a 8�s�(p��pO(�����af�ܻ�ֵ[}e�M���1�4��  �k)�H����)��X�c`���X� �@�c�gϝ�h>��ft$�{�
���F�ϟmH��"���6�iˀ�LV2��	s���Zѽɤ�X����1�M�!^�/ի����j��@_$�i>�Q��*���|6��1T[����ai}�%T�=�Cq�
��F�+O��G�����Ǣ�����^ ����p^�%w:����/�̷έ��ՏMR�:�nɡǍ0�Э�ʞ[B�w�;U�m����8�Nm%��E������T�"maf*�������4���O��O|��2�0��E�]=�v���a"�K劜�"�^W�D�ڙIV�F%���hG��; yWfC�B���(��:_f^�I�R��ei\it�2��eYR�*"[I��c�����<Z�h ���%!S�ݫd\��6��<�����-f|�sӸz�����޷g��u�7��߂�W����ͯ	���F�)TJ[�g�HD��6�����g��]w�����^��3�HH��IOz��6*78���@>K��	|ޏ����{�7u^$T	��H��E03���]Xܬ�ѥhKl��(Ƒ�Vd��6���G�	�9��p���V鮧)R������mS�<��L�a�ZMR��Ȕ�epBn}+��'h�%խ��q̎�P�^ƕ3 ���v7��#�%^��2{}4�\/t��F�H��Ñ#G�;���yNt����ǹ�i�����,Z���5A�L�˯<��-Q�p��c�T#މ�������2�qX�����g�2+�`���w�7����ٳ�N�3e.��F��x��2���j;�����'��儕��g �2�;�/�	�3����<0����[�;O 9v+N��L�r��q��<ٻ?q�� �%<�F�ػ��X,z�L�V[��?[�9�{��l��1s������޶�=��pŦ�%̔�=fCH��Ns|�@���)3��u��+��\MP�)� �-�:�Ϗ?��ǎ�s���$��,yox��1Uo4{o���Np�\�[[�x��e����:{��J�Ƞ���J�V��xJ����5�|��
j.\� ��u�f[�J�V���߻D(��Ozʓ�y~ˋ+����E�i�G��D8NQ�>�<��Z�nФN9�ħ�Uz'�;�;��9?��*C���;ؔt���.Aqt���_��{/m��ՏNԫuD:�o&(�e���W�� ISiv��s���{���蘘��ЉZ��7���}T�6^�K?�G߾�mO�y���)��M�1�c��(�կgdF0RV���J�dts��<���T�"�#���M#BBjW�Tx�c�Ź���cGo�F3�VTJ���X�H�Fpey�h
+%����P"���5ē��\\F�!���U5�D�ZI��3�E�8��C���؎�� ����U׮ �cf"�Fyc#)�V5!G��������s�p��G-���7#�]t�g������w���|�p#S.��c$�w ���IJ�����]*!����za�ޒ%��j;-�8�M��c-�=ҡ�g�r_Ia*��Bs�,=��U��1�Hg�sa�ǗR�ݒ-!������*R�B���O���~���&GP�\D�]ӱyݬTИ1��⋆���h��Ј��W@K#��ʿQթ�н��"��ip�=�>��fS9lo��%�s �%ׄ�h�=�l���oEX�c{f1���K��<�Q�
���g|v����p��������vog����4B���$��xQ�"W�"T���)	-	M �J%��F��v��N����z���x��gý��e=�~��k�5�;����~�wX��x<D �9���t�bXk3;k�#���\�z��)*�̜��V<C�jٌ<}�����s�W���[@์�1�b�;QY`3#`�tM�8؏1��B�q;/�G��½��/��	�Y��iP���Ҷ>��W���X,���!_O�q��j{��VIЂ������2���o���C�-"@d����k�ڹs��禔�RNh<�R�bF���ujꔶNn1Âuπ�[p^�C�?�yŋ}�}��/���=3�c*2���|8��uLS-B�̳����1�����v:6?�^�'=����[���n�m#��/�H��������g<�6�(���a�� ��ظOd���=��e��[R�ЯZ'�b����K}����PNG`>��%���Ө:_" � d��Q��3^������O�����������[��0��d�e�i�b�-n��Q�ƆE	ĺA��}�:AoU��L�2�Ԭ�!�5ޭP�6X���#O?�������W>G��t��u�_�����4Z�ie�`���Q����pf��83?�=	�d�N=�B�0
A}�%kz��-���˿4/�XLi��c�@�	��C���|�a^,�x.k]��[��ܥ��P+A����E�L���oF%�a����o�:Ҽ��:��H�6��- z�1D��N}U��Ym+i�hA��R���E�:�-/�;o���)]t�j5���x�_g#�qٔ4�ٱ�L�"��{Bcc��# 6�_Q������6>2���jviM�dA���z�����j� �	��i����雲�F(٠nC���?Fi�6�@;��P�����f�G2[[`����H%D���V��p±xWՕE���]���_��Y���F�Z^8ed<̳�Dve�>B��1���OS�ҵ+e@�?ak�9���ȉ�<T����d�ǇF�ϕ*Q/!B��<�6��x�s\��Ɯ��F4D}(��A�D�F$Q�9 ����-w�H��/sD�By�c����f0�hjt�����[�)����PN9<� Q�Ŕ�Q��M��_Y1�bLs�*��N�<8)<��쨑�GP�e���v#��-�a7�^�� '� n�wx^x��a(�-e��`(eꑫ��J�b	{�@()������0}*ZY]��:�#B#�,`�.z͈� ����zc�QVǽ�Nx^��shF^*�x��7�0��1`|�<g��5kCLH��A6�;Z7I�x����Am��ʊ�߯J�qy�l�������t��I���h��
#��<htxX}���y��(~�����P�þ3�1Y�?��l���ҀNL�+��h��T�0��fG�ʈڤ�t�LY�#ߌB�(Qgm�]�#�R@؄�$������S��'�B�l�_��-(�N7;��^U
j�H�S��
ݐ�P��ZV
8(�`[ӻ@-h����= t	a^9p"�R!8���/9�Bn���k^0݌r����I��S�:�n�fau<�D/b9Da��Y�Bf� �BӅ����(ݫ^����׃>h
뵯}�	��o��ʽM=��z��.�P�Yg��s;=OLj��J#����:5��FF"mM54��A
T�!�o%!��؉X�[Q"f^��a)t�����u������:�8���*�`cj��$�������wߥ���U�R���n���cx�^d����͓2�M���U������NNY��/_��:묳t��س���Uс��:2�n
}f���NR�k �ǵ4;����%�����O+t�;��3o�{�S���cǛ'd�y��G��?B#�������Y[Q!�S9+m�S�[�cޣ��NU��fB��9c	������M�!�X!2�����Q���V���P噝����@���8��!�+5Mp��9?�^���w�I��?�&���!hzt@Bńd*���������1�y+`X�u����w��!�d��m��w�!Ӏ��`$3f�Y5����r��-56:l^)��O��TJ'N��j����ޢ��pM��"K<��p�{E)0n�~�cu�h�{�ʕxR#���]שּׁ��d�%FF!~�۸0�x(Y�E�� #��X�R���X� ��⼭%z8`�k�-Z^�ZU����|�����ذ&\9�����PC��� /��Ȋc5XϬ���9�m;l�<��!�s��Uu�A��߳�3V6K�8ꛭ�ur�S�7g�H	���Y*�"3�J��ȸ��W���ِ�c�!,�����F�0:��ђk_\ԙg�m��z�.�*]�S�IBA������Z�O3)�Ri�9�5�4G٩Y�V~Y��H��~Z�O�ܩ�ِn@�=�:!�~�7?ph�]�^f� ;䊪uK6S'��jo<��
0��E����))�������t��Ŭ��Pv��Su}Y[�hyiJ�R�z\��U�-���Km-hy��N���!�X�t>��F;X�lV�9���uJD��c�����v��fsaa~�Ƀeaq��-��=b��_t��������/U+��R=��|��Z���W����Q�l�l�.-��agh(���)46��l��/��ưu��	k�b��DW�d[�|�.����-�y��z�EOQ�YU�N/��)��ڪ���gt˭7kue�j�/���p
��w���ԋ.����;�zр�Nؽ=|�rg�|�+-���C���@����gj����~�n�����Ik��1R��Ҫ	lT���n� ������g��Q��u��jo)�i���� xOЪs��J�Q���eC9XV�C��{�c4�X�W1S���s��jyxL[ǆT]�Q�B�C����􋟮�?��f�=z�*�(��{�~S.¦�l-�#T��2��(Ϲ�fS�|#���9zI��&�P �~����u�=\�<!��r�3a�z�l�=�+�ّ��e0ŗ���̴�f�-� E�1��\rI �)����o��>9���1��P���3r���QH�-Z]3��FS.0�ues����V��3o|����/�0�0�� ��I�C�����t�O��n�lN�7~Þ#�t��O.�a`��L!}�;��ԉ�5��Bh4��W�J/x��ۜ�w��"���1���k�S����fG4�M3t    IDAT������Ę�9jF���$�6���:��}��_��͡���]3�׽�uz�s�c�u��?��%�i��뮻ΎaK0>/	|���ik�cQ��sf�2����{}���g��r.�.c�Ї>d���x�qV�yj�/��7 ���q<���_�N{n�=�x���hԮ3�����3���旭1T:W�&Z$�(]#��ƩL��>�9������Y�1�,i>���IC�SR�$-n<�.�xR)�c�^p��>tp��-eGjkU�5�k�Щ�<u�ա3Al0��)�N@'{��� X���ڭ�T�p���fU��3$�(aɃg��W��M%4PHh�HE��h��5����M��"B�J#����y��r��ow��/��+L��;�� lm�|�W�^�E]x�E���}�h�y��y��ʗ���r#�k��QO�S��-�["�Fh�@^ A%b�P{	C�Y����*a�86�����%�A)M3��K��{*��ڱ�O}EBH1�:qX�<�����=��C٠��g_t������،�w�6����{�'6P�h�533��;δ9����c �X�i�Фv������TUN�x���[��&'�(���m]�֛X�t"(DL �	�.�n�xd����K��!�ijf�����:�|vnYtQ��WØ��)!-B�Q�먱��.��꫺���9vP�'k���V� 1���<3�H�z ��Ba3O|F3��i�>�k�.��o|�	#s����yG�&��Ю��U�#WĚ�wK��sα��(B]7�L���dp�������=��ݜ���rqO̄��+k��[~���� A�}���i�m���>n^��Q�8z�� D���;���|e#��%Ng�}����wY�ɯ����֘�����|D7�x������܄�u��/�>����{,���2�d,m���o����:k�%t�K^��#��Q`n\�nvt��3��ꫯ�=w���(�F���^��ٟ�y�o����A�3���������b��V���)��U��]f�``���,+��v��aڶ�/��=t��k^�]u�U��s͉�m]����կ~�F�:s�G������7�)�Y�4�u�I�׽�+�Z�͉���=�y�^��W����;��9�o��}�oZT��c"�#���|�~���i}0aB�+Dɚf�\y�5;3���Q=��'Z�6ԍ%�A�J��Re�HǨ��u[����|�SOf��ik*B���ݦC$\(��ɓn2�\�h��I�C7���o�C������
=�l��B�:u|C� JD�o�<�ytyh����u:�S����͚:��r�'��� ��n(_Ω٢߲r��PuaZ�3'�T�������BlxfdD�=� 0C���Q��������:��sM��(k�5S脾٘ ^��Y��w��?n�sL�2�镦:ɲ���֝�Wߖ�j���dT��r>�[�B��E�M�ȅ|��5�k�(��r3�S��Y����1���+��k*�����RVՕ%�8zH�S�y���<���\��%U��j6'��c��~:`�3��/^�fӄR:I�*���{��?]�����#�+�����<�UGNNi�o�Z���4��UX� �H������H�z1�S�K���Z���45}L}%���ȑc�;_]�9�����I���D��,��u������$^��	�c-]x�6�����wjJ�V�*����n0�>ք����y{�[�bQ
��ں����}�몫ޤ�'O)�H���:j�Q���a�y��[��ZU��T!�����?�i+�#7O/�_��J��7���z�ޠ�����w{�_:ү}�k������,��;X����^����'��@�^��8�ܳ���o�Zb� �SǞ�u��G?�QC�=v���Ĩ��'>�	�}��A�H*nƝu�IM,i����ϑ�f.�g_��͓�%Q+{���n��VS���?~�պ��7���uB�/}�K���>g��L��7�]��]ܪ�)�����6�q��¢�4���^����ր�SR�N��(D�n|��7�Y��Ϟ{����կ�����r�J�``n0ެ�d"f4�o�ݫt���-�Z���|���_���x���IA8�s���y1Nx��u��-s��g<�Y��?�S���D�o�q��g���[��V3B9��ɍX���q�o&(�����o>`�Ǻ6*Z��_�"]���C���Zo��Tħ>�):x̺0"oZ=��EM��kfnA�bIM�"�:x�_ԥb��LY��p|�*^��\P�F�00k:�W��gﳇ�O*��u��ᡣ��i);�B'�΢*�Boa~�Ѝ$�M�4��C���XF-t3�����֤y�tOkQ��$�Z_�Y�uHX��V��':�+g�QS[+Z�=��G��aK $[��MGÂ���+�՗[)�5�5���k��_�+��e�]�m[&u�?ҥO�8t_��6%C�F�Bx�<;�m|b"����ߩ����oߦ���
�jǳƊF1��Q�vB�+K,W:�u�R!�B���`��A��T;���um�ܪ��ұ�)�K��C��oѱ#�͠�2>�Ǐؼ��Vt�]wjz�)���[&���$.��\����F�{��2�-[��+㡑D���0�ȡ�vg�}���A�.A3����Gz���b�>�W֠���ؘ�ͮҹ�m(�7Vk'jѴ�;F�I�R'fy:�~�ƚVVgu�S����v��l�n��a}�K7jy��N;��jC�gl32
��Q��wr[�F����)��k��h�ݖʙ*B8o�:YZc��������/6�F����y��wgax���4�׿�uz�k_g�Q��/.�[��@���˿�����SS�A1����o�/��/Xn�2�?�0o�[o�M�_w����L�ODg���������<Sc"�@iXJ������=�t�M����Ͼ�K�袋x�@)_0J[������t�-��3����k�7�@!�YC�z�զ(����xY���q�v�w���t�]wm��Hϐ��'Ș7"<�����w�k�ɮ ����^����/j'�1�#��;!w"rD3�S������I�_�)�L��Z�àg�
�@{�fx�k+v<lr�����7���}���\w2`H0va*���ݪѶ7��0��W)��α�$J�5Z�0�`��O�{gx�I�ƃ�ʱ<3��^!�W��xn�!�b���q�Gk���}�ȏ��E�)&���(S�eX; N~C��3n`Ң�AS�ҕ��v�ܥ��?a)�uk$�0��x6c�g�B�
d-��	��Ǖʕ�y/�����ܭ����)t ����N����������w�z���Z�Wi��TO�8�DM�R�R7V��I,�$g��)��ܪ��\W*�Q1W>�6�"=�!h�t��	k�23?�����T�imԩÇt��~�i�amk���⥬l�K�k��Uo� ��Vh�:��җ\a��v���g�aBp��Q{m�%�k֨RɮQ����Ȩ�}Ú[k�7߭��]Z�������)D�0ɘʕ�:I��b���ۤ���Jێ=j��!s�RΗT!��n(�ZU����^��Z_�S_9������.~���b5�K���>���6ʕ�����LpaH��Q$�?�ӯ���<h~�a�_2���x�v��8rƄ��Ƕ��Ǐ�4�M����ubaU��`h�Z<�� ��*���aej=��ti��6����#B �M�^]���)�����~��.�������ݨ�n�S�j�Zf�T#�lݸB��єR�6L��kjW��\_���a%�MM�:�g_r�Jٸ���cF@AHt�9dyh�\����PV�0:޽{�i߾�&�Y?0�`#m�7اm[��2P1��W2�AW=z��-��9��v?d���VLf�PN��9�bP� �@8p����{��ff��X�P<N�A���)��6�9(
�H�焭�A�f/��|�������sȓV-Ε������D&�n�@��qv���f+0�5@�G<�`p]R4��1�0��s ';e����?�\^;�3Jk{`�\ܨ8�K���YLn��'��2��]�xh�"� �#}b��r�}���FGH�93=���wX��gG'6/�[Yeo\eO��6�^�ci�M|�ND���"j� �v��e	߇�x����}[�c%��oT?�kk������&���8����� �R��0�KD�`�é�=Ǹ��r<t|ެ�(���>+��/ �}&�b! ����
xpxDO�s�������N��s��lN�g�U,�Ԡԓ�AVe����pS�R���6Gς\Q�dΪo؃O:�;��|�?ߴ���4�������� ��}�g�a$�,%������ȇP{c}]��j���+�i��NsY������kJŌ�� Iss:x��I�����*�(����GԬWmX�ԟ"��5z�,��k-b��a� �
E��VK�zֳ���߼����%��+��L��o�,s�3���	+7�*��Pk+Y�7��}=���eK�%3�VO��?�cX԰N�3�j�f1�����,֩9�7��h��Spۯkh0���!�5>T��j�\J��:� ���Sk�Kz�G�;�J���`_�!��S�-����!�U#f�;�~�2��9F<��^��U~��a��/�`D�ʠV	O��~x����^kiey]�LY�Bž9��e����"��$==l�-ct%
�ψbZF�ܟ{���W������7��;���[����X*���1�%���e�{m%y�a{u��o^��?�Z�_���ʹ����+u�]��_��}�=p����Ep������s��v4�iR������h��ɴ��Eh�	�ެ��+X�Pπ91-/.�P���O��=j�V!Z���	QD¤--,E�!u��ؽN���^`7�8'���RH�.h�T�?5��zw<+�;�f�f و�āb��X挺5j���t�`��t�� \�x��k�T�1�>�N��`(!�P��e�$˸�>���;�bqaY�#�VҴV������>�<�nG����1 @�ܗu�"�a=��1�����>���9��q@ ��T>�I����6���y�;��H�v%T2p��R���K��|/��R<�y����0﫫+F��������@R-QC����^	�/�/�/7>�>Y�Z��r�?��]�&��Б����>U�J�O"֖�Pֳt;���-X�t^�dF�L޼�.�����M�h`L�O:�o>��7�9��'�Nyl����C�,`qz�6�mjX�@�@o���I�#�P{.J��ꬮ����?�R����:���+����Z�N��?y��	YB�P9>���u�F�j��,T��@���ؔ����� ����IPT�F�O��g���LPvX����-gS�*���KIK��VK1O�P�oD���)�)�40�z��*�k{H?��e���1rcԱ��N�'%i4��$��J+ե�M�h��]�[�� ��)_H����J_V�'Gu��ǭ�<�(�I��XU������)����q:�%�.���7N�k[�,�G�������4�Ɂ��.-��#��4�_<UԹO{���LO�� ��ߪG~\��:ݤ��@�����u:f4��V�<-:e7!���q��wʌ.r�xp���ʚ�|Q}C�j��:�k)�V�J�NW�^M����T]��|�f������߹I�=t�^�����ҭ?���5P�Zl�B-7���?8��������V���B�F���!����(��,�m:ه���RWH.9�����O+K��+��:�m>��)�Pp����!Y�,	��S(���lϑ�^v��̑n\@�k5�Q�=���/r��1g�Z�P��~wc�{�㚼o��h��0rC��8�����WH��ٟ�%���h�bv��#����Z���?��_���s�<7��(�6gN������p��s�Z�o[7�uq��G@�ߪ}��	&��ĽL��טCOe���y�:�ܺA�b�F� �*�Ȑ�xVK�MEL}�:C��g�t/����ܶC�N�hϞ�Z�7�V�r5����p ���*��㮵��(�Ș@�O���R�5����N�i�z��S���Þc���VL��zP,h`�dbaj�BG��MD�Q�+%�ڱ��S��H������k��|寫R�il��B�\��R��p����he)(����K_�����F��\2Fx���`Ųa�:g�����
M(�%����R�R/ܥcYɄqXpx�놪����A�YDZ�b)((�����)�(�2�E�LޔK�[W��w*�ho[���NM�P����0����`Yw'�M���̩�<`��l���eW��<k�PA'�2 �P�����T_[R����ʲ�� F�H.�<#s���<,�GPA�S��Y��ڽ�Vk3�J�#*�G4<2�\Ͼ�ť9�MO�Q��z�g�&t5��I�"�Av������ga���O���5)c�����T�^[(fM�7��;��B��������v�W�]��s4X�����'��o����99t��<���T�:�[��.R���_W�T#�B�e,g�^��#]���q�s�+a�o���ެt6+]�S�����9hW��/��JϿ�J�C���0>�v��vcÿ���s��T���k��^} �Bd�x��u
����V>��ٱ>���Ct������(j�&>WB��z��:�a�"fR[O'�i>�6�4���C7���v.t�W7|�����݋>�Pü!;�g��U�yZ)W��S���Ai�+��Bd#�m6H=}@��71��7c"j�ΟV��.|�O���L��~�F�[�jh�3��ϱ�	��y���L�/��L��T^��;qZ�[N�n$3!�ڋ�M~���BS֖Q"W�:(�t2��S蔭�����ǎ�ࡏ�������0x�Ч��k�^��RG�1�9:?(�9�lJ�em�����/��+W�T̨� ��E��4(hk:�N�Rf��+����{d�G�If<Fm�+t������CI���Q
,�j�~&��T-b�B.X�5qiyy�L��4Mb*��Q�Z��jkeyM�^��UWB�+��${�6���8h����{����8���&�4i�Q
�[�M��	*X�������٬�fT(b�J
��GH��R1g�T1�9���S�+�u��O�~ �D�9��x���E]Rԉ�d�U��Q�hE�d�9�#�5*0vF�LMy�du��~]v��[U��G����T�%4�PS*ӧ��I�C�Z53v)�A`�3&A�qiSKIb6����FC"'�O�\�X����[��C/}�B��������N���W���b����5������_�/Whr|HǏ�z o<N��`Y]	}�]�P��!mr�s��n���@��9a�9OKSE?�=����=��^+�q/��{�(3����k�=��Q+����Y���r�h�cf|�<���ýxϣ�"q�������vD��¼�ܿ���01y?~��1� �� �b�+�X�ʂ�1���9�g�!o+��Yq��OEx�'W�f�����$t�
uC��oP%��\�����8����#s���}T�)d��ح��)��w��b?�f#�Z�l}t�c�ȍ�1��������j!E���A��+�#�
�;����x~n�����!�i��xh���n���x�����Q����/��B_ t�x&T-�ЙG�a�G�
J��	Q&s�(k#�w��^پ!+�1<6����������w�|��ڟvz}c(t5�M����8�l$)�� �h}1�Tm{��
���Z`�B�	�W�e]�kR�����ҋ�P�N�yO�D��l,��C};`ue�?����������	"���]�m���t{~9��    IDAT�I)�6���	Y�cU�M�n��t� N(Wjap��8@Q��P2Z�g	������ʐ���r�A5�I�ќ��텤z	.����03B�(���E+��@u�}�C���Y�K�+VRD�7��ۜ�
/t�X�O�xb�쬯T2�/q�N�!��4Aw }*�IE�O�k �G�s��ڔz(0��5[��M*��B|)��~���j���m}��ާ��ff{�򗾡[n٭���R�~�O�T"�����Z݆���ܬ�
o4��N��J)~xC¼�NL+��(�+��_����8
�M">�T
O�hO���~���c��{� /@п�#5z��?W�nM_�������g\�{��(-����)���Ʀ+@Sr�<���&�#�2��v�����v��:E�yHҏqo�Cś=�͆�{�ӛ#�"�Ϙ���u%잔�?���B�D+��̽��޹�>~/��{���6��H-6�<mPd!b�څBG!�³� 
�ܩj]�,*g�uh�9� ��?7�87�+���(��p���x��#3�ڹ���Sk$�w�>QA7F�'��z��l�!<=��13���z@l�͹?����ݮ���O]�=xP��P(w�+�xr���
9w�&o @r��$��G�����}M�z�HǻA�{��0z�@h�d/�CqaPUa\����b`hH��9�f~�	S��X�<��U��� ��)�!b~�'3��2R2m!���X�st�I���h�W��g�����\w�70^]o��ڂ���@���n( +�(NL�9AU蟰��U	�[k]�X[�Ы�x��;g\t=-�Ci��^$��<�,#W������ǭyc��O��N[�l�����Y�_ͅ�(t�u{�Y����*,kC��s�y��\Z]S&����ZOk����nֹ,�/���Z]�նr�e�}��$쩛�B�����n$�b 0B'1c�]�P�,|64���Y����>l�yxp@�4-(��4�ק�m�� uPsφ�Pd.l�m���Me�	��`-��M�ðG����K���B�$�TL���:9�_^�S��ߓ푄��/ܮ�~�_���R"UQe`L=H$� �6��Ž	�.���S_Y^V��T_�d°ըYY<�3S�����U�z�nM�xOM�?�г�b}����������5�ׯ����z�����_x��r�ٺ�޻491adA����� �˴���ҌD#
���Q(�T���]�B����R���+CW2?����.X��D|(t��{�\�Sq��Q��
�����. �g��{�~}�����f���{�s�{��N{-P�FԹ��m�C87���?S�Q�x�����f�sG[��n���w%�a�r��E�QK��fC������o#��xk_���"�q��y? wCh~��m�����������>�����C(۟5��S�k ��{���S>����9:�k�4�-.n�x�k�:��_�`\�׶?�$����\���9A07�vl�c��g�{����z�}Z\]W2�5�� �UQ%qa˩R3k��0�cz�<t�8�� ݳ6?O:b�Ggz��3
}��nopK��1���2��H��O-�B��`�����F;Ԩ3i,9�K��b��3�+z�k_�ɉ��L�)8
tg�|��@�,�[2�&�\s�q>�,����+�X��o�,n���A�A�4�!�ټp���(�Vt-��Ņ�Y�d��pM8�)}�QϘS�Ht����2�Q��1�detBM��؉���A�����B�l�6��\.ivf��T�$�$�1�6�-�:r��͒��t�p(u�Ž��B��u��m����
��o4�"��"��,k�2Bc43`Lf�l&gт����~��$|�+�cz����e������7���nݭ��_}��ު��@���ڼ5�1Ao��	C�w[��;�b����%ujuU��-����Ջ���1�I"����ſ�'>v���oilh�z:��?�M/|�3u���t�}?6�xx���`gk�Z5��Q�Z��0��i���b>c��J�m^ �sl�f�D�fW8�=@W�`��{��p��d�^�\�q�x>�=/�oV�.��R?�z8�kpNC!G�{dD�~V�����̕I�ЙgJ�P��q���;����a����� �2���#��Z~ώ�	ϭ�4��i�Y�\���\��s#.̩�����U,!�o)�(d��1�ޮ�=W�O��s�ȁ������'�%�5]�2.��c�k2�<���(��y��$_;~.7v�_�~�f�FUq1�UQ��=Z�*���@f�
P�t�~�yO1���ji�j
T{�Dv]�n�P:�[	��7�;G�Ǔ�C��K�e��g2O>�N����~�=v|�]�^�$
���E��B>��O+t��2��d�l��ZƩM��ÔM�9ѧw��J�ZK��2`��ҐNt��@b�P<Ԅ"c�paj�����P�c-���ѽ5d [O�Q��l�hs�EEc6	�8��sv��{����Nlы/��"�o����ܯ;�ۼt�q���w`1� -l�����K*�hn���Ū�#���IdR` �vW�������|�q65��y=z8䪠�{@�I��Gbh�fK�T���n��s٠SS3v<��|Q[�]@nAq�'c���5v���; �F�Z�Z/�(����[0{�ܣl�@(��&R��e�^��`A�+���i�s�kJ�˖C�>�m�e5��T݀����|�y|��^�& ��L^Y��:g�l��U�0"���x/DE��mkLy�Л����|����u_Q�P֮[��8���?�����u�E���@��FU��S�I�\�Ѽ�z#�prVA�/�s�geލ`$����
���a��B��=S�@B6(t��$����s<S��{�/�r��µ��^�;�KQΞߎz�\N�7�K 2�9�{_�ύF��0�����e�\ÿ����aa��E}�+J7�1
�&&���;��r�G��]�U�P9Q@�y�D��o���V���?�7{�1��+���5�{����<��Q1�^��c��3�HS �����c�@���@�9��x�/�1�Kw|.<j�Lp��a�2.ƈ|fn �q��SF�6 ���Í3_���/�y��ό�x ���H���B_\����5P\"�1>w�\��a1��q�tb��/�6�;m�[鼔��\"?�T(w��}��ÿ��7���j5��M�����k��.��\8��X7�0���{e�%��:���1��nաC'͋��:J4�u�����׿�8��*)Q��)ш��p\X��[������AY#�	��7��[����s(M�_X��l`|�N(�����~劗�|��v�E�÷�� 7�<�W?��Rt*�~�NMNn3����	�v<�D���3����CO����������	��K#ZYZS![0�Y�Q�23@s��;ݮQwҔfb��/.��67��n[3���M�@�B���c��RZg}�A�3UD)iy��wxga^������bcۦ0�K�љ����Κ�����/?
�o�%x!tI����m�y���e_�iqeY����.k������oC�#X���54h^��&3'���3����e��E�0D��y�zCC��>s������M�����ֱI�}�V͞<�}��g
}����d�y�4A�Z�����7����C��.y�`��{h�͹��9o7�\Y��ܬ�]Qq=�i�M���5н:W��7pQJb��*�h=��9\���C.ؕ��Ϛa���Z�%R�\���.{�RQ�7$��
��Ǎo�B`O�`���5�?�2�n���;�7ƽ�/F�S~����Fډ�wJs#��R��Q�����2�ߞ�R�t(�g����ϛ}���9��w|�r-��)�����şO�y�(��3n/F�Gx��|�{c>��<��u�!�����3��]v�̼*�V�%���elE�p�
���{d\�k.%���7��znD �aۣ�ϡ�0�m�G a@q���{ʅ�����������m���P5��@C�blb����s�Jgʗ��K��Ζ�2�{g�O*������Yz��o��5K+��c���K��BN�B�w{j-�i�h�fN��@^;wn����ވ�<@�~J�^S��)=��I��_��rB���o� _��v��<�|������u�!�� [��L�V��7t������V	���k-V��i�֍/��ڿ���?Z2�.��)��J��01�Ug�8�<n+�H�Պ%���N,��B�wxF�p��R�1����fq~Q�L�J#�N�ծ+��)��Z��
��}�:95m@�銕(�)�铧B�H:��R^Ǐ��C�U������{^-<)�C�ó���C���7��#/�z��ME
���`FeK�'L]���,պ�!��ToJ�1�S�����s��F"��֛���Ȇ�@b�5c	��m�R�XU �$�
e��3VC:44�B)oh]lK��E
=x-R蟽�}�ǯ|U�����׹��k��A=��^]q�t��	�}l�͑7�1A�Mox��k�c��Պ�P��el6/Q	�{�� �mV���"�7�M(������Ay��	B0t�������z����)��u���#�����滞����5����m�.��7��ρY\��1|^}��l�X�g�Q�cQ��x�e`�#�u}f����Mh�f=��J�q{$�c="�3�^9b	���3��5�X�����<���H�����9x�g� �I��u��k?����E[��6��1-�+�=�����Z����i����}��<�䩎`��L�V��C�J�4s@��`�%����{ꬩ��'��+�V�7C�Ӳ{^��σ�[o�u�]X��(���B�d���ʊ~�u���������?�Q-�VU,���̩�)�Bg�OF����kϿ�����������X[Tm}�<t<�ٓK��z��`.���)�g�_~��t������s���5�\W&�W9�Vc��vm�[��-�dT)d�MŭQ9x�c!�Bo��������M��&+�V�{[6gǵڡ;�[�������p��;E�X��J��e/~�v�:� !W�Tq�Ո#{snq1�bY�,�N<e��Ԓ�q�j��yU��*F(paRu�_P�޲�>�x���ZͪN�<n�cCC#�j�Z�����͒���y�ݶP��W���y;|�@aP'҇x�B����²ż֬7wh���P�`���<���Ȋ��S5`�U8�3��^:���z�S��HN&Lh`tH�XK�݆�3N"BX�<��E�C,c��-n�aC�����L!�������o
}����y��x������!S觎�7b�ѡ�榧�B�ʸ	c�GL�Ľ.֝�#-��7���Kw��B���~����$k�Ƃ�{#B�G}\��$���fA�Mӛ�!������|��|'��Z�vwCPb�4�������Q��������W�@=�X���	��P��9��^Vű�p��,fx����q�=糏=��@D� 7ܠ�{�~=��υ�L�Dt���漶�r]��B��1J�O�)��� +(�bf�>N:䘀�y8�?�Ә��B���� �лGQXG�G0�B������cB�@��Ζ�B�>\bD@��}A�;���>�����\�+R�����d���B����25=m:u�t]��=��v�JS����s�a5!Yx���C����y����;��n:vR}C�Z�6/)E7�t
��^/u�퇯������Z��^7�nu�M����Ԣb�H���*�:]��+�x�^���48"���o?�}�|�]��Rھe\�ڴ���֫~C��EsI�	�C 	<~Q�ez���ɇE��}�B�8�<p.����"L�0�1�h�d�����*fs9�_��W�t�#�s6u�,�{���<s>8%s���оc��7���妊Ó��J�wZ�w�F���k�UU�fLQ:�O[����sv��J����f�-�47��t!�-����M;��O�:�,-���Z�S�P��B`�9qZզCI 4�6��t�J0��Y�

=lSB�27���P��VB�>��t�i�aуK ���\)��� ����qp���ǈ�B15YZ��  ����9�WW�}���o�_ӳ���M�(�.$�\�[���}������WoR![Ԯ��Q�}�^���irlD'�6�7��ny�N -�<��<6�D��=`�.<]����a����֔���x®�s��g➾��?�t��R'QY����r?���������?�zH��f�cƅ<�9Ɓgu�x=��ʓqp<�4��Hf(a?�7�Y0
&����^9���>4���>E�Q�ڔ���b��G�G���\~ots�8o��e�Q��S҈��s�s&18HmqO܃{�Y ͳ�8�y<�2�W'�� ��ȳe�8.���+/GΛa�
�u�V��) �,�uI����/��c2� )�������sa�D]<=���S�9�Žr�n�r-�ml�Q�?�zի_m!����S� �\%�22bLq���r�cJfs����B�J׿g=�R�q�#�o�y� ��'U�	������߀X�o����}`�����m�����S
}���!�B�%DmQ?e������&'��Sҧ��I7�~�ҙ�ƆL����_o��46�W.�@3����%r�,Ґ��"��'�5��	N@t,�fP�fљ7˂�Ń�^�N�h�K͒���B�l�e���A���,46�:-q�[n��:�3ZPx���~�#��?~W�^�����U��c=���Zԛ&�b��,5]�����_ܪC����43���jC'����v�RQ.O��^����O(Q����������j&=zLM�ݶ!�iSi9�x���D$��"O�m ����A��as�斃���L��C�G�;Ke��LF���m��H�-$���R�֤�§�5� N���@�Cg,��� ��=4 YW<�4}`hP�33v�F����P���-S�ܧQ���_��2ɬ��6�ř�:��#z�󟡳�M���C٨C��CG(!�<���D�p���^���+yW⛽�`���� 
!��^rmr�A��a��"���=R_�;�koV��g��3���x���}�ၒ� �ߌ�s���E�1���<��91��[`<l���s��'|)<R�<���ӭ��j9�˹� ��"�!bOcLx��=KOy�8߿��K��^.�!�=&�X�����Mr��'� C�Nt
b�$
�1;vܞ�2��=X�$:xqNc�o�,��YhÍ��)CR��p4��]�L,���&3)�X0��F��#!A��HkƣQ́G3H�a�������j��w����F� �ӣ�Y��S%\���>�y���민������g�07(z#p3�8�6nٺ]sK�V�^oS�Li\�����Љ�q-��^x���zt��o��i�R*?ys蔭���_}˱��[鱉ե�:��:e�Ԣ���B�Ĕ�k��q�M=���i9�'��G�[mv�c{M5���Y�Ի��,&��@�f@M9M�/���Wr�|F������9l��)͂s�W��+
�CT́)���%[d��Z�~m,Z�~�/�T�^z�@ײ���ِ,rB�,��q���Ǭ���;l��֚��+�������O5�%�l=GUW@�� �RU��W���铦��ܱEW���i�"��I7�`Q��SZYoi��R<Ū,]@g&�jJ�N?zO�+���A�X�9S�t1�� DtP�}���l�ը���Q�(}�O�,k 7�fϝwZ��))�x"#YT�c���(Ƴ�Z���ι�Q�Ɉ,�,t��fX�H8	���2#�{����̆�3���9�u �!�����4\N�s��s]���t�?��J���G�����������3R�    IDAT=���G42:j��*�/�	�ҁUn��\�Y��t:�B��˽��Fk�C��y��� ��p�ys�����x�ω�7�c5/>Jx���ɜ�R�3!�@g����}j�=�c�����lw��eԹ�{��v�=�ؽ���!�6�B����۲e�x�6?�w�6�D�u��g��s�a?���|/:�`X06ΏG�r�^Q�	(���.0E�<s��Õ/��;��=<���5�ϖ���_�P�����5��0.��)�b>h�j�\2f�c߳j���￹�W85.�!#�9�&82�3��p�7���ߎ x�T��/��3���� u�0>�����
ȍ�Q"(�sϞ=�I���uP����q,�9�Ƣ��"��6��!mGw���am�~�V���#?Q���{Jn �an�5�/�/�?�aiaE�LN�r�9b)0谾��٬5��}���CG���/���o�A,92^]m�]]��:l=�<�Э��P2�檲�e�[�*��N���)S2��N����I�ܥg����I�	e��}�|��	���<!���v���{�>������֎:���Қ�έVБ,B��L&���b� 3��ir˸�?�lU�W�XkK9=L����v�x�T��I���3w��Z���^B�?z@��۷k������ڒ(8��l[y�@9�k3W�dOoy��EO��t������_[w��}�kvnA��[�0�p���n�B���P1S���>p��!�Ŭ�}%#�i�`
�m��a�xC�Z��u��)��ݰ�c�<F�j�r�^yH�X+��u�������B+X4����D�H�@,�t�"�e$���wcJUc����y��C��Џ�<ZH�c��]�gHW�by@�>i�Ϸ��n[�ZK#�����{��k�����z���4{B���ſ�,]x�.=��ǡ����&l��_��́�O�$u`��\~#&�!w�yoV��Q���Jz� D���� Թ�U#�N��q�*�\��p���e�^�! ls�e���F({�׽G��cxЌ��*���Jj̣\�c9J��a;�E�}��m�7D�Jf�#�QЬ[G_��BIEC��|=���E�����C��]��ܫ��s�xnxќ��a��;��{p�=B倷P����0�������ఈU�e�g��� �a}>��c��؉ �#��x ��9/\\�޽E\"���t�	}�qg,ڈ�����#������C�n \��p�L�t�g�1�}x@�(���Glp�a������!T4�����DҞ��1C-t����ڶc��͎|�q�Z p�j9�R����f�nitb��]�Yo�*=��zM��1���ς�Ji˖�'�B��M�}��#�nu+�FO�ڪ��@����u贀D���*�SZ�;���:���:�����,<��H���3������lL=r>���(���^^�F;ϻ���>�����S-!Axӈ`�:pJ*@�#������gfz�W��-7�urBoy�U�����yįy�kl�������(Ӷ1�7�P��1/<�W��c���ܭc��޲�:�c�մ�?���&����֖�tƎ	U�TK��瑽*��5���V;�yḆ��8�Lc�3���+��y���>S��Q�ݮr��*�ecO�
�G��ܯ����z�V�Ox�E)^�PT2��F�<p���^�eN��5��j�=�n;C >�NS�$
/��M��n'P�6�`b�Q���V�X�F�R�����BO��]���>`�?=3g7�r�r�~�c9u5:�ı�[�j4m����蚏F_��?茳�V_)��SG�4w�����1�=�<d��Ľ��6�I�v�i:��X�X��H��g��y�%������59ƅ���2¹��}��5��2�7����!}��r#��z! �B�À}�7/+
:4�@PUq���\��PQX^�t�%��Bu��wsNE�R߱������εH	��r�
O��0.����zE �]c<>�s�%�3F!sG��H��_l�}�w�9Qƌ�(�I���V^(H�炏�7���\y$��s�`��M�Ƌ��c�����d
MKx^��wμ�<��@(��H@�#��֕FO���
����C�K@�;�##�� �c.,��r�χC����?k�k1/�yx*�#���@34�k�c��OMp`�d�������3ͳ��z��+�=p��WT�5c�v�W�3Z[o�����!��(�@�������r�ޣ��h�8f
�����_C/a@q&7��jWq��I:�$�¸m<1��R�Y5�ft�	�ş��*Y�s�s5����c'��MY�n«�TN��ߣ}��^\Z^P�T� V�F(Ai�Xݪ4aV*Z3�Q���ZU�++���@�^rً�O߸ш+(���
���'Hs�V��t�q �}��6����p���zɬ���;i����.�Um6�Z��y���)/*@��R:������Yx���mZ�F''8���3B��T��fbx4 ����Z}-x3���p�Y��:�ٓ�t�S��׿�պ�s��8���E�Í_Ӄ{�ʳ\S*[��L@�ֈ�t�.N+�骘��]���Q�(��k`�b��pZ�X�JO ��|L�~3\h;K�Y}u]�l��~}41I���fBn�[W���©��]��}��+_��۫{�W�lF��z%�:vtF���S;��~��S��q$;���������?����]x�.�M��ܥW��E�/����f�sC8Y؛r���Ҽv[�!T��)���5Pϡ���P<��߄p]@:��X�Q	f�?�y�^8��+�r!�x8=���˨�Sv�ہ���yݛw �!n��x7����3�)ap^�\�`wc��|�
��!D�z�v�
�NH#�p7�3^��x�������Z��
·�X�x�I�Ox�{���=Gƀ>~�)8�K�ayq����� [|%Ž�S)� <��϶H���}r(4R��b�020&�gݶ�qO��
�������<x�!ee�$�hS��n ���^2cF�{5���'�(��I��F�1r���s���?kK�D\��W��Q@�m8���=���^%a����f�rg��Ƙ1�5��N����Թ�urf�z9��i��cFc�����r�\�Z ���9k�p�LZ�R���"��Ir|�W����U{O-�q�WChw�0�-ip`�&˨_�J�:LV�<&WK��J(��*�Zՙ[���߿R[����܉4#B��`��n�Ls�&�����~}��3!D��\<*�ht��V�)Af�Hf�!7�oT����:-aW58C�B�XҼO���#�Kk*U�O��3�|�_�R�:��pI��&b�e`�P�T�tAK�5�֫�Zԡf��P�XL��YlqX�p�h7KyXW��V�лٔƶL(�I��ba�8~��ֺ��&FP�Y8t���xY����9��9��wL�o��m���M=t��u��ipl\�;w�?��n�m�2�՚�@��7o�������*ro}}���%�Ծ��48ܯ�撒�X�z6v�+^kp`����1�jm�n� �a( 4����Mj�Jݺʦ�z����o��K5P�~��;t�7ꜧ\���Zq�r�Z�Ŕ�WCi�	�1Iƌ� ٪���?����Ǯѿ�t�)����KS��i����y�~��;��8v�?�!��<,z�G]�,��\qz>���ۡ��ߛ��7{�v����#��`�!�\�"������G6�=�Y-��L��T��v���G��y�﹑�1.��Qx���� g|�G�2Gq�bXr���Y����Fٔ!n��	w�w��8���t��ω��lC7���<������H�����)���-��y9��P �˵����d�Z5 �[�t��8�ύ0>gx�|Ǎ=������3GF1N�_H;����S#��M<��
��E
F��	�>���n�F��#�50$87c�~�87��0^^<g�ude�V�J�<��µ݈t��������K-eE;Tr��ˡ���2.�g<�9:5�`(w�e�0�"���2'�IV��;A����Lf��!-�dV�w����|�_o�ɥ�uz���
}�z�M
�G��-�OzQS�yT)�3���/#]z��z��@!�b.�D�j�k�d��;gA�Sp�� ����{v��-�Z��t����q��4�ڳ�X��:�
)C
`��G������)��	��ZX^S�<����F�K��R�QO�
�Ml��.䩢�����M�6Z����W���R?;:4"0 �,\��1��2B\�[&̃�{B@�8a
��lk|dT�|F��r���"�N��|l�)��+.����Z�nj��O�2?�;~t�����ӥ��y���?�;�ݣD��z��2��41R�[��Zm����=��?���9=���v�G��n]:���0D*<��W��O��C�N���%��+�]9�˹��ݒZY H"y��&y0&9`��klcc� �c�Ɉ [�$��S+t���z�������_�?�?�V�Z�^�WU��{�ga�ˎb8zl���`4�{|��(*^���i�L����*����X^t���R�\x1��Q�V��B��nB�{��c3���H���4����4�\�m�3X[:�ZaO�p7� 5��и`��N���Ky�,�
���f���q��,�� 7-n�A~Na�GyľC�74	�pc��H�r���Jotn�
�SxD���Sސ6�.W�^eqF��_��@]ǑA��%��1r��]>���Dx�C�b�s|�a[�����uC �qy|z��.��y�u�$lyyi�H�q����yz��.�J�������y$?�7��|f��Y��w
X)o��Z 䃤�U%U˱�<�~���y]q2�J-�$��
E[��+u��i����1e J@i�#�F��T�շk���	�V��_��L�� ��k��na�_�е�U�^޽Ҟ2�d�p>�`�y�VV�Q��ݣj͑�Lg�xƥ�[�M7݊X�$g�y@���ͨ���D�C�!����S�C�/���K7�m�r��;��$[��C�UJ?��ͪ�\��e�t<#l�܋����M��}�a$��X�r�^��x�I�u<Wgɒ���c��|�=���?�ϾH���l�v�LX�e_\��^$�B��md]�x�9%��z������`�k���c/�p#��(�j����bش�t�L��b��i�|,tl��[�n�n�X�A_�шa��]�;�F.|@��ټ� ���B�#���5"����E#����ԛ5��1�62�B������ٸ��]�2������0n�������1��|���Vm#���6G̉��)\��o�Hȝp�R.��\����8�o?�ZM֡;/���$�qsc��Y�zv�:����z�G���߄{����8㜋�����J�2�V�ᒧ��7��C��^�U4j%#D��h�3�!H��B	�[�@�E�����������W}䓸�C&����cu� VO<��lg��fMl�aH,l�:����m�'Da#�/z,�2�yM�abu�=���ٓ���6�7͹�.�'�%e.����w
��k��-� s���U̍R��1���H7({�1��X�<���+�+`���Qh��B����1�SV� 	�/b�Ho�|�9^�8�e�>���9?�"�|O�v?�R ��(mFW�uj�g�y%���.�ݲ�����Nb<���0�9xM�K�x��Si����K��e���ҵ�H����0�V�ۖ����1�(;OD4���W�a#��GF*�9��y'_@�ևB�"Ur��4�ymJmp�i�{�O^�����q|}���9��c���Y��$���p���[��c�B4�����$�V��Q�&�g=��Ѓ����r!w�G�t��]��Q���h��!�'{����A\	��y L�:-�`�X��g�v�������^�r+�G��ZȤ����R){��	+��������9���ق���ب����R��Y���du�b���5��f��C?f���4��*Bስ�KeG14<���("�ZF������'�i���$�Ћ��FM�D9OBm���CwY���7�y��P���4=c���c����2հbIc�3�O�ql�j���g�N�A$�����W�R\r�L$�˦�,�������cC��:x��<��QL�n�� &�b��?�C�C=4�NS�֨��8ݢ!W��
,Ο@�^u��k)�
�?�o��u���d�pl~�ӳfQOoڊC��a��#��(��R%e��Jy��A����������\~���q�C�bz�t���HNoG�5��������/�->v�?ᚫo����ٵ+�q����8w�.�q�p#��87�g(�h�/��;h�G��7s����=��f(�(�yy�������z�p��k]9��ܧ�o�	����T��󧀁������A���t�jpn|�sJ���7d�ϱ(����y��s��~X�8#��	��z��K�E���sE�? ��Wy�J{褟.^ �����[Z�V�H�h�ؓ�Bv��.���fȹǘ�/�:�,���w���Q�]� ڂ2�\��E��\q��L�u{#�E���r�R(2B�\C��8#�
�N��%�pp��{<��@Exh��,Q����/Ej��йy_%BT��˝��r�dU4��q�gU�e�W��Z���h������`ȝ|%��C�� �!�~$ʆ���`��������t�r����8�ת�;9t%�ȟ@�eh!B�qa`���
:h�sx�3/�[~��(�.��{p��!!9�0�F�eĕ�w��ҥ��G�IG��xw�}�u
��kM��C��.W	|�s��sC��a.�d"m��X�G1��i�6$�i's�T��湓GնF����-�$�X/U������A�I�Y$3��G�h��9k���1���YB0FwϚ���OL
��J�N���y̡3�N@�b��b�����8h��l����G�P+�����'��Z��e��ҁ���4�DƱ��ø�w��R^|�MH��a�^�P2�׽��DH�\A�TD����vnA(����>������l5mw�G,�a�����ȸ):�m9�R�}���ܧ\�b��;�����H�nF���!~_�����9|�d�1����o�>��kϋ"><���f����7S��za��#��>��O��OC�a�ڶ��q��O�<���>�k�v�UP�V!s�T��r|~}�4��~��f�¢�����]��n�sc���r��;���t��{V9�ꑝ7@���*e�x����r�"�i��]���`xV�Y��5������9>I�*�j��HĮ�ת��@���g��OҤ�C�s�k���G� ��2e!/V���2���z�O� �����Tp��l�t��Q��j%�~��e��GA���)�y,�@�Kn�ƒ�D�U�>�Gs�"ǃ`�Rqh��%��C�ºP��*��`�$D���t�yE��R���y&�$E����S�E�*.:��V^Ǖ���x��]?�� �06f�U�/��Xl��hɖek�@�v����ia���FWN)@��������VJ�O@g���5�GGƍX���7���Aup!��)�EI�z�����ҋ�Gǫ����P�H5��`���b	M��l�A[�P&���CXX<j!���C63f5Ձ^��+w�E9Mn���35IU&2�]n(��[~��Q�'���d�m��D�Z���v�q&����;�G���f�8���z��(��,<D�%,��:�څ���&3`�=��9�肿r.�������O� �5��'}jb�<������ab|�"^#�Z�>�?�E;�1��B��5P�o��c���'���    IDAT���*ֺ	�� ���U(�8z �T�m*�D��P��|n�x�F��F�Y]<n5��X��͞�_U������q��x��_�]���g�����X���pC	]� ��B41���ҙ02�&���!X_Ca�(�!`�T��w܃r+���k��z6Z�	�")�Qt�ģ���_���ᓟ�<>�_���4�;�4*�8���8��mNceei��Y�Q��.�=Z���*������iʐ4�������$��yפ"7<�`N���X��dՠ�������AGb�Ե�˳��! ��e������Ǔ���3|	�酩F���wM���!ο�w�m5/�'�A�%h 7@ȿ�X���xu][.�f�S7���N������w�_+L=4�1��6��z��N�t���6����zU��xE\������{�6���P���q?�A'Vk��q�u9���+}@�2�N�>4W�� �y�N�]�rV�p�*�Z��!����?V�l���~��"Ez.8_��Ǭ����ly	4?6o�3)'�C�j"aZ��C�޳���>�=+���vR4f|<�9�;r�G@��N@G<e:�}J�����/�.U����� ���F��M@7�� t�,��*�c��	��P� N;��l�d�
{��M���
).�"
"� ���&v����Q<Fϐ�N�Q�#Y#Kg��v��䘝�0����!���mTv�Bd	�en��_�������7�)?��N�&[Gf�m�������b�z��FF�vw?�w����"�Qx� J͊[R��A�1� �LՐ3��&gN:%Y��o4P�=���Y��P�h�B���؄-�����\#�86�nF1�C8�B���{��V\x����h��D:���On��
p���Y�a��!�b(;��� �n�hӣ�U�ؼmw�s�:w+B�.�W\k\�\=ɛ`u%�H<�c����C7���[\�J�DȌ����bxj+�� �:04:�V5�J��Gߍ����Ǐ �Hu{��ý=�P$�PxH��ʠ�"MY-F@��}�e�g?�^|�3W�ӟ�
&�&�s����<���c(M�j�%G���qz�ʃ���5�p�y~�K���)�\{�����u�~ t�&sz,���9לj���A�5p�!�±:.�/���0�2�Y�=/�?=U^���yS
i�o��͚c��	,
e��_�'ߓ��Q�6}��US.��c��J�qV���䵹�`�_�3�����"ּ�DOv��v�4��;��+<;���7#�os��;�NA�F@��9�[��|�Q%�y��S�ԱNDDΙ�Wiv��u�k��0x��w�^��4t�_�Ĺ�MF�"*��T��_�N9\�
]{�f���Je�p��8^��~)oM�n8;d@���G\EŸ3����լ��wރv;�Z�������9:Y��� ݽ� �:Y�O�S�C��_�ˣE�͍Vl��h��5Ѭ�w0scQ��hR:�tz�X��^A{ϼO֫[��>	j��������!v�<�f3)lߴ!�P)/bl$�J�8��[s��A*6b�8=�E�@3h���6>{��p&=d�I�N����$^���]��w>d���qg���~�s]=f���ب5ya?o�lC�z���7ⶻ���vT� Z�$�2<*�1��Ԅ��p:eZ��FA�7؝�R5O{jf� �]ی�u��)��C![w�4��N�n(=���it�z�2��E���/}�ٸ����Ѱ�~��z����W�����|��#�-�ʹD��nJj��7��矍��byq����|���@V�N`jz�ھ�HD4��,
�yd3�`nlu�����_F'Ŧg!5<�|�I�&�MΠ�`-_��-g��N&�V���'o�򁇰p�Qt�u����}x���f|d�����7��"���&�`����h
_��{�w�
��F���#��������K��0�( l�s& p#�%����e8b�#�z�
5�	�_�'_����A�%㖿�P&0�w�~���)�Q���(w�MU�)7R��),���胹eG�W^������B%U9v�0h���@�`8�%�O��q,��8uL���)��E���=�w-�d}��QM�<Q���� P ��>�ؔץV�rּ&��Ivtw�?�k����L2�V���/6��3#E(�����"��<���wd$h{՚��w�e�(
�9��d�p�Ůw^����������n���ϫ���%���ַ�s�{-b��2>-;вUQ����>C��<=t��M�眡84du��>��4|�K_���:�'�̑ Q�����Lإ�~��P��M'�J%P�>C(�53�����_�����h����k�r����b��>HGx��{� 7�>�*�`�u�Y��J�Ȥ☛��W��Q�!�o����{�E�.F�k���ajt���`uє�ȵظ�>T���n]Լ��ُ��/~	��y����i�����]z� ���6���&�K�a:7�J����VkA\�͛���eD����Xv�IY蝞�1
��@w�s#�z�rAvzhV�F�s�����63!k$�5bq��$��G���nC� ���ћ^��>{7�����ׁV���+E$G���~��k�%'����Z%o鑏�o��OC���=�r�D{����k����)�Y�nv��ΐ;�S� ��2J�*�m31"	D��Ǉ�DM�@�%Og,�Q'c�㘻��kȄj��_�����ǵ�M&����C�Xc��n^8���,Z���4"Q��t�D�k������>����_�	��0N��F���ؾe�f'f��v�J��'��-2W׭r�im�"�ɫQ'/�J���B�bsCb�H�g�g�=q��Oc�����b�s�
���鋔��"Q���A����Ks��)��͛�KLn^7�0�>C���2<ˍ� ��h�50:B�<���e8����P<��X9b�[��O	��'�L�'�S%zJOp>M�>����i�q\<S{������}�F�O� ��	|�}R�<h���ދ�h��V���dPh͸P��"!�ᒃE��S�S)K]�,w�������С�Η>gy�bq�����#��ce���a��x����oJO������S���q���̓��s��� �"C�º�`C&��Q)���O�K�z@��B2��2]��A���t�?�vyd�l:�P��~��8Z�~Wz���O=t���YP'��uEӋu�u�P6q��d"�P�C���^�F�X��m��p��Q�s��j�W�R��m���N�N��Ұ\����f���]��l�R���|9F�G13�:!�A�4;�!��/�Neq�Ӟb1�����q��N�C+��a��z��H�nB;C�M�	�F]�~����������u{�*Uc���Ǣf�Rnw��!��f����=��{��V���3q���E���W�czj�}p�u���M����h�0��4$)�V����{���vcm��Bn�RO}��ȭ-�O��۰0إ��|7A�d�Ͻ���Xn�L���b�Qct�q�j�:A���b��3��fM� �2��=�=wބ���!�Nq��x�z��E�@|dk�ť!3>�Dj�����7��F�z?>z���u?�Pf������&l�C:�i�o����m$(yw\K"������ɔmb����'�q�RH�����67F�뵉*GI��F"A����_��|�;�����8y�
g�|���*|=�S�6v<���u3���SF��M��@���
W/l�h8���p��|��A@:��aȞ�j�Q��	�
G+t�<=G��RF�t���4�v��F�ב�!T*%#eQ+�F�Ͳ��.�̚�p����>0��=`n�fPO��'�<p,~ͣ{�P1��$]�H��S<��4E��;�
ϡ��C��l��6N1]�%�Kz�|_5��j��E�\����}����9J�DϚWU*���*50��Oa�y�ܜ��KY<���v��	��US�[X��رT����`S������lͮ�t3TL%/���L\&Db {��L�m��S�C����G��[�^|���mb�q�wzxC��uTs)_�~c�Vɣ�f�2�2�z^�nc���Z�h5s����1�S������XI*<���7�pQ��9t;ƒ���?\t&��`�Z�5��͠d5��\����[m#�47�յ5�ڹ�V��4�����;���%�)��A�G���[����*H,r�y�:����z�����F��@�ga��Ih�d��~�TҢ�j�k���k��q�߽���ݸ�K�����x�kd�[n��|���H��^|���>U+k���'o�M\��q��<r��XZ]���]�X���~��8�o�q)Z��F�h��ѣ�r��V��$��E��0�"ec���:�0"�ʵ��&�RA�+�x��G��Cm����'���y����@le�����fؤ��D��jU�Nf���}W~�J|㺛0��eO�����؃�b��s���ȭ�Z���#���z�A�7J�r�b�>y7ƫ�K���3���Xǖ��9�Io��%h��U��h���t%���X!~�]P���˘�+� �ߕ�+��qT^%�P�^9]��T�� �g�r0n�����ש�l�rI`��x��3^?�A#��C�  �s��wd9���kU���}��*����qs�f�9'8Ѡ�|sS�񾰰�_��_�]w�eF��ϼܔ���!�1m�<�t��e|���4����V�hQ���M��.o�W~\������pEB8�|_����`>\޾3�ܩT���4H��e������w�}���H!��l�1H��/�\{��ok*������O�5�t#�}��n��6l۾�vۺ�����Ë��̯�M}��v�%��#H��0��0��$��.�?R쏼����ˣ��[���H���B�~��>��Z�2���!k�e�X��� =�InWQ������^������	�w÷139b^z���zm�n1~�cȦkݲ���0Z����?�sqq�V�}�P?�"\�sp�Sγ�5d>��
�����K���l6���M7�/z1&f��ZپC���o�J��^8�b������
a�Cg�6�>���t��i�0�^�).���9�-�����c�)PӔ�6�I;�@��"Ca���6�)�=��C<�m��D�ě�����Q��?�.�0:w:b�1�KE-4+k��#�!�blx+�Tk%ē�MO`����IU�PyB
u�@f�c�H����6T��c�!bqĳcƳFtk���@s���t�����ID0>3��䧸�_�E�B�Bvr3���B	��9�j��m������������k��H0��?�R���܁�����_}��^� �{n��x��\ޫ��k��k�&V,;���q.����;[�`���e9}kzH��|�(�)m�V����8^���1�{���ƾ�<� ]5����j��MZ�m2*�|���1��!��^���3�e��z�^��A��a��0OO�@,<6��ҥ��ss\
Ws�����g?�3��ca�w�`l۾�ِ=����,J±�/��o�w�w���4gߩ�Z�қ�3��{!v��W�qGT��LU0-}�ע+���5��i_ss���p�ClwF,�Z�zN5O�+�)�g8�4J���k�:�j������ .-~�������\���x 2r�ٶ�]�h���B�]Y]Ŧ-[LXfߡ�8pฅ�	�L]����}|�������Zr�t6j��N@F��f��R������G�ޛ�^d�?Ρ�O��� �?ђ�=��dm����W,!�ct4�׾����睋�p��>��=c�0��*��2�5+y�gJ��U��ι�he��^�gi���<��qj����=�̡��%/D�V�E�6�-&������]w��!�I�8~�*������D"_��4���-](#3���D��]�Nǲd�sE����&����k�;=4JeT+�SSV�֦�
a��<¾pB$H�� �Ѱ1D#�����E�i��Goy=���D�J���Qo5q�`�\�R��;�9`=܃�4�u��gz�^�z��3��"�r�ض}睳��c^*7�����s�!�����T���+ijd����+����#� �C�b�7ahd�1~�U������-�97��0��pC�ø��[�� N E�F����qk�h�_j�J8��������������� �h�<�}�݇�ݍ���ⅿ�Kط�	�kzm�J�[�8=��sM|�,-�*+�nP�M*��[��_Lcn���ˎ�I���`UB�2/y7��kSW�\��<��.$���N�[�a<�E|���y����2&t��w�v�^��8/��1�M;�.�[�����!�]�^���y?������|��-6Hr�r�2*�s��sA���g �LXİZ���$�/-���x��x=����b����K�xm��2 y�SJs����J����pye'�#��{�rJ1����p�����\?��K��9��W����?�*G�E�����_��5%i�5$��o�_6����#��?�`[�����M�ࢧ�?�!�>���-��jw6t<lO5r�+[$�9���:=�^<a�)I��o�?���~�]Ǌ��nx�,=t�[�N�g*GN�3��n����	��<d����i�,��ǖ-Y��ͯ�3���$a�x������F&�D���J�:^�Nk&�D�d0�B�.�f�!lz&l���q��b?s�4.@Ww>�׽�u��_��}{�������ãXXZB�M�~�ʥئ�u�dUr��N-`���1�To�g�����IM��l#�����m�F�f�x�����+[sD��I@giN��T<���)x,+a� ��|@�M��� [�v�܄t���H%�����ۯy����"�b1=;�}Gcd�������%�㣦��c���Cx����I?��V;���&ǳ��ģ(��0�ɢR���4Y�W�0Ɔ^�r�����M8����&�7#g���廇ǧq�O�@85�~0cVv�]��Ho��������[f�p�����Ǐo����B!����U�\!��׋X�޳H(���2�ݽ�����}���1��3�z�n;x?�ڵ�����{����/�1�����ZB+n4\G�¹q�y�\oI���!I�D�d��Ir��y�7�<�~�;�:�W�Y�����k"hr3U�φ��1q��������<}~���M\�w���[y~z�|q��I�%9[�����IΧɎr>8?�?�5�{"�9`s� S�-�eи��P���F�Pl�۾p����Ӱ�s��Gܻ��Cg���slg�w���7o�b�����x��T�M���J�\��J�2���D���z�"�1J)ֿx@�8�^�\�^觼��9�u�\C2DźW�%y���(�V�Q��rӻ9n05����Xy	�"�^��3�Mgl-��
�Ų@
ˌ�M������X�M�=�J�{�cf�G��N�n5��;=�S>���r��_����E�u/���[���ekYDBQ�׊Vk���]��\��ɒ����çϲ{(�E�'��j�cnv�~�3Q��q�O�E��-E�.C���~�L���Ix����~�Mձx݂cܗ\�:O�B1��
�6d𒗾_��7-����MV����Z��:8�̳0<>��ܺ-�F��Z��H"�X:�ɹ���'J�����u�F�Rܰ C
�JN�K�|Q�=@��v�E{H-�GV�����q���C�FBֻ�Rv=��B*��������l���m��EϷJ�=�>�b��W��7���}���7��K"94���f睳���#�a�^���Ǚ+\���(#��>    IDAT����J(����lQh��K������Vӳ[05�وp�U��Hē�2�ѭ�cr�td���f�����o{>����]-��sva5���<�Z��-�w���5O� ��R��p,��������H'����������g>��|��/~�HϺ��XZ8��{���ho��7��;o��cHUb+�1p"hs���j{�sg��ֳ���=�������dܠ�W~��� �Z�E\�4Nr܀Ur4��9��x)��cs<֞���}���X5�򤌃��`�)
@&�]�ay��'���9Ny��F^�c�K":F(�>�μ9����3bMk<
Gs�֣�O!�d�h\|�yL�>=i�+	p�W.������N���Έ C����]={�tw�>�t�c��Y�����.��bK��:��|s.�n,̓3���G����(ͫ�;���-��)9*��b�d�W� ��<J��^s=����X��������7�uNIb���T���)F�Z�w��r����彑��y��ß�w&�u)��I��=35�mo�!�p��N@���šc'P*�0�����9ˌ��v�?Y��d�g5���>�9�����9�{V��W~�[�=�����	��͞F�V�p6m�������ћa��fbiR���L
}��������s��mK�N'�@�u�	\-�!m7�l�Q��[��Ǻg��ۈ�	ڮ�c�J�±M����xN����x�X���Uˡ�&GS	c�S�f}y��A�`Ӷ����8���"
��L���׼�)Q��a{m�|�����ex����iүd�V�(��!�۴����დ[Y���k���:g=�{�eOӀ���V�Hg�>�׿�%����#��ٗ?�ο2�+>�|�?�U��F'��Iصz�u[��U���(�ȷ��+ȯ��x����{E4F82�@�욲\*����^��W`q9�#�����2>���USڣ���D��.u})�Q�-a4�_���#��'?�76�5�h�P�s��BT�]�w����@�Z������#�(��[]��>z��cW�#�>y��L���s�D!�����G4�����e&������Fp���t��hd�h�"P��J�x�yi�I��y���)N�7s�yΫ�Z�!
d]�թ���_�|m0'���ğ���
�˃w%U.�.Ä�T�h51�(�������A/��^�"��A�r�N�@�腓��ۜ(r!��S�w�pQ~�6"e�����@��9t
�����mIi��(�g	��?�4Y�����PXǉ�ƂgZiii�>/e?��)*���~��h����z����"�2�4�2b�\�yۚ1�9ʹ�=]#��օ���""K�A��z��]�TMa�O��%��h��-��k�1u�c@ 	S\�C
��~�F�YaOF��0�?X�F-���"V�H%��uǗ�O�W�E?��.!B��/�d���N/=�F0�B�������_�����^S�t��Wo`4�a'O�ry�+M��o�b���[n��$[i���T�15��a#z�?�Q		ud�yA�PcZ�lb���n�:\��@�k����l�̒c�=��G��(2�P�ٽ��Ƈ23<�a��l��y��1D�I�9�0�M���J�N����4�d\��ȎO�����x���Z�$�p�q�T�B�ϩMnc�ѓ�Xr$R��^C)�C4�ܑ�'�����]���4���g^r83>�S)̳�㢳v�Mox�Uԫ%�;x -��s/|*��a��u�E;Gf|�r��ֹq��������e�-���������'���-���EHRk؃�	�̲����XYYá#��q�nԛm�╿���w�����÷~x��I6Yڦ�C��ࢋ��W��=��~r��n�s��(Z���>�b��-[wb~qC#C��=������/��\�����[7܀k��I��/��-?�톇�v�B�]�c�ݍh���.}�#܄xm�ZyCYL�6��ʣ���eҤ�ʖ<οu;/D�7<�Ε��g��{P�E9`y��>�Eώ�b�\�偮\�f⊜<����
��3����@$�Q��s�x������5�y�1 Pn��c��I��yz�Y�5
��P�+�S�Y��V���1hp�]�]���A½ǁ�3�e��&�7�uJ����̌�=�E��1�9F���sL�[d2C����Zn�(I�T�=�N�1����k�p�b�ʕ�����h�����(��y�K~N�t�)3J�0���H����}�OgT�6T����xO�փ��Α��<h�|Vx/�O�x�\�2`��X�>���������kL���wb~a�+��t7��=�N0�P4�~4�@2k���SNX�����|���5^U�Fbu��n;�9	�Eg�3��!��5�.;.nv���a��l����+�"h34+8�a��j���i=�QH��^�Tj�?v6�6pg�s˫Z?r*�9ˬgF�3�a=���X�4�N���Z'8*A5Z�u�a?�&��,�@��<��wo:�4S��/9�^�L5bs�Q�Z:n�Ԣat~O�+��lT8�t��}�=P6/��6�F����+�i;�N��e3zl\���	+�����A���N��)WN�i睍�|���k��������On�mwއ-;�ž#�f��sox�e�Ic<F�k����6�k�+���h����Ӯ"�p�)7��y�O��@��ۊ��i�s��dabr�^��~p��8}���82D���=�g\�4<��M���޽���X���vl�v&��!x��/ R���.��i�y��7b$��?p���q�羈����M�T\E��ǁ'�����=07%�M��`ܮA�en,
r�W�<ܶ�A���VuD����ڴOzI��9���ǵ�E�o�?;��]����67m���N@QZen|_F�lKm��3$��"E��
�+l������� �p�n �ʯ8NJ9�yu�´\g�*��sDT����Ǳ)�����~E/���,ǥ��As�9��<㌝v���/�*�����4Ǥ�	���]E��@9&44�?O/��!C�g��(R��?���9FUb���8��n����}�g�:�<E{y �����urr^\���(���D�vWٜ֊�娦��q�.[����Ӯ�
�d�e�_\��j˹������'A�̩��[���7>4_h��ލD���z1W��	��^�D�J�����I�0����h������0̍t��s�@7��/�sMLx~���GB}�������"Ïz}z��Ō�JD�y�]I8
��^C�$�O�@"E�V���v �����b���G��Em�Ds۶��|'S�1ی:ݾ1�i噐Lߕ��ܫR�<l���xa�����E=��_�RX��m�4��.=�k�;]��Э{[����� �H�ڨU+H��8k���bz4��;�v˚�����qǝ��.��2Sؼc'�VPc��U�p4��u@h�^.#�(�WG2��(��6�p��ɬ��ֶ�k���sg�O(6�W�@!W Ba�3�hV��cj�n���0�5�����5����X�R�#C�z4Ø��҉���[�Z����f���M���xe���,�����q�W��V���>�g&�ӟބ@�ë��+���j��C�F��s�_dŁ�0�:il�P��_�$?Ǎ��(�D5�!c��n��X�!���<)��Mǔ'�U�17u��	�dTXdŗ��X��{Z�<֓��PxW�*@W�����	qц�ݻ���h��x��!�ϱ���x�`TN�3�5���'�Tޱ��(	����9/��Q^$�#���x<�P����
�ø�DE4�-u*d�'���3�1h�=�����}�L���y�����cSJ��c�D�u����ľ������N>�,q<�&<����RN������'�9Ǉ��{j�v����ΐ��q�I|�W=tz?������߽�����^{剒��z/�5;�Z�D)_pGg��Յ��J���ų�}~����߂tv�^�^�N�tO�|�qζBj�����ZN#Ɋ�h_].$p�D��e�~�vˀ�i�^�ら�D�t	N�$�!����m��p���@��Ǐn��pM��"�������-�Je#o�n݊A>����I�v<�R��5ԙ�c�d�<e���BӃ�"L/�m�1���mr�Ѭ�Q-�#�b��9�����ı��l��1�`��}�x�!c��c{�����yj^�`�KF]��!��1��O�Pm��q�S���J�r	�j	�d�r�JcɌ�R�����լ���<���09���ʊ��ܧ��Iی*nҼ'�X�fӄf��ch��HgFl��H��Y�	,-�[��T6�7	����Y�}<��g3�D�y�J��b��z�a�t�N?�jC�,�k��*
�گ|�^s=n���HD¸��p߽w����&b��a���(�;�Qʋ���k+�,@�����e��J�"�#�T�����;�N�6� =�!0s!m��Цi�_�L`�\��<����څQ��*T+�A�Q������s��.�?e��:lc�B�߰�s!��yOn����;c����"F�� �f7���ƒ�'y�k�?y݌v�3"�� 0����ܹ��I��ǖ1���s��OP�������A��1w*��]�#N攝���E�J�A�<[C��2�Dp����<�kJio�~#qE�7�*1��x��t�י��9��קT�ຳ��3�sdc�}J��)Ne~���M�0�ș���ɱ�~A=� �r�8�	�F3��3N�)�w�J��|��].�^�@�`�z�!�tn�v��RQ�\Z�ٻw���;ز8~��C�Ԅ��u��tC������@����ΐ�m����9�ޖkg���X��ud�v�e�b�ayF����}����z^��J<�����;�ׇ��[����a*�˧�B��^b��$���i�_g'�D�p��%}˟�=F�0q^��<s-��痦[��T�-�@�ը�Z�!s!w����9浕Ut���Ѹ�DГ�.z�҉���m!� �azl�$v9w&Y*ddj�	T;]�=v����Ma����U�kc��6��M��Q�W��p|�	���Ex����9�����0Jf�_��} 34�f���Ms8<���ci�bI�D��--�@8Է��^����D��(M�p�T
�U����C@/�x��#k�o�}\��H�8��y対Ǐ���a���/��A��҃^�`x|p��(�d�?�߷�l�����A?�H@W�U^��Kb��[vac���f+��^�4�h37D������?;�u�i:̛�:��U��?Ǡ�+�)��ǧ�kyo���N&�ɐ
4��U���BW��c���]ˋ�\�iQ!`�����F��3X\HZ�d�Ô��wynΕk��矄E�8��謆�="��0:�[v�v5V��� ���`4D���t�/����62��;ﻈ�"�ɳ��4.����ɠ.cM�4e�g5N�Z��Ω����9#R���tI�f��WsH%G,�i�����9�ˡ�6 ��C=�S
�o_��������6{�@�ٵ.{��f(^Di=g��=�=z�=����K�g�*X� ��|����I}v�Sp��0Ӡ���!��9���;��X�N���'��E[��o&��=��Ҍt�M�Qɯ"��`ۦi\u���1'_��V|�S_F�ME"#�u�L�kvP-�l�'9��>�l�M��c{ט�z�ф`M��XjB�	�]pD?��1���S�#����.Zuz�x��(-jz$n9�~�mz:r�tE;ˣ��cTv�G�����'��c�D�����̖�q|��~<�J�E,D��C��C4��Ms��H$�(����lձ�p��YLOc��	x�Z��mt4Q��M����Qo�e#�P�P!�O��ѓ���{121���1�W�N�$�������љ^i�\s�d2�6��D�Y�Vꨖۘ��A��1��@��ё ��N�<����8{�N��]8>��:~�^�n�՛�U)7\�Zw]�h���6xy��Kjs��*�Yya��)y�px�Muك�T�X�$`U�]
o�h˺�I��R�j�����X�)��>+/O�L�\IQ� 8)Ԭ�O��U�{9AgЫ��(���<��y4����\��������6: wZ0���L��T�/��@�)3+T�#p�[aq��<��lԣ�@��X�y��]����w)��o<�~�{��p�(�"0�8���#4>�m�+��7�RY�`$�s��Ґ��x�ϵI���$��3�����y}ay�Hq��.�.@7�F���I�`�;�{4��:��u[���o��d\p��	�+���������f3�C�Y.�KgȽW7&���0�:���E/���o6E�v/�n/�n�eZΊ6"���ϭ��M�0s�	�N�����/��U�:+ۤ��V^Ǳ�p`ȝA�H��@��g_~	~����j	����x�CV�Fb\�l��m�ԛ&�s�潒@ǐz~�d,}���b)$�CX�Jۂ	Z�Ǽ��刬'-{����{�Z�X�X@81@wd&G�akYz� �*3c��qڌ\x���E1:HD�z�ݨ� �I�3ع�Lx�-�^m!5>��b�F�@��8f&'164�cǗP�xhv�,u"��n�3��,-���sתe�>0mB;��&�aC����Ǣq�ҹ��0#���ߪ�E0�
��%$ba�{J��y��d"Q�a0j��@7E��Pf�O,ct$�P���C2����<�J�C)Lf3S�w}��
^�ꗠQ+�R	����&]��70�	�s�p%00�ȗ4xMγ&��V��|7�g^��"77�S17+�`ޗ��u�x�(��[�]�y�@�He���x~O�)�7X�67��m����`�@Ӻ�U��+?+ ��s��ynI��Z%23
)K�@՞snu?X(>��B�������j�ȊR2c���۾#cX��1���I��`p���I�q)�%�g�}PA^��2��9�2~4����
�#><������/����`�Z��*�Ces�*�lPZ����j��up>U�?��q<<�I�����Xlcl*W+��ۚ��ޅ���6<��u,�䱸���}����YqD@��6p?r��w�mN9@�k����?���./�z�@8�A�P���a���X8q�H�<�p�m�(��p]��B$�2��H����8ˉ^�-z�ldQ�&��3�s<�ڸ�J2���An�RS�<h<EkL�<���~��x8�h�2�$���g��:��T^K�$i�x�*:ͦ��Q�9���\�a�Ă�omٴ��r�)��,Gf Y���[��6��JAhd8Pp�s�]_�D�6��N�Fu�]!�?8����ܗ�D�uLE.b�p�`CrM*IQA�17;��|��ce�(���|q�'�\x�E6��?/�"��W��\��O��<�f�01��4E�����	Z�7Q2hbtF����;�XF��p^=���ZmW��u�� �h��7��0����m��ŋ��Kرy3�N�[Z��������������,��q��V��+���&��������K���8��8����z�S�o���P-l�v^%G��$;��ԁ�S���-����@��Y��Z��`�l��+77i����&��(7C_ʯ�sb�S�C�v�Ք3��1:#��pWG���ug�l0�N�����XDZS���;��T��3�.[boK�D�v2*���Wy�@������	�	}�H�F���~��%0��T�@e:~��"�����[��J§@�c��Z,���\��<`]�"����^Ɠ@Y�γ<X�Gea���j��F�w�_�n�3~��U��P�    IDAT_�S�1�S�s)�s�kUjH�^��߹Ɣ�44��a��Ȉ�����e����7��$�� ��G�03��Z{�F�\C8�@��%��l�b��v���$�Iz�$�@�ҧڧ�ru�wi���W_��b�V/��+ru�q�H�r5�A+	cٚ�la��_1�F�D�QiT�'8sڦ�B����!'��a��I�c��yݬe���%a�4c��őQo�z:C�$�����Q��`u�lOJMx��B�k�Lk8�quHd��v�ځ+(�*������0;��'����A�A"\Xu�cc	S��ȅ�̀�աl�~�@��s�I�k�X��ʗ�:���m� ֖��R�h%��p����� 8@ǿ?X�C�><��}:��ηcn:�Օ"�
2��Ϯ�����g���c�|���W��ZBzt�V;�؁�L�V��ٙVh�l������ay��2����\��k�C�矆�~Yը�a?22d�@�xM�VW�}^��"���	e��������؁�����L"=4��@fd�P�r�@ّ�U30Bѩ�h4p��Y,ޏ`��raoy��Q*�l�!0�4���6c�T>Z�@O�6~�[�ꌹ)s�Rm5��	$|_^�͗_�r*�6`���8=v3���6�a�J�.��¨4$�*�2O����:7�2*X�(u\�S�o�k���������X����Y`) �y��+5�sX������+�+'+���(�  ��'O_Q04ry�v�L���=+��xΖ����(D��h��z��LU��MM�]�`�A��d�2�8ni��3�k�{�0�B�ڏ�>ӽ�1����WD�ȃ)��ׇT!b�ɜ�������� �CC��}:3d�^k�q��<*�JZT���~���������;wn�%quPBg����~���?�ׯ(V�算��"�U(�B���R��HP��iD��H� �P˼\��]�Gϗ1S�q��}@��o���
i>Y����9�P�'��&�L��_��+�ny)z�ѐ�{7U��GG�Dj1�G"�@�тG�z�^��WA�D��fL�Mcimňjg��/x�0;1�J����$j�����R1�ˎ\4xh܄#�!W��㦭B�<[�~C�4������%��T�R�,���K�h�+���d8�l�ߡ�N��� ��6z�v�܌���]�D�xྻP���a�Zv�w��щM8�����p
��Óؾ�,3�Z^��*����`}���wY7�J��3w����Pr��H8d^6�L,@�sK�n��%��w��ĢX<v�����w�e��T��XZ8�d"a-k������t�y��{�ŭ�݇��4&��c����!6�A?�C�Z�\{�\A��רᴙI������x�zן���}6'��X[l]��`�[?��=��+����s�tej.$�75>K<�_Ոu|���8�5)�̶�j��at��xn�
�+�gJ�''Y3ꚴ�;4��o�����*ϩ��$j�=E�!8�@���'�cKmO ����p�}2��#��6��)#����#<�$M����?ߓA�k����|v��%��ny}֐�G����Jp����[F� X�9v�B΋R?��v��眿K�)����9ߊ�(7�5�c�ZyO�����C�
�sli��S����)�����{}^ڠ�"�WZ��f/�p���G����k�ei����-�>3��zO�=�R�C$���N�%�6Ӿ��G��~�f���:���␇������ P�`�ժ�7���2�p(f&5��z�Y����^0�kA��z�@��
�j���%����P|>W����\����O<�Tk!�"��w@0g��Z��<�v�<5k���I�%_,+�CW�TP���-G�f^�eaJ�����m�AO "~�5,p!j�h�귝A�׶Z��̰�4Y��m��naj|g���*�Jz���3�R\Бby`6�K�u��S�&oJe���f�f�1I���БU4��y�H�X�x�����<:k�5&n����an��U�1�C����D�<��V�ѩU�����Iĭ���@(L��L<�kl2����G�w�M��]�v�,�#�<d��ҭ�M��k��G�����R��dr��P�x�r�do[V	������Sw,w}f�m��M��Qt��w귭�.�b���*�Z���[E*D*������s�f���ż	e��p�wa���1^yWiPu�at{�ˈ��Xg��Ӱ�G0A:����_oëֱ}f��Et�X[=���篰o��f8Q���dn�4������qT�i�t,]W��w�K��
�&Gc�s�ߝԪ+ˊ'\N��޷�_��(Λ�sS*9mw�g9&�y����x�7���_�B���8�Aje2�xl�8�k��;��kS����� �ʀ������ѣV^��Xغ^�?v ���v����3�{�����%�*&�B�/�G������wQ�����?�'�),o��/6���&s*�1��օΥk%+�Phj����c�ҵ�p�8�|i��9�4���"-^]�6�&yE$�w�0��8E,�5c͑X����(R��ս���t_�<��Ѣ$�����)H�o��*�`�}n�V�M�ٳ�J�X�y�|�,����8�q����OC��~?[�z�����~��v�}F�՚��z��{���4�F
}7+����l!�/��=�ᡇ�]����K�|��/��o~Y$��H�3��56:a�-�e���Z�E��j*�10%�s�lݲ�B�6�r�l7�J����s�2�N0 �?u��$0v�T�*��%}Z��m���B�v�?6��'��Fլ��o�����{@YVV����T���s�i�D@���b�qt#�g0T�Y1������H���r�u�n���=�ٷN7�3����굾�V�[u��s�y���{�g?�٭E��١��H�#}����<����@R���R}��p�"�M���G��T����a�#��,-]h��7M��GR�^�˩OCϩΛi�q�����y���j�ШOZ:Q��mգ��5gy��5�������>�=���7���m�i����%˗����_]�E^�����;��Ѫu�,��Y���L猾�C#c���m���J"cu�tXD�IUԫ!��N�.\�|8kXub�2V�y�Su�O�؂��K'mlxH^e�Olx���tڂ��l�cZ)�	H�4<X�E��m߾C=��J�mɂ�R���l�d;�%QSE�
٢MO��x��6�s��m��Ġ��ԓmr��蜈�ˏ�y�|����N���H��N�DN~�]��b�B�R�-�=+ț9�Z��t�w=o�/��+�<zdn`�<'��Gx!�M4	�`z'��[�s�h�P�$"]F�g��=�v4ɍ�G� |?�2���p<�w�7n,��&?8C�W�*IŸq༝U�cGt��P�$7����ҝ�_�ip�=�]��~9Z��厀窹��\���t ��px���C�޽/�4L��x(�����^�c�2As��9�>fqă�plG���#��)�38N�4�=uG�� �xxd��qH����p8#���#A�9 w5�ID��{Xb���*��g�)OںuO�9�.Z�/�j�J�Nrg=��S���yK������A�ۿP(��og�i�\ny>�os
V�oA<a�gy���11=0T�����v��~������Y�t��{�젱<Y�}��+���Q���\�1`r��W�[Ʋ*�5ʕ;Q� �32�*^�0ye<�] ��L�����O�J�6u��#��ֹ�l�>�h��4{ȍ1��熹����X�(HFa&��yc�ł$�D��.$m[[l
�vu�r������̳��1���u�[�*r����X"[��=���Y2�_<���4��U&(-���Od�'7�A��ר�-cSַc���6���r�M���z��1�O����謕��6���p�����Wy��/Y�Ng�Z��"�bK��MU)��k���M��f��%?��_.��Ӂihz�8�4U5�'���)KOW,U��<7nB�LY	���fwwX����|�����,�~�:���w(z���!�I�ct�b=s��Xy���v���~[�n���vYK�])�d=a+�.��;�X�&K%jv�qG�S��+d'�
k�^(�J4����fh4D��S7�ى"ڰ��:f6G�����زq!N�ѯ��<Zu�6�К�#k7��|�?'��Q+��SfA�mȭ��4o���sq��9o�,=� {d���FŕƜ,����GFBj¡sH�qh�c�5
nn+5�؊��yZ��I[�=n�8?�AOA�R���N,�:���^��Bd�4�7T��8���Ѥ���78V8H�-���k�{�b9>��1�9�=��<����;�q΄��+�<�qn��8<#��A���S-|��U��}�ݧc9Z�{\@F�7��?o�˞C'5wh�n�ǹr�Gq�l�����5�@��w��{6O���[ڭ<U���1�>�n��8����=�~�<������������O�k�C2���T*����h:�"v��ٶ3zo"ak�\o��_�DL�t*DC�C���?\�<�En�9Q<��ʘ�s��Ӹ�`I'��NSn6�?+SK�0ɯc��=�Q҆���ZQ���G=�tE�F� q"$Kn� �X��2�/T�r������A�$�e3�&������������=^.ےEKm�\�-��Z}��]�0V��'��3�̒K�[$��� MZ��N0�k��D�j��S62<hV�ɠק+6ݘ�B����y��x�J^����R!��;lἹVj�ۊ�mŊ6g�|ۺe�����t����Q�LhP3k�<u�۶c�z��&�%�6�o�z�C�J���$�}���2�+S��"�)�� ����V+�tu���Q�O[6A�!#�������뱅K���m�>i��,������0O&&����|R�'<&�j60<bO?��,X����S�w������H4DË-���m66�o�lݎx�a����َ�;�R�l���R�5�͞�*���n6��J���c���V�Az3�b��~��1�Iȉ�Ɖ"U5/ߢ��� ��>97����oS4��nti�B�qժU>��4����{��!D��p�_%��W�QT�y��a|^s����(����c���>㑧�U8*8���*d>7��#�<���w�f3�l. D�g��y���n��x^�}�R����O��I�n�&'B�6��p��ktG��9���UF�}	*�Tk��`L��~�)�8��{���wْ%K,��I[26�n��/��Bw����Vy��߯�O;�9	����ؘ]x�rt<���y��3�hvN���R���׾f<�����������:+�
���c�����/�Ҝ�\��k������Ur(�2Bk�ڰ�����_�*~ZoՐ	Oɠ7txl�iJ�����`�/������׿�b.��b�R��	��w�� ���c8�=���Wƭ��*A�w������˪�'�ڴ�a0�le81穜����r�4�'r�t¦j����C${�|�`84)�r�~��;��rҜo|>9i�A�7ϟ��C�j��І��&bc�3"A� ���I{�v�i�`�qĒ��!�)� /_�B0�3O>��y��TV%k��{�jtd#���Z���6ɧ&Rt>�4�l��+Ԍð'p-��������*��T�����Y9k�N[e|�*�#6�c��Z��-[��ҩ�X�S޺:���OLXoo����[�q��[����lgߠ�}�I���,[�[�T�bkQ�+�*ض�1K�,��cI�z:�
�<ڬ���M�ӮM�,�+Z:W�u}�jS�6�+o]�I���[�<lC��mv{�V,[lG~�-X8ϖ����ܿlRb���ў���c��_�L؎��홧�Խ���;��{���N������/���oЏ��AKY޲����鱑1���-���b*��q���G}����TӘ�1Ƴ���!J���o軙�k��<�Iڥ�\fS�P� ��Z�ys�jLC~;ag�}��:)�uy~�K^b�y�{�����V��4]�T�_�R+��	{��ߦ�:�8�2�[����Fm���������!B�!}����5�:��õ������FF����[go{���0���+����g����?�oCC�\�l�HE03̈́����hxp��E]d�w�Y�A��MZ�.m����鱟_y����Oh/"�ó�1�'�t��X7@���[2-�c���7��}c�R�8q~���/�YӞ��>���hXB͞J�-��3ϲ_\�K yz;������������/��T����e4����׿���^9�^a�h_��/Y�sԝ'�Z�T���~����J������W`���6gv�*X���ݝ:ϵ3�>��	q�Jƈ���=�.��+җ`�dO̤2��g�<��dì������V��|ݎ����c6o�|��~�,w�Z#H�ܯ�~������Q�
�}��BD�<�a��S�t([�s�J���N;lr�{5B���{��~-���;11�po4�-�d�?L`g��H�M�����O=i�c���8�/[�M�������:˴�7��u"C��^�ˤ�t �@pcs\�`����j�:�"�%�cL��0���]
��=�y��0��"v�iT�D��*���P��v�������D`D{�e���H��=Q��x��kY��ɀ��EӰgĨ���,W,)w>��Ix��v��Y�\���ꢉ^;:�V��[r�t�떨���Ԙ�tw�a/|��ң��~3D-\c�Ȍ���&5�=�&��6:2f��C6^�ج9=��Ï�c��Z��Y��+��Tض�����:�
-ݖJ�����6+�ٜ�]�o�����o�~����\������w��Ƕ�>K;mz���!+��V���N>��v�����M�m8W"k����ަ0,ry��A�æ�?2*���'��M[6y����µ3p<v"W<Y�=D�f�*Gĸ�ܾŞs�A��ם����o�َ=�X��> ��iE�	��;�-oy�"���� 0�!��n_�����r�ixb|���a>1�0ڷ�~�%�!-����j_��W��AX9#�c�Vj�s6��d��
���7�N�=80l����1�c����(b�;�ܝ����`3e�6�è�w�y�3��9��#i���þ����Q�Q�T�UN�	'�����U�i3�t�-��?���v�?�ȀF}�9����������Ο���T]��M"�3>�ׯ��o��U�Oe262<dm�a��) )`/a�	,�0�S�&c�����[o���`0V�ߕ+Wj<����\L)-Z�&��?���om��w) B��%�s�ى�~�-_�Ԇ�Fm2jF��Ɵ���;���o��_�x<�y�3�l^�1�^x��!0�$S�s����^۴u�u��Y���J��Z��*{�_����0Q/s'�y�%c�zضmK�qT��`�.Q*��c'UD�G�˓� ��Iڣ=�u�,5� 
l���B{�ˎ]�@T�{�I�����j8∣l�A��w�m���`��sm� m:)�+<//z֞A?���W2Tь�zJ��rꋞ���Y>��Ͻ��o�(���<rT��	E䮷¤����t`�rs���=��#��Lt�;w��榣Z&h�9S��0�󐛟y����3Y�K���EDl|-��"���$�cc|�����dX`��d@�r��N�u�w�Y�u���'y+��L���h�<U*�nJ!/�}�} ���,�tF���p�L$�I�2��4͋"�m:Y��q��ڕ�跉�!���a�YK&�IY.]�jeج1aGy�������'K����s���u(Îw�x2���l�'���Mv��j�㟮�|���;�,��f#�S���~��ۭ¤��    IDAT�:�ҙk�c��I�a����v�q�m|�l͚mv�E���[&�p��A�ӝ���qء�����f��n��8�%x�i��<�.�7-j)���=c�����rP�\��۾�W-d)�?o���Ҹl�K�,�[n�E������Ѐ-]��V���x�>�%�݈������택�f��V�ͯg��)G�9d��x���5���U��w9!������z�z-�Fr�'pvҖ.]n�|��r�P:$�c���R	e�8m�R���W�P�&��Xy�"�s��w�~60اTd��JU덊8%8��C���Ï	�R  �([U��_p�R��*�(]�>��|t���!P�§�*e;��� ��#�?�*d���f�=Vj#���6cɸzi�7_�4��ȹ������P��\� ��r�?�F�3�M�4:>�n����.����oO=vuv��'Rؔ�bE��N=KZ�T��;�p�[l���6��GC�Vj�j�f5D�����d8ps��~�&쵤�@ �X�$8��3h$܍����Fʣ���A.�[Tjk�jeJ=:Zۭ��B"a���o�X�ag-��0�!�2# t��M4η;uBy�)9�n�IyҤ�fR�%�"}r�@��"�8r���K�i� ���D���K�I�s��ۃ����xX�9{q��b��̐�ºBE:��/iV��t�@"�����?�����������SMp�r&�WJD�,�;�f�d0���������
e/����kR|2�QI�k7����ϜGܰs<7�Zl������7�q��#��#�W��ǐӏs�ݟ���F~�U��#����j�-*)z�DT*j�P#�,��YN@�"JO+�~КG/#�\��j�B�5�2>x�\�2�i۶�i�f�Ҟ���&ldp��z;�-������)���D���,>ƮH瑪��gSd�"���m[�ٵ��6ו��g<������LY�r��?f�D�f�,6K�go1�*�9�m��h����5�����YWgɺ�3�uӣ��{��o�#;��h}7mV���Υ�\	�Z�Qo��0F�ǚp���Hk�YhMu�5Q�<��_ߠ�U����u*'|���ڷ�����T_��y���&�e�&���A2��&"�1�fI^Ƥ^������*�:kVWS�F�]�yx�{Ф�Z�{�L���<H��ym�}}���w��!Ig ���j-�VA�h�#΄��R�6���1mȡب@gg����o^��
Ip���ـ)��[W}��V.s�*z��9��c�o��SA���o��mB����M6j�CKc����ުSHX�+r��b�X
�T�gBN-η�y0l��>��-΁fB�<@$٭;�jB���A�w<-�ga-�m�pV:p,0Tp���CՆ[P>�Z&��:�V��P)o�;���R�^g�l�DO��:�5�e@ü��c�S�f9EA��QB'�F�6m��PL�"J���F����O/rc�6x��&׫|����a��\$'�[���:5�
"a�tV�-����MUH9��V�֦��J��j6��e�dY0��E۾m��4�:]�f�̳���ƭ��G׉��ݤ�T�R�31-9�r~��h(���ݠٌY
t4k�Z���5R�|���n��K�|n�0�?�G��!n��M@�DΠ��;���8��7<�N�8����9�#h]�ƣ�6���7W�+�E����H��aȌ����x�(=w#�����įsOH���;�`�eX1��c0������Z�e���^2�c��ʩ�3�<x�ne�L�����蝎d4�!b̧�}�F�u��w��e�{�ˏ�w���l~�խf�ccҫo)�:� \v��z�'$~���o(i��w��)F��Vľy�6Aa�n���s-�i�����l������!ڨ֔�{�k_+���O
2,O���X��2U{��V�kN:Ύ=�0(�66T�驆�9i��5�y���Qs�;>�0蚓4�!%ӻ��$r_6o�j��v��{����'&'��3�D��
���+mdd���Z�?*'����{�����؇�f%0��vv*�n-����xS�Cd<����"�rw�Z&��Z O���dRH��3��m�3OdCSr����!���8:GWo⅋�Z/[[g�xW�_�8���I�/7`���.�m�ҥ���G(�;��k*M���ӵ��c�jՐ?N�t����@�s��|��D4��P�򰀠��r�q������C�[��8Y�2&/�z��^'�����^�uI��R�&��7���=�kڤz.]�Q:��0@ή��qb��`.��a�x�M���(�#��ҧBkUwʕ�Br;rd�W�;J�\�uΛ�C���ʱ�{��/=#�.��:�Ϥm�0��Q	���a���q�*Ý"'c�z�:<%��=P�b*�F��v�Aϵ�j͆��l����'�W*N����R�n6�jX.�ٚ�x��'�u��Hg��-�Z#E�^6��u�玽����dVS��e$yj!�3I+�zd2�Aפ��l������'�������,f�	|#�O߰�k�?6�J��A�~l�1�fc	�흭����\���ռ�I��������f$A�އ�i�#f/MD�f��`*&�Jeظ��{0�L80��|�4�)�?jҽ�ʄ�_y.��F�l�t�:�KV*�mx�������;��V+d̶o�j��E�P�9�f1�8^�<���Ę0��~g�$_�b�)�v�z۸�ia�r0��\�ML6lpd�Rɜ�
K��������[m��mvO���)ٖ-����ڇ?t�=g�J�<�H����>+�5R��Y%F��r���4��\4ȵ�M�eJ���7w��[�e���Ӷ�� `���٠aS�������~�~٨\�˂X/8��:��9<���:S#�Q!��艏5����,)��MLM��=�J������E<$��+���s c�\�D8!�X�|0P@��N��$1(�'�5��;Q�7��s_���kQ�$ 	�Pn����`:� w�~���-r�x�Ѧ���-��0�	�����:�6o9�pz����gy>��Бv����]�nh�ߊ�B��fBjG$��c\H�8�2�Pf��Ip^����07=bn�Q�T4��|}?�X�f��sF���h��w>��)j�!�^����k~ϕ�������k��Qb�kk������v�;�8���	()`��ݹR+4%�=k�ۼu��OLV{d7+�VDQ���Z߅>��%�5YQ�t��W�|��Y�ت<�^��Q���������^�J�V��
pP�@�b�b`=��A��!����}�	K�ܠ�o�v�CN^^p?O�Lg��
5bn�,�cnt�ДE�B}�{k�(ϿT�'�8�������A�#�n�����E)
�}�@��58rx
-Fu�
=��}�A�����J�Z��:zU�S�.&mV�w�,���j�m%�S״O<��8�߭�����~��խ����A�v|g��p���_�K���� ���C:��7>c�7o�|���>+OL��7��dJ���#C�mۀ�u���%�WX!�fmm�62�k��ڝ�l�\�Ĺgۢ��>LW!� 7��Cޮ<9A�����/�ih�F
�~.Ay��v0W�U��~ɫ_��?�SO=�tQh':!�2s������;�����q^&�!ʦ���F$߿�O9k�	�5Р�]7��R&���Q���k��3RM��� c@�97\�GV!��%����6M	l ����u�׼�Sb��A�\�3s����אG�n��sHH�5�&�$�9��fpBpbú�5>�=R�*#��2���z�S{,	{���~d��4�����G���]ʔ������ż�!@�����-#_C�7���Wia�v�9��L��q�/D�Y�9o�Ü"r�\���l���Mg!
��1�aL���}�n:�1�^��Qr�bW"E��U�D��+\���=�〳���w:q�m�;A��q$���ڏ�/�G�������_��6e�A5���4P��1�Ц���1�/�c��hF�p�6BT&_�D�m��O~򳯸�뿘��W�^ͦ�*CaCp~��K��(���0֮_g��`�8s�Y�����q�Xt3�{a1����s��,� ��"HAq���:��pMN�E��7����l�3��0�
UbG>:V��B3L@:��|h��bTW996�X	i�ŋԵ��%&�Ԧf���<�8�r?�ڔ�ѓ/[>k��>KT�?6�o�{��y�-�O��Er���≄`�9=�BA��� R8��'��k�[	šL�Z�m2T@����=�����u�Rο����u����Y�2�=k�eS����ł����}���n�9�նi�F[�p�f
%g�d��G��R-kx4���Q��>��@�h��z��?��>�+�;ٚ�����y��frp2*������ x� Ϟ=G���op����''HY��ggttt)��p�s9�rJ�쀖E�>�(�I�2J�п�E\��zJL�C��,ɡ;%`�JE}�A��dLo�t�>"t�Ux_���qr�t�*���>����Q���g�A�"�pò*�׆xSww�I���b�)���T����Q U��-㜀8�`UN��܀�:��"�!Q���0.�.#V�7�PK��C� k14p�!2N7;��)�ReR���x�����y���b�1v'�p��������:���������xnd�7JR#8|���nw��\v�Fmm�nZ��5�������J��$�bA�>v<�#]�`q`"'��^�����q�>\S؏ܩ��➤3!M12jT�QYŜ�G�'�&P\D�#��g�}fKuB@�u t�^l?�Tq��ں�Xy:-��5�Wr�D�8�S/��֛���޾*U�@vb����V����C/�c^�#�=��Ơ{��p7�)��1�39���65�#�FpW����|#����:����#��~C�Qx<:�=R�'	��0=���7��!_�� �In��AM�rSH�����u6�@�<F��!�iLU�T�����"��	A����׬P���V�R"�i�X�TY�1U����w$C�,j��a@8O����Ժ��g���ںm����-۶َ���?���X���4�9�T�Z`�������m������_��X��T�F��r�B����2Em������s�,z�܇ 6T�� ��D�䓽-f W�tHu*lbO<���p�v��7)7α��4�Lh!�a�m�}Z�d� V�uVkJ%�� Ёj��կ�7����o~m���U���v�#l�D�l�aQ��x�u��,���z�%I�u;���:�0��o�2u�u`w�����jL�I���+��w�R��'�����ϤlldL��ԵCb�D��)S�u�8���.z�|��@1ʐ�7¸� �x��&Z�^H� A)�BP���L(Y�㣍�Ȭ�Y#�՚�
E�OU�s5�VVA�_ZN��mn4�OZ���H�tth.y����%t$�F0�S���
&����&ً�r2 %N�,�MIϙ�"(�i�#�<Y�d#a�R�Z�%�A�	m�A+�b�$�]��_Z��G��:�HX}lB{�ip)pU�:�q&*�I�gH���r7iuD1n,-'i/���4+���2�i�|aƑ��(�Y���EU�,��w�X'ڋ8�d0��-�#����	�Ad��#%���$�&3�������͟#�M��p�Z��b�9U������}�~�9�8���o�B.�]%/�Jy�x�N'�\�v.���GC�R_��.أ^>ñ<�ozlʇ�`&B����XH�#��i�Ct�=7���<�þKT|�\f�`sD�7�qoW�����r$�/(-<����;Ԡ�o�?-��MTW�Ag�QϝL�"@��/���h �'��56��deT��)ki�Zmjܾ����q/?Zb1x���	��3�p��rEH9�r�8'6#���G�э#�EQl��dh�Q��#�AI�n� ēO?�2���|�l��vE����p뚽�n��۱e��͙c��	�����=�����W��E����Ȑ��| �W���8�?�O�SO=a(�-��@�T�TBf���p���5��AP�Jg�����9�T�"���G?�'�|R�H7U��h�*�P��3
���R��3g�mX��<p��񏿷��;lV�,{�O��|P��x���w��˝��|���)Q� P��XZ$��h�ލ�|oԒ��ǉ2�=={9��r"���\6���B��͏�߻_�t*B�FG�l��e����~��J��갣�:Ҟذ���6km)ʠ�1Md�I�\6�/�?l�S�Qw?Z���ș�	ׂ�!�K�u��%���1������s=<��������X�*W��(��"Db��V9�$H]�s��	e�����_�2��7��S:#��`�������	ֺ�c��C���I�ҧ��lmR��DdJ)M�	D��8�z4-<������TCd��ך�=���~fұ(�9�+|��/�ݛW�,/"3NQ�� �c*�?�za���rZ%���w�a�[WO�m��o�\ɦ�mR�d�V��8��s_~�Mw\�Aw&�,�ա=��=��j����ckk�/LgQbН(G�--�ߎ���EӉ��I9D4�z0�@�Uʰ�Vj�{~�߳�M��Y7����͏���2��?t*��#ڐ�H퍒�f�Hq���?����4#��')�C�cP��#���Q��H�9I{K�&+#�Ϙ���W�9�e�]�!����T�{o�A��T�/�A�i1���Ο?_����K� �D�ZzW�˖�pn�^�Ɲ};�,nuJ�5wڶm;l��(לLf���Mo����b���F;��#,���!�_eg����v�r��m�vE΅b��9����r�:|=����x���d���f5��ܙ��R�omm��g�ŎM(��fB��5���h
.ɩ Ǜ
d%�*��p0��jHw0�)�\��~��/}��̝m##Cv�i����<�$&q�`���#c����6hI���{�;���|)#���98
��P�����g�ϩ#�6�`���*f���=��9�\���#�ZY�l���y���m���X:Y��}�=��C�u�Ӗ�W5�!
_�d����	N�L֬�g�-X��͞;׾r��m`d̆�&�Z#j�26A�Y��qܠ̤h�����!�HU�c[�=��ݐ�I�;���V|s�S����w��p�0�p'�%I.Xޤ� �ɱ���Xώ�F:{��q���!�q�|_ �b\Ik8"�`�`,�C�,zRO�4t�j��G��~��):n/<�Q/�	l�����#">
 ��Io�&�A?A��-T?�~�-[b۶o�[��n���WZ�X�}CVGų��ҹ�hй�s�9縛o��+�НA��7r���χC�j~���6�k�`�snН$�{<*�^��g�n�Xd���-�i1�������č�G)��L�Z<�ѭ�u]�}��S)�퓂�ߏ�1輟��c�)Ny3�t.���d"^i����4>�A�797Q���	k-d��3�������ll|�ZJt�
�+~y/e�i�v0�3�?%��y	*ߺU���">D��L�����hC�����&c��w�ޏD�7�h�>���v�q��_d�;��7��{l��s���p[���S����˥�6<��ڂ�G����*ET���%�9b���o����.���;�:poy�[��^*34_y��)��>�;�A#�`xtD��㏯�v4��@c��&-xm���!ң'BE�?�����Ȱ���9�(�я�=��#�sE$Ш��"��04W�b�+%�;�'��a^�<t0��>��Nd��y�����E�!RQ�� �o�R>g�L�N8�h�ٻ�
y�v��U��}�X�-��pv���d]�lGo�-X��Vp���s�������w����ќ)pz�Gʕ��G�@�aQ
M��B�h��G���E�w��<"�7W��    IDAT�r��A��!�]"Ԙu�=�S���/���ݐ�1L]o*ڹ���4葡��|J�\=�M��e�AK @�I��4��C}�l�輧]%�\\B;8*3���%0����m"!1��t�*N@���`��q��I�"��#��2�pz�;5�zw�k��y���6[�F�����ދ�#�~��7���|>��	 6�O�x^5�s3�g����X߄����0q�l������l��rw�=1#F��3���ڍ�O�g-��㩀ݣ������/��#����Ь&t�c�c�1p�����[�'�or~8"Lɳ���i#^/�F�Kk�h��9Ϙ�p����K� x����C���(�*�>���4X����#*�;�C;�V7u��,	ģ��[�.� X@��~��P�J)a__�m߶E�����v�=�q�=��c��Ҫ�x�O���m�[o��^���?����Gϴ���$�w�m��'����1_a��DB��W\!�: ��:H�50└1ƌ���XӠ��I�~g�J`�o����,ۯ~�+�����D�N�eG��#��@��`������Tb�2{r����HTI�MِTC�SX�!B�7lx���a]�E�@��|r&"�HY����cJm!������}�5��J�P��9m��f�H0SX,H�^�����߶~�#v�=wڡ�bK-�����k���y�.�̡���n���7`�j�v���}V���U���%���4+������P!�B1�?�!��)��6�Ȱ���p�"�h �H)�)��l�<(j��{�Z�M-����8j�G���?c�B�?�}�=�Hd'
�|Od� �Ŝ
�h�B�.Tn:�P�)��+EêL�?R� ������H������S9	 +�@��}���<S^QE�N$g�G� E]�"�Q0tP��TH!�MU�K)�-X�Ш�9JY�ԡ�Di/�C?�s���[/���=�j��t���'�\nTV��xk�3ɡ���C)�k8�N��;��ll�e,;%w*�|w�4��dO���#���<�@��G�pk�P����@�;���S��D�2��A'�.�Od	''Ր�\,c`��OM��^,��>�Qb"_u�b�4��iR��{D��A�U+���\n�8�ejBR,�{� �����81�C�C���*��NQc�e5v "���_x�΃��8��f�-?��s��[���m�4끝���'��[oY#E��s��)��fk�>f���;��c����Z1#��g^����a����D����ۥ}��_�Z,�V��C_�°y傐��< ��  �J�	r�[�n����7Xa!��Q�6k��t�M���H��b�ר�E
Tڔ�YK(?�w��.H�.i��s��>��K>5��Q�*M��M�En,������w�]�G�('G������L��3�aOس,���szvy���5����i{C��.ٔ�++�ۗ��y+��v�9���JĹ�a��+�N�����r�/��A�����Z	�jݶ��K����Xѐ�t�Bbw�ĉ��&GG�:pܐ�z����!�Ǵ���aP�l�o1�7�i������p��	�7�ܮFj&X	��N�U����cx�PȰ~�,24��U�9n�=B�A�CʋH�Qd����Q��=�l�͓�=%
&"��K���ߤ�ݠ{�b��,BT�H�R�3��|e���{��l<
Z-ͥм(A��NL�`��6��A(�[9t.���{��7�ri6�;��5$�``C�� ��$c95u���A�|y�Б��=*WH��מ��:�u���C�>��	��Qozd1Hl�h<>���l|����=��;	���{�]IK���d��4�IFz[{�r�2�Ţ����M��&���6]���ļ}�;wR����b�#��R��o~�3�w���N�n2ec�L
�(��� �#��A)��gm y���Ԗ-[�T͜IT�e �
"(AG$@�3�t�)�3�cc��3O
�^��	��o�Q���h�r���z�[m�k������}��7��[�x�Tj��/+�C�;����x�F���1�+���Ƹ,�Ҫ�tϒ���߫����7o���=��0��������< �Cf��K��G՜Q* �@�@ZD��HF0��6U%U��Q�&KCu $"�B��T�I6V߈f�%\���vs]��g;�3���􈯋ݍr$�w�.m���I���!�U�3���-�ۚ5wXg{Isi��N[�h�-Y�جV!��Zz��xc��ٸy��wu�hyB�p�Ԗ��Q1D¦4��DV9��HF\)�E��r̼_^���NЊ"���Ȩ�S9��A�G(����Q��Ս|:*v�:w)Úi7�
"�h�i��#��ϣ:�{98�in��aj
%�R��Pܠ���m�5Ƣ!�A�p&��m�#��.�%ʣ�)���;��en�Ȝ0�i׾�[%���`�9����P��H�)��b�M#��/YM�� �
)��:�쳏����/���:����%D�Fǻ��5LT/��[�~]T�>6A6~&<��\Q�{.:ܴ1������51�5�ͫ�}��("���	���=�o��?��O��D��ݺu��ҿ�rg	�HowV�lN�$A�ʂ�{f�����3��u���ښ�j��7k�	�kҎ�o�r�ڥ_��Xf����3� �J�-f /�k��J%�� G�=c�a�0���c���#��FQL ����iaA6�!�ܭ[�x�ي��7��w�i[�lS=�qǾ�FƇ��;�����Z��;�z,�$/U��Ĉ�ܹ�.���l��v��'�!�<_��G��bZJ*?��_�b�J���v�u�YgG��#�ȇ�O���~���|��U3�6n��leɵ3.������f�����T^6U���׷�)h�"t�� ,Dޖ~�D��Hl>����D,D2�H�NL��Y�W���T��K�l�nD��ƝҦ�TĊ>�*�˾�=�6m�{H3�9����������.�Zm\+rT�[�i�	E�Y6�ʄ�P���Hy�ZZۚ%e8yT,lx�	E��RQ�Fy?DP#�V���B5�A
�uz�^[_@6p�@D(�A��#"��h��ꑈO=�"% �P~�eW�嘁v'���se�A�sfN�#��)�m�n5	�;�Uf�н��L�r�@�.��]٤H#ڪO�0d����Qyrd�)s=�g�cӜ�Ў��4��3��7�l�
%� Jk ���>'#��fv�e ���B[o]s$��G��B��~��FҲ�9� ?�|�2����v��������/�{�G�r˭��r��`i�A�\'����;Z��1W	V�xni))���W1��h����
�67�~�8��:�1�����[��!�jVYV�"��;����=�]��Dܠ3���M��Og.DA�#�SY��ɢ�zۅ�͝?OD( n"�r��.{���H����o	�ߥ�9" �=dG#�-L�L>c}��p�;`�J�����+���и%�^[�~��e�,�!�0CJ��Y�0�i	]u����z�[r�Gu��_}�ua��SO�B�ݜ�5z�<o-�1%GO_d�ٍ7�lW_�A���W�ƶn�l�����SO�|��A�B�ϒ/ok)ػ��.{����V��w��^����3}ϙ�D��Їԧ����5'�'��^}�ډ�����~�/Pچ���A��q�3��a�<��!Y�ӟ�d�+2�R����C��fF��:?�ß��Ĥڻu�u	v(���P���� ��ڪ�B����FDe@�_M��H*9�(�(�����B������݄9�&n��<w���£Jr�@/%��Q���Q���H�p�9Ѣ2�l�$�k����BӐ�	9e}��I��q<gJ����X�3�g�b�QÙ�*�:82nĢ��:�g-�
F��A��U��z��8c���=�3Bo
n��f/w��d�q�HI8���7�����k�N�
7���)S�Y��G^s^DppW��Q�Ce�8�S����O���h���DN,i7���0����rŢ��s�J�"���EI*�m��"���Fjz:��9	�T�I�b�&���o�ZlO(M��zP����Yg�}�;�\V�VW�h:bFu�L��y�[�I&���ԈTi݇��Am0��J
6z��O�d���M�>�.j9H2��Bssu��-	݈�K�q �c�����ϻ ��
��ĉ"�E�H��������PYH#{�V�đtv<�����;�5�[��9=s9?��f{�ɧv�ޤ����J��j4�կ<�>�gآ�s�@W�D�|^s����]"���S�l�w������d�ÔS]��_�e�]&x�?��?d�?����g>�	�\|��v��G7#y��Ѐ�+�'2�;�� '����%�|�6n�l��-�#�8�}�1�����O��ș��ɨ��v"��O>�N|�Ծ���>�tF�k�w��u�Gy�}�#�����A�y�f{ӛ�d_�������?�#�8��p��A$ Б;��sp`HML�����/�F3�G�Lэx`�+�ěR�$s�J�:�T"��=�΄nN���(u4mƩ��F/�# �����2� +�|W�t�M�L�ܜ9rX�֐:ŕ��WR��;
:�ȕ���:�*�j>�6�Y���$G�jET2цXHHE�Í�p��C��7lR���r� a�"�]]$��F�n��R(�濺�)�����1˶����� Uk)�΋Ac!ŪSA�(�I���XP[���dĢ�wY ���J�ҘH���H�D�]�����>-@��� ��!�i��F��j��jMd/�Ix3"�
�IWG����(�P�[Z�"��<�}N�M��.ΐY�l���h~�MP�d
�`��t_1�㣣��٩{H�a�����m��mo�Y�ݶ���R,��Y:���ܜ!~��T�ΨM0{�*l�62��L��O	k�m#4<ꚭrR	w!e�3�0ٰ��t�Z�MUR�d��0��d9k��t:�,�ꉒ%��L�X���gqz�?�Ú+�	8�t���dp�5����g�y����q�e�db9�w	D����B�%_�'�̗l���|0����d����Ρ�2������μf��ݎxN���{�:����u6iw��3�(n2�R�y�$^�����p�ٳ�3&�P�֙����e9sY^u#(v�I�^5�4;�:�QO��аMV��T��@t�}#�*�c��1�/Y��לt����T/Mkj�I�Qn�������_��7����ى'��h���s�����?���=�\{��o'�x�Z~���W��SN9�>���i� gl�;��VWG���s��t�JƋv�\���o�^z�"�ŋ�ؑGe�<��q�mv�����?[�'^<}�i4½���7彿�ŋ�Ӿꪫ�(\�׿�h��������Dd�Gy�>��O����OZ�f|/Ft��_���qU��1��c�	�F2� ������{���\p=4�	�Z�֋"��Awt)��Md$$�~OѸ'ڬs9�� �Yk�Z#t�S�0GFe�D��8"�5E��,�����.E�9��R,��Ҝ����o�k��C|Oq���j�]�գW7p�_�Q�����e��K� 
P�c��K�w2��WĔ��7i4�\������۹>A�	�����������ԐK#�#ڨY��)�Ѵ�x��Ѓ�Z>ע��Q�;Q1���nu��Y�;�s��D0�Mf{mR�:m�V,)=��w������a�_�q]�k��yYb��~%uF��y����Q<�E�B>���lYmX!��Y��-�S
Y�)��z������F*�s�U��U���^���u�� �RnukV�`�c�d�-^`#C�
X��!o�\�r��jr�ptK����! �1U�Z��F:���k�H����������e�0�����m��Ŷ�{�p@獳<Q�v��l���H��{����T��z���}������d"3:<6�oht��X}�j���5K��R���T:	
](�$zH�J�8�:�&{�^1���������.-������˳G�M�f:��!7��D_�6�н�����W%k��$�EgS������>9�.RR���GP!�U�a�Z�;����N�إQYP�^�����3�\��ל(�sL����߶ozMX3���:|'c���p��6��ˠ	�M�Վ�D� >�i#��)2訹I԰ְ�_u����l�K-�Ȣls�ϳ{���9�l��o��������6%ʩ�9��6w�|{�[ߪNbD�D����'U�d��OVc��]�i�f9],|6<��u����elp`X�z������v�z[�t�����;�C���϶jT�����)�!́3A-��g~T�t�rm��q�	�6*�kzJ�/�x�;t��x�+D����[u�ѹ��CH�ײ����.�dt$��`�q�z08
�4?w�ݣW�be��2�2�IP�d�G��E�*]�)�0��J\�'ʇ$�R�&B��j k}�̳d�|�p��+ ��	eo��U˽��3&]�%��*� Ș�R�����{�(�T\68+H�����ǡ��⺅�C���q�)W6��'�[Z��
)��yH86X���9k�'HRkG��I,	�T���Yg�l��9h�^�u����mb��N;A��Q�[���a3z��\D"*�᡻r�>�X������G?��+�۶-�Vjm�R��8 �F��|��g`sGfH�i� ��5!r-��C�es���)�n5�h�S��,`.@������l$4���:\�dG��:���Ȱ͙7O��A�0��o����a[�h��رSץ=9r$�����R��*�\���]�����G��Ouq~�ϬY=��FykU-�7n�i���mW\�7;דּl��+'w�n-[}r[:���XH���ӭ/y�Q�_y��QG%"&T�翻���7>�}�C�/���Oɦ�ǌN���wu�n�D���v����H�I٫���q��}�%�\n?"�d��=��Dn����z:,��Q�y ƅH=@�rQ���������=Ro�����)K0�ΪG4D�.��m�rJ ��X'*)!��"�Ot��}d�a�;��%M䚹�m[w�����O�Bn�q!�A'����z[�;����ҩ��2�CC�R�MBw;���CH�S�"������'�l�,_��^���'7��"���>'�%X�l�6>�I��ήvm�0�1��Q����2������x{�g䌨�,����ڸ�t�b�|�@(q�_6f�h>s�]��w����`Џ:�X{���d��9��v��Gex�nR@�Cڔ��ݳu����huGs̏�{��CJ!D�I��8��XpF�l�w��k�	Oj$��iSĠ3n?�(�R"U	��ƀG�l����ܧ(�7�WJo0�Zl�R=i����;���P��Es5���XG�\g�����15����H�L��`�dD�2��Dnô"|����]����AJ4�c*u,
�w1���a3Нg�A87�����^C��x�j��Ü*79����x��i���0��'$"�mپE�.�wߠuu��x�-V��5��-v5(����Ҩ�)���/����q��"��"BoSʾ˖ے%�lld\)�<*'�4郃�Ƒy�K����{h�����+QzN4�#v���v2�qe��Q��� ��zs��Ozz�'�����t�snWt�w�@G���&��Hߛ|q�;�:Dz���Ino��q�B�,<�M��R�ȃ:�(@:�RNj�K�j&�f��P�5�*����n�+~�S۶}k-������u��;~����׾�O���������?^x�7u�}����{�!����Fʦ(�-�-ZK>�����>��5�^�H$�s��9r�:^��=��Z�L���wh�a�8�C��b�Gr����    IDAT�m��Q���g�!3#'�x��>����ql���^���$\�;'�)��n5���w&�q���a؄��;��7O��W��zab؁;�~#��+O:Q���~�s���1ai�P8Ǩ�G=Q�VW�k72�{����'oKϷRVu��/Zh��;m�]w�����uutkÃiJ)��X���Cy�Ϲ�ʠ]3�\����hT��*�Q�)�aT�#�|��۔�ƩY�p���W(B���5v�Y�!�J��&݋ �Nkc����8&����l����g�����T|���{�v�iB���8��:��?��?�����Z�d�>ØSg�w�7�0<���{�Sj���b���A��`E��]b�Aǈ�$ep R�Ȥ��g���J�Q�`dt�����L���?��	�WW��\6o��������C��]�>7�M%��,��	�tAy��H�����ƅ���)U!ʋ�:�%���f.�XKg���kr�X�Ir��M���@��?"�48<lm�-6D��5�@�TKLOArʫ��:�!�r.������f�L���[K2t8�LV	�f"�-��EFLD�640(��jh���Mӵ+�A��(�}�4�b����Q�Ż.:/�0�\MOU�� ��y��A�Dklg/�"�9;�6���|�I�sV��h��_�<l�Ã6{�����FkJ|�+��D��=�[@p�(�lXk�E������_��V�L��3���Do�~r}�L�t��Ĕ͚3����Z�P�R[+�k�:Y~�Q�|�������}�����W_}Ǖ��v��7�rf���ŕdv��tڲ�NK�l*��^5�k��r3�Ag���pyvQ�9967���ha��q�&E�Y#}w��ȍ�<.�����(ݽ�]8�e�6�x$��bg2�H����o��ҍ�nJA���l�l.�B������?4���Ƞ�GD�,�!�u��׿�m�(&�Tǀ�O$$pȡk�:�q�/�"9�W��{�O��{����=xr����S�~�ӟ�s�s��'1�\��~�3A�?D�tLc�Bx�ǵc���w_�� ==��z^]��Pj��9r�V�������Ï�G~�x�>{���&cI_t�B�s��Pi&d�1��މ�pF0،����>���=>C4!�c���~��J)�Y�F� C�u�����/|�6	�yt�}bD�#�c��@���)EE-����O����w��=� w��5Ł�Al	��=m�4�IH�C*h�����TeR�?�*P��SW�m�#�6w�������N�Azc��8�r��!E��.��ς�݆�b*���>1�#�8�q���3oC{�9P 1Y���d����Er�{c���M�X�����uvv�Tm�jպ�'sfϱ�;vX:���Y]�����h�"���l!k����E���!��γd;!n��g:iS�r�*{����ϧm��qR ^X����1vt5$����+�y��W��"%�*�I[H���C��"�,�9�2g��ɡ�f@��2�H�\_�}
��t������~��������ۂ��^6�P���`�K��je�J-�'�Րu�SԿ�/�j*m|r��u��J5 /�[7[[w��s�a�4utS=?�24���'Ӣ��-�T��m��&�c�!m5V�A��u��yN������;>1&�Ṱ���׼�������N�_X��n�T����_����j��_���:^C�
~E0�r��ɡ���8����4�ɬ���^��ݠs�պA��s&�c�=���ĉ��p��p���h�F]�<o$�8*=�G�|��i>�f�ם9�5/��8'�x���q-ND�G�oXq4��ϣ6!w:xCŹhq������{͌�;��Ë�Ԑ������ D��d'������;����iˤS֘��/>����ۢ�󬣵�� Þ����_�M�1!B/�Mb'����g��w��.��BA�41�ꪫ4�_����?��~��_�O�����'�}C�u�ю���a,O:�P�U�6��;v��!�aйGs�γ�>�֮['������K.���͛��c��p��)��>�1E����O��+��B��y��p���^H��`�cؽ��{��^�k��#<����e2�>߸���P����3߁�ߖ.��Aۂ��״N+�r�hه����Fj[���������ẉl���2Z�8��o �H�ٝ*��G�HRi�A"�N5��)��l�2w'X�rM�'������2�kZ�.CQ�Pe½ŉ<�c���$� ��֕W�T��^�*��Y�8�7�t������U�W��d�N�Vɥ�����Ν�v䑇[!WT�b�h�LF�g���p���ب]��_�u���
�mbwi�������������Z��))����G���R�X���%N2!�H�wk��F���8��@�J�a���V��47b)�AX�*	̀���=�pkEh*Ry��Z'�$:d���o/|��l��+��_�B{޼�s��9�::[�nٸI����J����z�G0�o~��^���q�io��?^��w���]���y�(�E{��/��;L�w��۲e���sy��zʛUـ����9�ß�Lz�=s��z���r���g���M����s����\&%�(Ɲ�K�,�SNy�-\�خ���v�5��i�.��jet���ƃ��w�����v�����]���+�>���ή�v<�@4o�B2��A?�3��������Һr|<��94g�����������0�^㰙H0�b3��̉ĺ���tҌG�>�n@���d�'�91�s���0;�E�è�Q^� � �F�`�n��i��"�t�q
��d�]��oj�W��K2Ec	k�x�~��a���/)gt���A	U�V�3|��!j����Ӣ�R�<� �緼ٖ.Y(�.�u������yJ�0��`z��J�x�t�Ia,1|�#����)�Ⳝ7�`i�(ca�sf�Q��b�8Y����m;dЁ�1�|en���O�;����Vڏ�#mҒ��&�@�� 'ǁ����e�9B2]t��r6� �Yg��(���/;�H'�a��D,���0y�|��T}�;������W_�R����*��Z�F�jQ钬WDZ�uf��&@�Q�\nS�`#ZA_o�:R�ɑK�� �å�P�Sā	�8 ��	T	T�hI4E�-�(�=���m*�1�jͫ�����5*�3��g�Y�� R)Ss���a�ONJ���}�~�]�_���/s��O~�#ݗ�����O^l��{�P��N;�>���ҥK�5@����~�#��e�_.��U'���%9\��G?�Q[�~�]�۫e�~�!v�s�k?����?^����N�5�EhF:m�����m��裏����V*!T����/604�ySOD:鴈����j���vk��$���G$px"ޘ1�����9�/d%@D��k�1�m�<��=�����Q����=����c��ן���������Y�4�㒯~�֬�˾��/��B����W�z��_�L��җ��>���{���ؕW\iK���\|����R:��;����~�[u�O}�9�T��е�uٿ��]j|�=g���)���j9f�W�g������y=���.���^���)0�����~�.��[��>�ڷ��}���~.�%�#Y(�7զF����ν���N�?5�|���}{�O���S�Gk�ʴ�j�%
�����3?~�m��~Y.��O�"'���/j��%l�*G�~6l��d���<B�=���)ʌo��f��s���g�����wэ��D��pa�E��<�A������;�Ht�p8�ʏdj�_m,c��A�;��A�5�^�!O��sζ;Y<_�غ:{D�
��GA�ٕD�'C7!]k.�\��j�b�{�)����z�:�ޘ���6E0R��1�����YY�t���=�Q9��3�LN�c���G������1h�s�e��������@BU���`�{E��PAAP���
�]�+��`�(�H/��dz���;Y���=�=>�9����)�s_�,��ޭ�T��*��+�=�9�͙/_s���l"���ZV^!��}��H�~ܸ��KJ
���$�]vtǆA��1��3A�Ю=�Ν+I�#7t�#+}="�1���K-Hy��mu"����(0U$�kv����u�y{aQ��	�_Q���������5��Y��PJ��ZDx"���"�%Y���@�h"�P����%=����`"*8���ziR��0T򢾶AQ��
K����j��:� .�ﬡ���h��J�w��I|��hg�q�4��j�3������	��ط`�7�k�9�\��9
����m۠q�^L�1m��$�:�\p�r?��,|�]I�֮[+���uLD�?�x�8�f� Fd˖-":4��+ɟN$D���̕����h-*���~=:�6lB��2��)*KYU�+Ľ��!k��}���/-�i��e&�c�
�����t)R�1e�Bœ)�1��hv��uײ�j��1� �J��H�����b�#�E]�7��2��2��i g�7�V���#��q�n���n�ʯ���ŋ���ob�o��C?s�t��5���+e�VW��AÍW^oq����}���fc������^��7^��'�UE�y���q�q'`ƃc�u�c�}(.m��F�$]+;c��w�h��F\��3g��a�ʘ�Ӈ��1�q�Y����W+fPR1�ҙhƈ��^=;ݹ��ז�7�9?㻭[�z��u��ݙ��+�n���nk����Z-qc9��uu�۔��g.^>@���TۧJE������]e]�����Z��\�Z�L]�H5xO���q�E���|Aa�E��!�0�C�M�|��l��骓��,=	��*L��q�\��]����Fca�s.Οg��dɗ�9�)Q�����{>V�2C�+��~Щ�^ֱ=|�u�:�?�t�V�<�n�&+��V 1�rz�G���R��!e�C����7˦u�q'H� � �ky�Ygaٲe� ��q�TJ����<�Y��5ջ��+@]����}���
Cr����>��6�>�A�˓�{:+���%�=+w�j��X�kJ��
�\8Z��g�'�ئ&9G���3i%�J�M�?���$B��9����Ҋd��x��������� �;O�.�o�3�$/9�&#�	�-Ҽ&Ǚ�1I�DXE��H'���Y�(�TO^~�~�T�w���+��f"j9�48b ���]���2a���ZI��=����צ4�u��D���2�*�H��p^�}�C)��Z45��Ǩ�#��3�I'бC\��2��ޥ2�W�|}�.��[�Fޝ���|G\ ɸ`�ƠĠʎ!��K��.�S��7_�.^o^>^��WW�̳��ò;��
h���d���+v1�p^������G1Ｓ +W��D�sq�;�J�[��t�DL��Xk��ʜ�k�p&rY�*�G*�t~[�ja@�X�P�t7&���׊�������}0Ќ��=g�u&��f���v����~��>|�k�ph��H}�љ2�z��Gѹ�B�x~^�����_��Eb�֭�6m�xP����`��A�ɬ����T���M��9/c�9�ԹR�ݺc�o[䙡3^QI��r�!�"�	���� ӧ�-�+�h�v��̳Ͻ�޽���SNǹ�]�=�;J�#�D��믾h�C��n�ot~�u3����꟟k�em�Ft��RܤI��^����k/"�u�ՁMs����ۚ��^ �7���aKZs���tk\�r�s�� V:��9���Lt)�[�<^=���芚�/�΀(�Y�8~O��������5J���y�w������"J��}Ὼ���Z}��v�|��Νg��-z�_���@:=����F�2&dL��20-����/�QG��N@�,����\XU���^8����-�8 �� z�����İ��H!o�J�o���C�6Xy=D��h���}�I��1;g��96�:��*���C�s��,'�C?\�y4��g��{X_['`V
�W��	����~~O3 x�x��<g��ֻ���`�����Z��=ד���-�݉k��A��e˖K�!�GQ�f���BUuL�.7:v(~8[�R-HwR'��l.DH�2)Z'���R�<�b�)Q);��c0h�<:��N�y��!�t1�5�(a�*!;��R� ee`�M^�_K^���j��R��D	��2�lCi+��J���]$�y�[L^���ЕJ(�S"��w�GS�^QR�Z�E��9X��+���<�ȃ�\����+��~�T��$��.�a�;}2Ra`�8�s�ƦzL�s�8�qn��{b͚52�)i�+�]��O=�~�9�^�.��#����V֜���!k���H��4L1����&)�j�X�Y�6�	G?�D4*�7�'ـ�{�{m$R�v�T$�!�&X�7� �r��f:+v�7���n
��=M�
�Pd�bFsM��q<.j����\�	��ŏ����1�
(�����_,��O?/���6����=�N<Q:tL�n;M�;f����_ ݷkG]��}�`������u9r��^&�8k������9x��1祗е{O9x����]X��[�c)��"x�<�Ӊ8�>G�SO<A��˗���oĨ+�De�����V���+F]������N�>C&��s�θ��S���o�Y�~Y9{��/V��f�N���k�6s�����U�|���b魜�T�FW��AOK�� �+l����?���X���
�7Pϭu�[���־Z�z>�[N�st0֋57�П��򹕷���uB�g�:H�&�=�znGA�V*��\J'��.��9`�օ�69��!*�q�#�����|k.|��"���R}5��<%����;���,ݨ�!5�v�����t�T��o�e���:���GN�_���-���vvuu���q6�`+�f~�$���2����G_�T.��4\������9��ի��/�z�p�r->X��l�s�'ʚ�pW]5�f=����V�8��"��ب�l���<?~�����geşgK^��[dx���"uόh,"ׇA����~�����x)�7sS�o%7��Z#1����Ͷ��#�ȟ�8E/l�w�{��;���Ċ��%�)1�H���z��sp����?!V��M0׊oV�SP(�J�X&Or��L���ʚ��-�q-�p(w1̓�Ϧ
誒�{�-������%'hM���YL`��̸2R���tF�xn���c!�{�L�����~�2V�f�8i�$Y7�Μ)L���;G���_��n����"z��_6B ����Թ3���#|��b�u�D����hס=n��f�<y0���hBF��WϻQ���ZT�JP(A�GA�S>���p-��ȈO���?��ͰBW#vm���*�r�wDM��7��f�[*tV�|���F��\�O�x$��6��z��hWR���|8�f�}y6�}�)L�1�;���Ũ�W�s����G��O�)Sp���H��g��������Γg���ݨ��:
�_p�6�q�[U�~L�>M�p���}}��gpޅ��!�c_]n;�XUuu��ۄj��D0��q�����KQѩ\Fv��v�\���
<^7��؋�wLB(JeLbKbH'#MCt���_�p�.�b��^/�S����L]0sR4a��?ЧY�j�&���V����@�.j���0nn��4׬�A2e>x}�&���`�������V�7A�fp��t����xt"׭W�?�2�Q'L�Y�+����s}�脃���M9C�$j��f��@��(YF���о}[�����࣏�WP$����Eu}<��l�ՙ.�����8�Xn[\_}=��ܸ��k �`��غ}�2	�J�r���x%Xk ϟ�k&f�֭�8�+ϓA��(Ap��s���h    IDAT�*Z�˩����Z���J2D��u?�F<��
h�xƬ@�	��L[-�?_f䜗2��ضM*k�(�e�E�<��{��+�^k@����w���@f�N�2��"¹���`��ɧ�K�׎�[Ye(c�j�Sn�&8]D����G��MB�V�L�2l����`�<�TQ#�moS�>��1t���H�	����/���m�)B0FW=#)��/5z�~��NYX�ڤ�KdR�h��6щ���]=���UKX���yk���.#1�e�
cF4�V�ԡ��ԓNĸ�7�M�Bp����?�r�f�7`� ̞���n|��8��S0w�c�>�9�}�e̟?_�2������5W]-�(����/||�1�O���}{����/�`��WH%�[q�(ͫ�-��6;��s�:�vB���d�y�й�Z��ib�%9A��0���Wv���["Q�Z� )@ֿXV����l�3Η:�j�R�c� G��]�7t1SR��u$.��B,�b�\{�CW�ك�G����Ʊ'���n���v��O�)������g�~��<o���s1a���h�|�%��ݍ�/�޶m�޻���`աg	H� ��C��ُ�^GE�N�|_����㏘��#���K0f�X��7�u�أ'�%�[ZR���j�3q"��CO=^��~�5F\~-v�ޅ+F��U�\��[����F�I��r��L�W�o����s�ճ��[�_�o���Ӄ��x�5�������[+�ɓ���o^0}X%p1pȥ�� *��Y�����0y���{�شB�~7W�*`렭��:Y�U���=��s+~��?�s��r��ue��n�k ��Xe�P�@f?���Dn�Ǯ�凭�~ u5�/��"�D66��0�:����K>���}���
�WT*3�]���fsJOP�9��
��Bi��B2�1��ŐF�>�,�ɧ��k~���fU��j�V8�xN��h�P�?�*G(���͋�=�����cT��Y0w����5�]+�.�ƍ��'ϛ���t���'��l��4�;D��ggz~��?]��1"�RZ��QS���xL<6qI��<�=g�ɯ�O�o��ن������A��g�2����W]u��9��9
h��=� J��� ���6j��6L\ںt���b�;��GzM��3��V�W��P�_TX3��,�� ��]�x�g�:�;\0�m���˦m+mg�
��̂�G�6)n&��J��U��JVV�I�CWk�5��v����*��t�E�]�ٍ�$�2V�8�h��p�����SG<��â���d?a;����3���\��s����� 6�m2d���	�����p������ċ����&a��{e��-m']��R���,|�=쯭Ʊ'��Iw݅3�8S�]�T��i],{
$��b�IMs�hOAM͠o�ūx�4l@�v��"�9� R>��,N&��УHP�n��aǄ9�*VTB��9�a�aE�N"/�@��A?UY���K��(|v
����Ǻ���?Ɔ�V#�|��rt�섊����kx���0��s����c�m�Ģ��+���Oє��oźu{%Q1�|����`�P��z��M7M�I'���;˖��I'�_6�.�Ε�;�.D�������vq�磩��=z����wv����p��`�ͣH�ނ�s{0r�yX�z&N��ӆ��zS��K��F��UÚT�W趼:獧�9���B������3���PV�������6g9p>��ڬ�t+[�ƹa����_6H��2���ZW=7��Ur��Ź�N����Z ���C�ѝ]��d"��g�U5�9�$A�4_^'��y�q�~��{�=����**YY}g�M���oݿ?�~IY�rv7�*�b�νh����y�X
�7�7���U@��YmF�8�u��7!��㱇f�sE��{��JQ��e�b`s;�Ч�j��X�+����۷�(8�Am�X�y-��T���z܊������G=�H\:�2�𙱋HOL�ω���(Z�6���M:>D*3��֥��=9�g�ۧW/�3F�9���%`3��sy<?���PW��:Ya�ª_@l	�	
�-Z�yy9W����W��8�7�e�
��TNkY��t�(ݍ�����͛D7�IT��=Чw_̜�2i��|��#Ɍ �2������v4����B�=q��E`�|i��u��Rս��bX)p���$��v�����U�.�h��M�3/A$ӊ~��U=g�Hk�i�X����JdU"r`@�xJ~
�4	����ϼ���x�u������sg�p��D4�D��k�)�ֻ0h�$w�PPč�vr�ԡ� �H�㫄\U�b��*쩪J`ܻ���N��xP0C���u��HNv�i9>ۢ�B���	���N���1�h���M���̿�Q	褐r4��� �/�䖋�P��&��f@Ϥ��GA�4B�#Ȓ.s�wѐ7#�N���M1��vmJ���՘��x����6�С�#�n~�m3^����O)�/�H�7zL�6M�K�O6o�U�g߾}d�V^����E8j��e�`�TC��^���t�Q;�GO\v�e�X��kt,/Ã�>�R(��h2���&I@y��?����"�\X��stl����w��+����߭�����d�W+`q8KQ>��)2�_z�޻�u�2��/���li��^}����yl i4��}ڴ�\�b%���p�r!��5>сKg��z���*�lC�r�ݻ�E�T(�v�����ٿ
���-�ߓJ��*x���5W�9)HKE�`��D]s��\�)R��� 5��y7oTe��<�UJCm��4���Q��rBYʐQ�zY����ओO��A$�%Kp�e�f�wR�q>�JtPs^-(�,KK�f�I�-Fx�6�ݳS����}�~�3f�/�:�H4�JK��ܢ^�*FW��1�a����o�z%�N��L)�)V���:M8{�V (v����N*[��F�:0}��r�ާOI$�f���i��*b1<������v#�[�p$�;OZ���������EҖ3i�*�@���%�2{���*ry66�Ċ�D�U 5�uF�Q�8k�p��~�j�2��+1�l+6B�2�^_G%<�l�}9DZ�_~�N<�D���G��1qf����b�7=�#Z�f4#�i�����aäMIu>�m2 ��5��g���� S~1L��A����,I��8�����,ۻlϧ���U��Ox�������-�p9��,�M��ZR�s��r�-Ⱥ ���9���m1M<�(,)��/�\N�����C�PpO� 	����5�.5�a۞��������ed#�bJLA��N0Xl�:]�[���TQ㬝k��ky��1�3��^G�!W���ԉ�)c)P���@��0	��B�#�5ˠ�.Z�rM	Ő�&I�Y���VI<Y��U��B~A�v����L
02��&�"�uQvF2�(��G��(/+�gI��v�.�G���>I�#^W#��
`從L���Z��y`�^��f8�ά��E �\OT~��r�c2�u��k�.$�Ē8E�-,D�b8�`obl�N����\�$�;�4���c#�E�|iBm�^I�ڕu��r��Vx�Ѡ�j�}n3���[�K�\>f�k�����33�����l˽�!}��8���_��)��~0-�&�f��^��T�����T�V�(1UU�S��Y�9�P���k�]%n!s��[��V���Mh}_m�R��5/�IS���ӴAP��߹�J:M�oe���լ��u���MCU�����&#rN�����@9BV��"��%_`��j��"��-3�.e�3)�������G�����&�y�{�HRt"��l����p�=S��'�PDǎ��E�����`�����F �<%�x�y���N�ͷ�Ə������I  � ݭ��REmߵSڞ����)S�Ȭq��[�kl��Zq�Ig%k��{mu56o�$nj��9;�9i���E�_ b7��O�2	�o�C����J�O���j%�ѯ�3S���-r�$ȉ�,i9C�A6�Dm۵P]CS���h��w�^�	<�p���W,��3	�|�	l��E}��!���k�J��U����8�裤J'ņ��YO>!UɝwMƌ�?F^a1�Km�:ڐ6"O"O�a��MQ!�>ݺW⾻&b�k�����N���LE^a!n7��b�N��m�ǝ���B����*D�"�.�)�)X ��DV�LP �\{��9�շ�uyM�)��t�v����:������YmMi���hWR�@]�$)\s��4�m�2M��ʊS�(�a��Y�u��SQQ)��{��c�2��׉*�^��c�?r�?����{G��<ʓ�˅H�|}{V��]�f��^�D`b� � �u`�,j�Ի�E���e�htkc�`.g�4�$��=PW/I:�6��$I�44�۶���21�&z�� �]X�2G-�Ѡ�hi��}��̰Y���*Mt�{J�({yēhWR� A���0��;"����NgD;`5�� �Jȵ�Ю#�����'�HRI��V��7�R���u�u�Zk������y
D�b�J�z0����{�ȳZ֮�h��Uҩ�"����k,+XD����w�{8)��f����O�_�R�'�F�u��ұp�lH�Z9��ُ.�o�5����>��uk����Ρ���:�o�O=z��?��n�֘��
�7����.^��lYs������>�ʯXq�U�J��x!��C�ϳ����A_W�j��k�x�	:�?��O�i���~O��5�@��uW���.�ȝ�����T Tl�N�މ�%���_�jC|��D��ђ��d����t�4����p9����a'�Ո��*�1�v\{�5�'�Xֻ���7�9Z��-F�����/#�2�P'���v"Zym8�mӶD�e����(�&���+*+�U�y������z���'0�cO��-�D����eK%h���kh}v�X�O�|V�\.#���}Q�t�K�/-�4
�l�����a�Ɩ0]9B ��x�U�X���uP�b*���6���\b��l�gu�p�QG�5cׁ -��+йKW���<4�"��] 	�b�;c��`�!��,�I'����y���ɧf��5?�^¤���􍷌��[��������p���51��'�7�`�=�'6��֯߈Ɔ 
�;��,@��P�Mi�K"�]iL2�M�EjRI8�!e��o��*�a�Y��4�H�i1#h��Yf����j�#�z�;���0�-�;j�s_��B���y(�n={�T�)�]���P@-�@Ɍ¨H!��� �3t!�/�`���]��.���WW%��v�s�cI����sLR��p���3(��TP7*5ǌ!%A���_K�E&C8�@�YC�={�!��SX X� G#f+�|�Е��ό#��H�a,AwɈ|�	L��I&+l&�86�#!�wĨ� Gϕo����x�ba��.v,k��wn��&���C�\Z�ND����+���h�� >Z�FC���xmb�D��핮%^W&/��eG����k��d��Ⴏ��hm��!��!���Az }at����2p�s#����]�=KJF�5��I��俠�D�Y�����8,��scά��}zx�������,0����e�G�LNg.d����O�>n܄3֮�y��j�Ζ;7:�u��niKk*k���������B���`6���s���*�ʝ��e���#�k��Q)Ĺ�����5�zn�A����3�Υ�x^���V42�漘�(9��(%���LT��8k��bT$�*�}�AW)�]�LD�v{&)2�l��J�k�$ۘ=�i�ҏY[�r>�y2��U9�q�T�b�Ç���c�Z55)0�"�"�uʭ^t�e�J&h����J�v(�;-U�8�(��M*�#��E�-���U�ˇ�3���,�.�f�Ģ����ɱ�3��I�|v��9���yՁRNpB�"Z>H����b,��e2��u���b�'����M\�a��g���)>Gl�ةdF�)?L~���	(�'�}Axϼ���E�3W�-|Β�tM�G�J�p�U0�?����~~a1"�V�#^xy��t�04���p�<<c@�ƛqư0��ѱ��ޘ��x{��h��a)l+U�¶�۳���R�� Q66��&"��T�	v� Ϛ<ь$��VyLޗ�Q�u㮱��W��h�ދM[�b�w�bޛ��C���ȚD��lnF,܌��I�O@7�޽�n֚5?	��neF3�if�9�P+���1l2���=�!����CU��i���2G���-c����J"����M�|�^&s���V[U�F��g`7�X[#�$��i{�5M�Cs}=ʺtG�dF�9F2�Et����D��`�hP�o|F����˓bgvJb�E``"�LO����ܙ�}	����j�ui�"�p�}�68\�h۾͑�� ��`B���"X(HDn;�Q������b!���#5���;�Ս>� !�>#Enl� M纠_��m��������ѶkO��hh��!��pP:/;2	8f	�ڵŮ��:DF6M���q_�o��d�i��'>�͙�?������?m-y��%#Vm�ut�&`sfn�8l`��'��y�]����秬VkwΆ�
W��50�t0��6U�\_	V&���![�+�����}���~����B?0��ռ��k/t@���K�l^��(K9�����<�W�Xw&��hz����߭^�%���mf�I0[���"�fT���l�Q��&K|5[R�{�r�J K�S׌}��H|ڬ��#�f�vZe��F0~�8�r)�J�������Bt63A(☗UT�\V.<�I�W����߫Q��pD�X�i�Lqҍ������x�b	�ܘ�3�>UQyp��p2��}��j�P�v��N;���Ҙh0P��U�y�ڽ��[E�}����}��Sئ��ZޫMyx�������A:��|�e�$b��н[O�����+�p��c9J��d����4-�����Pt�󋊥�u�op�r��_LV(�s��Ov��oIm���F&��8�f`d@/.ȗv�5�F`���f�A��z�o��Ǟ@��r�.f0��\���i3�Vܤ��S'�PX�F���0�a����x?o�O>�2��X���4�ҕ:�2�I�Ł��S�B��q
���`F�j=fpE<�G�=��b�ۯ	�w�Cq�Eg�w��_����'[�|��4�n;�����;���B+v5V�ًo����xP��P����$���,D�6���M���� ���L8Ԭ���J$(�i�F�mN�գ�[x�W�EZ�j��v�LJ�F�����ET���WW���eE�� G%ѤfΖ�n�	f��(T�.H��`P��ť�2桔3�ڿz��}m�[ś�~|��@ �; ��G]����wj/���=�I9o�3V+��Բ�K&`�`N:�H��!��*��b�l��@�;���m���as(�^&�@2���i3�� ����0_� �ITv9�]���������J�����Z��#�E�H'c�T�A_�|��ƈg)(AMm���8�6DC�M�Lp�u�^4y��Wl�_��?����Z��K���b�#��-eq"�$��H������q��X��O��VKw*�P�xc���1��4��Du֧����4����]���H]�ZK������	ZV�:��iV��>v��x:�3�kl�n�� �'�CW����d���{�s�~๹��	�g,-��)F�R%�
u`@���tA�漲�:�I�j���x8��O��^__'Tj����{����eK�4��Sl���C`Z\dM�"���?��6*���p�V%U�X=�j���fJ����/J�r����� 0�ה_c���9�    IDAT��N��]{Dq����>KP�8m]2{�*�-VVv=h������d[��e�����̞@��<��3�"���q�TJ�f�{�$L�����%��C:L" BQ ��T@���Q�;� ϘqcE�4��4,iz� '(nΜ9�Dq����X��W�"��2ҦL�H�H�Af
������q�ЭKgL{.��<\t�Ew�L�g*.�d���4%]�"n� .}��B��o�)��4�mI!�u��7܊����aK��1u����
]�0�X��fa^���f#�2��0�ˉ��ţ�nx*3ω3)�������=�4�zlX�=��=��#�t�t��U`���(aV��DRf�l1��v�))D:��co����-������e����(F�yk��"�.��d����y&)�{2��(ʘ e�5�#	+WF�M[ �D"�Y4��ʇ�O`?�k�	~=���������O!��bH��s�^p..��\|pO9�������o�������"�1��?��^�K�xb!��2K$SJE1c@ii;�V75�d3�X�4��wI��0��v��+q���]�"|���0���`0Y1p�1h��y�N�إ0��Ɂh$ �ÆX�n�����-]?>�Ԙ�s����>��p
�;����:_�dn�N+�k�B��
H�PԮ_3��y>N;}8���8=Ű�
`49Ė�ϜP��A�j���m��a��6�{e.��<q׫on��j�G�/�{�}�-O�_�*�>�������۠�f۶��?l����_N��h�/)����/A�` 3��������w�i��3�k7fyz��/�d�Ye.Xsy�|/,U����_U���[�ŵ86e��,�����\��:�9�它�n��d&�z��$�>�>Y^:ϕ�9��}`Po�����A]s���%(44	��l�ɃD�"%	��������� �
�dV�~f�>�6B�<Ĝ5\��U�߻w� ������Xl����ү�����`EPXAA��BO��=k�6mJd��ʝB��D4<)r<��
f��
O�Z�T-�Y����:�l�$jj�a�&:�\�1kHÊ*�s&#P�#G]!����
��q�:	�쎰j'������h]M�#5��3�6���V��@����͓�S�E��r#d2����?���k�nq�:m�i�E�~�m�J���KWb�}o��y=���px���aiS2�[�9#X!Y�47`���[E&��o�|'�t�9���f���;.�h�t�(�Hy��
LŢ��p9��vP9.���pT?�VS�����6l����$�@�Y��Lf ���#�LZ6bv?J۵Gc("kc��A��$�d�ԾO=<��~_� ��������A}�[nG�dG4�J �9�	�GVc��j<�ģظ~-�xhʺw�5@��|�9o.�[ޓ�)+}v}�͓�D����A(+�(�x>'���`(�ͅ�v���d̊][����׺/)Ъ֪B�mw5?7!�Մ�m[pɈ�1~�H���&,_�n��R�ݻ�}>[�5��q��C<A�GX��PcB�h0H�M����z��q���Ear�ϤMP��x��� &����6m��/�ڌ��L��<��S�o
�YϠ�mGI�T-�<��u�1c�d��wO�(��K/>���ʏ��{ޚ�-f=3AJ�效�x$��� i��eB�ne��3(��mkA^N:��m�Ihg�������S-k��C�%��:�x��X����={���oø����k/�g���?���Ç��[.u�m�/U���@,�Ӟ�n3&>9��Þ��̉�0��^���_���x��?m�:rGuӠ��S�(l�}u~�ld�G���oi�g2�	�oX��6��yê%��/7�����(7V�t$�Dt����i�V�ro�`�U���<7��3�����$�N�_kI���۪���h��7��r���׳wn#�������>r�m]� 4,~�9P�[�V'X�35��H�!�X�s��g[�Y�gnB��,3��i�tcgv&��s3�^��t*��ݵ9r�pKO9�T�e�/hh���- 
H�D&+�B��Ӭ��σmx�m�c�<���/�*��x�<9S��p���LUO��/�p8q���r�7�i�Z9b�p�_�3[�.��qsg%A�q� �sy��X�vءb�z��YJS��M"�9��v�Y�#��p�M����f�Z�۰^ާ2d�DM*�e���~�Zl���*߸��l�"����'�}��[�`�9�`���5^��J�N��?[����01�{Md��IO3�I"�M��q�)��A��������Y��T�W`���0g�p��#�6#n���FA�ǐ���I�q��p�e�ổ����[�ن`(�T��H�\�	Q��⬦hg�3���������K��P�͜��F�[��MQG��P���ߌ����y��=����f�zL{�q��6D"q$ci8]y�bhȰ2 n³O�D���q�:IdvO�����o`�{�F���x�3�لPc�N���*��w����n�_���u>����%YI%3!ζsv����|��C�9�� �d7jm�[4�ہ��>Ķ߷�kF�n3I@o�7�=��3q��q嵣�k_�JD�j}D��ba$���X(��y ;9�Ri���0���F�bB"����`��p��0�ޱ�o�X��b<��t=��5�A,Z�f>��+�|�K�&`/�+�x�!S5{p�9�/��eб�_|�	��1�{v㚱�0��+����/�K��l�M�)
���7�¨�N�k�a�f��ph�~0�I���J�Ǟ��;��\:I8q&�-e�0�kqx�>����X������՘8y"l.
ږ������xt�s(*l�P0& a�)�6 ��h���֭��ag��a@�~M�"����������S��O�n�QuFcs� �����4��0�T��J�c�T�����d̷�~�9�oz��t�tɦ�լ�1�LT��Uk��5�H��F͗�\��
��wɃ�u�@���Ճ�-C��wfƬ����!�=�R�Ǯ~�-�����;7-L�?y-d��U�;0	��A�1�
_"*� ��舻�׮fNV�l��l��Ue0W�Y�Z.N%_����nFa� ����m�`���*I���h��B�xΏ�l/��%7�%P����F���z�q&��#��%�+����.��?� �˙�n�2���*��H[ň`4Ғ�p^,�������������y�b1t�2����n��<Y��Α�:�H��P��#y���}�p���ٻ�&�̷x<pZ8DJ�?�u��/3���V-{&�q.��
� p����fW}�Z���xM�h������9��[[��	�x����ٌ89��AA4m��L�3+1!�S()�,��{'�{�
�Y���.]���ISp�mcQ����q�	��\�R�Z�~��{�H$BX��RL�s8�`̜����@ƞ��x���8�Q3�4���K.F�׍o��5?�(��]��Uu���/��n�p��I*�f���=�4�q�.C�W%�	M�a����n�oxe��H-R)��v�]��O43RQ	(��k��!�`��������"x����u�/n�&H�v�[�>�77����#3�A���^��"���|y��YX���h_���8�i��S�W����G1g�f­�u���V(������I���*�~�y|��BthW�ں��8�����������^8�mߋT�$ M� ��c���8��cQY�I֬��G<�D~a��6mނE�{� FjI~�!\[�Y�A��]p�9Ñ���_���q�p�'�ۦ�O��H]x�W`�x�DQڶ�}��b��L���4���w����9a����z�-��-EMC=f�{_�X��_}-L�|	j#��]i|��p�8�oOL�g
��ۅ�n�a���sν\:
fg!")��|��.0Y���8P�o�n��r���#�?_�X��?�M�~E���҈{�8pݍ�P\���*D�u��2�-u���w�ɰ�}���u(_߱������Xܐ�6�6��w�����|�����
�������N��8ƕ'���st@8��_[ ��!��웬�'N�2l��+�X,]sYnp�l]������C�}b�a�K`�����W������״����S����Z����Nrix��C?���뀬����V��\�[mb�}]��^K�a@�/�J{����FD':Ac���Hs���m�ۨ�{vV��r��zFi����=d� ����Jd��
�U��$�2�^$R�a���W��#����jz:����LК2�I���\�������q��dV��D���[�3������;T�x��]+:cԕ#���:W�?�Q$(�WM�h���|-�V<ܔh"�*��SO`�1iҽ�����h�t��a�:�o�Q�A�.|OF}����Q�#E�R N��D�p%��n5��y0[��X��ki����s�;O6j�R���N�S�����X��Z�w�?�������c�XBP�^���޽�a���h��F�N��M�g�}�9��� �ʺ��@C|Bs�=6|��a��V�`����3��nD�`­�`O])�]�62)�-Rݍ�<���jkpť�χ���1 ��	���`u��u#��H���h,	��@P
]&<���_�����a��m��L���c�Kb��W"�ǜ�s��v�a3�1���p�yg ���D�PT�:�Ǹ�����PԦ�t;B�$�v���1�EI��GQ��B2Ҍ�G]���o����5!�2"���$'��D�r7E���C$�����X&���[4��A,�����0�pY�%�ųO<�n�e;�:TW�B���Em�1��Q^yοd$�؎SF
4�	�1쌓��c����^h�!����1��Eϙ_ �1%}�&�~�^\v�y���0���y�F��w�t�b&N9��7��������оc7"IQ�c'�B�t�=9��Z\}ɥ�?�pI��j��𡠸��_�yo��O�,C�bE�~yy���hn�Gۢ|4��G��];wƴ��F��T������������f��'
8�@��B��ކ�7\��/;O=�*�uV,���)s%em��ܗ���1��Wѱ� ��t��HB�O��f$�#Q�Qs~S&L��qNi2�8���`*��N&��x�o�qL�i��(
KK`0Q�X�(�r����>eʔ�K�Z�8��BZ)k�AMU�hB�q8Z�ٹ!�k�¡�tm�ɟa��0��*;kf�W-����K��������<0@K+5뜦���n�[rn�-{=j�q)���QEn?�8trDQʗ��͙�0m8Ѕ=jT�n��pE�)�*��Th�Ŗc%�j���^�I{t�x�B+#@<��Rg�V*]���9#_BI&EK������F�N��h�"ټx�Ts�3�ev� �-]���>��M7��eN������(�"��QJ�۷��4�SEe'D"a�S@�2�G���͔R�"˩��D��*{�V�\!�[���EP�����}Ol�����$U���{edС}'A���ˮ��-/������ݤ�ŕ��&�C���9u��۾��v��8��c1�G��\p��~����ʫ��K@�͛v�e"�L߄h\6A�ـaCO��G�uW^�Q�_�����Y�e��5����)G��@T��&��]3�J
ݘ�`6�Y�=�U
���1�ХWo��p>��x+܄���/�qfN�SQ�y��G�V�!}���>X�W��@��!?;!"��#��,�(�)?ґ}8��S1���(.)Ͼ���X���%����TR�-�JY�	ģ��(+�QCŦ_��'��s�:]�k�,��DS$.(�$)�F��X��Z#��H��EA���;�ބK.<��(�y�͉oX�p(j�	�hqX��5erY��I�#b�OP2#6�-����A��ګ��&�V+�#2Tūه�<&�������@4����������q��G���ՋfH�fd�X�I4��Ǎ�]����7�$�ﮝ�EU�b��@^a)j�|0�]��gb�Q\�ˆT8�;Ǎ��qפ'��G*��s�6L�~/.1s�}�Y��AAI'A���fB汛i�õ���!ìGE�6m��1��/��c���QS�f�&x��D<�� 鳁�t*� ��a_�T�t_���+0��s���ݸt��o�	���0ռ0ZmHѥ�x�f �G�co�G�!c���c��[`Ϸ���#��ካ�E4aE8���^$���P���a7Y�=dp$����PpGB���Su�d]�Mf�Y6�I��P�����`�j��qG��[��ɓO_���'�Y����ټq��ik٘��
78��T@W�8=W��8�Ti��~` ��`��Js�OI����}K�j�m���s������N4���Sc
%h�zk����f����j�_gK�(���9�U�cң�R�ь��s"�UoUړ��`�V�l�f%:������b����Ɏ�:��LN'���+��j���sE\y�8�3��&��wu�8��I$�}(	7saP*�<�sV K�4ȯk��ʎ���r	X@�R�����`��Q3���j!��ILHӋ�x��:���KeA�=U�hRXP���j�5i2�;�a�}�7�Ā@'&�9�r���Vf��7�"	b+8չ�~ݨ1Ta��i\:�R��>=k&�+*�{�o8h�`<��su�u�����할a�m��&o�H;#��K/B�6�g�|��2^9�
���B���N<4�iX� 6����2��<BI���:��Z��k�c�t��|���8�,^�#RFŵ���0����!$C~�j��d3�-o�~�p��1���R���p1|��Ddg{2+lVdL��oB,P�S�93�N�o�7�����#e��K�8�묈ǸN-��f�?���pvs;7��QW���� .�~^�	g��"Ē��4�!��$ד�i,�C*@�.��$��۳S���}�RAڝ6�}���|�*���)�ij���U��Oh�"b�Y�d:)�x	蜹s�ZDD�밢��
�:�-FXG�>=еs9:wꀚ�쭮�7?�E�?�����6J��"�+��7��0I����̝jhw�k��.D~I;�b)��8Pk��o��$Z ��:i�7��j�
���W���}?�N46G��[���i����t�#�oD�ׅL<�����h��tb�[�~����cæ-X����/m�ÅXB��)�����D��F�H��{3�"��nS�ʃ�O�.l�&T���k�v��5#�����ڔ�ke45���`�Xp�S����e�/hW���8�Ne,�ǥܧ�9���ƢrV�E��+F��י�6$�p�ꑂ�rQ�քD2���,��ڛ����膻����˗>a�X�����F��g72Щ��Z�{�9g�v��.�K��tbN0ϭ�u�>�����L�t�������f=�W�����;.	F�y����:Ӓ��sxu��ߥ�pL �����V�Q*trGIw&��<t��AB��ơ�0����-�I��u(?��'i�Oə����T)e+#
�ĩB����r^���7���&4/����M���;HCZ���|Qg�v�	N+*��*���t��.	b�] �8�q$��ly��t�2)�1� x�x�	d˝�^i�Ǣt:�_I�x�d�#�׆��q���ә��.{�U�$�]	hL��N�=�z�g�.Q��H�$��RZ��x���JF���[�W�����za��	�C�������Cs (r�D���d5JBU��'Ԟ��������~M<�׭_/nm7�r+6���L�kA{��yHʘˤͨL�(υ!G�}�v�z�N���~�y쪩��YO#�����dϤ���o<Ԍh�	e�y���L��c    IDATsq±G�]��v����K��P� �2��!��f���jS�sfSƔ�M�3��0���3�lۉN]zc���d�wГ)bQ���$������N�о�7�0��߮�/�����m�DVT���p����@�ċ�eA�a��D2�g,��ON�v<�v<^`��g���_�S�Q�I��d	��#A�ԇ�=�ʹ�l�u�J!(%<C�3&���Lʜ]dR�۳^�Y����.�ٹ��}0y��s� \x�Ht���?������!1�e� ��aNb���()*�?�����]q���1�����*(���ן��T4(���}�еK��cH1�ѳW%Nv&��q6����f$ɘH ��D�ӊh�'X&z����׀��{�s� ��?�®�m4��
�N	�6���I��hTX���H'�ع�Wt����s/Fy�^x�9��L
(�H�}
|�h__�>�a >@��9�H�	�MK����>zᘓ��)���3/���KW����8�P��.�3L��H�7��(���%�I�ƽ����N�JG��Y�u�J��zs��ϼx�U�-}��ɧ-[��I	�Y*����G�+5�4���h>�2aQ��F��5^W��\�-���pps��������+c�tK]oº��g ���U�~jn���ǪZ�ɁBǧd��YVnW@���7_w+4E��l���v"%�쓳CtV�T�u��R�k�BU/������c�`E�>V�<fq�C��UҘB�!�Y���6'[��U�j�K��	�K�P���� 5��:� թ���*6���bTR�: �&���N0	��n5�LJ2"`(�X���� ��p���
TZ���ʙeRm�4�P	h�M4:��I��䢡�N$"�{m5���1�D�����Hk�F�5��;-��x\D`�T��e�'p��s����Orm]|t&�a�0Y�"�"����#CM�`.j[;,��(��17�l1(��TR*���:,]����[d�4g#Q0,5C��:7t�Q��j�kл�!8d��x������)�S8���<�T�R����d8�w�zu�҆lh��-�/B����"X,.�,9�P$%Q�~�x��h_�@*D�n��&����Ͼ»�~�ɉt��3��m*�0��F8P��Oęg���=~�-ek�Ÿ� �������0����7���g=������w�}�]�٥�=t�v+y���X���i���)�)�S4�%�F\M�����Q�bDqg)��
ɩ6y�k���4X[#�j�E��mP�q7��c��I����.�m�`�G_b�k`s���:�dEyV4V�D�_�<���WDg��2�� ����d�RQ
�GhB�Deej��"�\C:�!������p��A(�P�O9��9 ��i�xh&~۱U��R�C<i@��PFxT�k�ُt,�L2$상��^��I���Æ���b�������N��7�T�c��F�׉����5�ܽ��e�5�N�}�$3�I%��JIb��)(EJ� �H�HP����  ��N����$$�M��dz9���]�>�yy�>}�~�˹�\i3�<�y���{���Z����t�����~Ь�0;�X��w��3D2E�a��I�Ew�N+�C�H`t]5�^�Ǵ��o.G뤱H��x}�j<����3���_�ފ�0�m�z�n�������$�B������&5�t��TB@f?�c�9�C�GgzϤ	�n��m>�o	��W���G w�TY��xP5��+W��,�*tM����6��%�l�g~�*}�U����|�J����o���w��?��F��=��'��?��cp㿑?@���שs�
z׮��.����C���<t��JMw�g�(ĩ~:��ҘV��s�#�T��8X��$+�?K���U~��,���ZI�J�ܨɳ2iK�(���U'׮��0�e��@�Ñ�[��4�)T�8�W��/�9{�g�x&�2d�Ns]If�5n_S�*L&��>H���$2=R���UI
�9kN������F� �BMQ$;�]��lp|�b~#�[$�唒DC��[����tVX����X<��J9D$)����X�d	�z+>�h�5�R�ДD1�� )Ψ�K�D �ہ�|y),\���l��O>���&�̳���<���~���M�R*�4�GbhX��b1�ɓ�I�D��ν{q�)_�m������[���d���dqO{S#�H�BH��0*���G��k/�Q<̿u�w`wY�a��t���хڦ�h�iB:U@$���)��G>5������2|�+_�I'��3�~:�t��;�Î�	���h*�� g(����a+�l��S�ǘ�Q�����sσ�W�_=����C�ndrE�i8�!��,	!iº��]8������o��Mm�����-��D�QB��r�N%�sİD���tVI+3A����p��k���y��+�-'dܯ�C�ߋ=�#�c�\�/͝���M5�~��{��O~�T� �-�<,�a��AݘQ(d�H�1uR3�.>K��ÈD��x2���q�$TF�K��o�T���l�~'�:v�a fϘ�c�,�a��Q�vI,�|�x�OB(���5����q��k�F�T_��`/ʹf8��r�Ќ)��0���lܼY���1)�U��uP~���A*�������r�<b�<�*��}I\���k ���&�
�24�)��ؑ��pX�3��4�p̑q�_��������\�mh�D,]D����4tz�3(���
4MZ�����Gtey���D��Û��V!6V�L�uz&�T�,Ɂ��5ο��[���#����*!�i�`�����`V���<��6�:�)L;�D�}�s�����������[�]�s��W;�5�����a���=>Dj\I�Ld��'�����h?�,XUb�Ͱ�Uα/�r弐6H��*W����9�T W�g�W+񜦽#�#�E {>/�U�+3�
PX��^�����sJf���y���E$�=sIh��!4n��B�de����
W�j��s�A�t����j��8�<��\7*Q��HA�>mv�
��xyE���LzDCaa�
�J�Q;V��ږ�{À.���+0�Y�����V2�%�M� ��k��Z���F<E>�/7��V�TD,�Q�w�23}ϝ� F+�^�N`)���PB!�<�YAr����p�}?�eW\���}py�x�f�v�3��lu�d�H@�!&^��K�%�,Q�b.���<S*�d6��(��<"J�/�Fz>B24�c�t(.�`9n�����Ï�⍷��eW����n\��:�k`3z�Ζ����0�&�!�h�s���ގM��;��>�<�*Eb�Ҹ���P2Q�F�����i
��r����_s>~�q����{e��m� �{����`z��Č��G93�0�%ʼ�����Q��b�wo��6V�~[w�#W�!P;Ѭ�|	yέK(����`��uy�%�K+B,'S�8�t��p7�s0�
0��FC�����SE���'�>Z���#x��q��DQ�D�d����1Au� �Ӿ�+.9I8y���W��+V`��Kq�9�� ;?����2,xE��e ���q�q�_���̀�
�q�}r��8�"|��3�A�nt3ں����IS1q�T���/�ms��Nc������1y�}}A���G��OB}��`��#��#�*��B2S�{C/x�݀l,�K/��}�"�����[q��+p��0����ƅ�l�+P/Z \�D���Y�0��H�0������_ڀ�}�8�H}������Uu��NCgt!�WH�٨<'�KD�����@yYj�dGeDZ�i4�Ɔ����6�����.S�Y˟���N>���;�KC���n����O\�z�]&�i,q�(���*�de.���LqH/��LmJ`Z`�L�e�����wQd����ڭ�,`hU�����ӠR�=����g�y�*#=�P��r�@,$��r�9�}}ң��KK$���S���s��&{�pڶm;$�9\v�rY
���4�'���k�������C )�m6�9��YH�c6j���QeM�iW,܊�4KK�VTHryV7f�����&߫�T��5h>���&aUNF��D�3)	�r�bh���q��M���P�t���:Z��xjR���r�(�l%�d̚y�s%	���DM�h��T��C��(�!*_3������##���}�g�Wn����q�J:�jk��%׃�\�@ �hD���w��G��ꔖц@�Zm'�t
�}���F����`8,r|]s���B6#�B!���g��I�&໗}/��<>�������p�(�0iu O�jm�5abO?��i��}�B	;wlły���{����Mgq�7.@��D�ȑT5}�uJ�\"$d�sO;˾~*��=x�7�/_����q�M7c��Cq��.��k.��bF6[F*��^�ƂC�՗.ǲ3N�p/�?�x�ع����'~߾d�E3�e�5J��}��q�<����=����O��g�Ĺ�,�c�>����\�<����뫕�U�̙vj��a#�t2�Ä���{v��q�K/��g�(��ʫ�?��xM��X�E�UX�f����=+��>�׽bBK��*] w��Y���<�Dzp��G��ӿ*P�6H"z��y��Ko���oCu�XX�U���b���Ԅ��.8�:��/��Y�3s<3����8��Ð/�p���i,"ɬ$6:�Mf��!�mf$��5m"����8Ɗ��<��^Ay�gX��4DY譴P�J�~��_CwW�~�A�W���,Z�K/>�>`׎}��K�q��C���S�nBfct�t�N1������f,��0���3Z��g����	s�����]ӈH����É��4�N�sZ���Еqم�ā�'��څ?��&0��Q8���d��lHK'�*�jw+1+&Zn�Ĝ���4�P�0�N����m`Aebw]�I=�$ϸ"\.S٢�m�e���+V^�dv����_������2�\sͩ���6��6��J!q�����h�c��Ԕ�XQ��+YĬ���t%����HA�dv0�!&�*�S:RާR!i,tt+�xE^Rn���Xz�h���|�g���C���/Vz�T���Tմ��ܕ|����G-V�.'�Vտf���Q��h���摔9nV}:�]�N	<~�T�}��0���OL�Y��
k���l����l.�MX,�A�����NoHf2�n��n�x2�v�]z��s�E�|��y2�qM/�0Ǥ�(��-ωϡ2zC�Z���e��^��f�f�H�].�S���"6!FR�u`�O*k���;\K���z���E��,�f�.׎ֺђ0~��0��)��XK2H�B��1^���)Lt"JeC�Cz�W�<y4Iv>�$�"�"?�������`0 �IU�*���	T�5'��s��J��X��l<����6�l*�(�p�I_���g��ע ����J�)�	'�V�(�p�q�����{��3��6}�[n�!g�D{�H��rp:Ȍ����b���4w�u+v�ڋ��[����o��_��.\w�����W;Z���n�S���q�	,Yt8������MX|�A����7�r+F���Y�.��哱�tbCڷɨC)�@S���u6�]���xT	�pn��v��ۃ���]z�$;��QTᄂ���b�x?n��j����֛�ą!=w����;p罿�3/����F!:�\x9EVb�q.D}�~�3�O��֖1����={���P<�����=om�0�kj��s��̡��p��+h�*3%J�6m�D�p��g�2�]�&@#��F�3���O9M���z=�[߉�z;ww#��I��*o����PL��2
'�Z� �&6 ��Z�G�z:���.�%R���� ���gk>�|:�Cf���}Z���� h�w����W^E��&D�	a��N�����Ȟ�^�	��D�Y�,���Ɯ��A��}]�x�X�q��d�z�Syx�"�LK�Q�(�S���&�mF����I�-��',Ũ=���_>�k�ISǞ�P�C����p?xU>���J�F����#���O���5�䁧�&~����0N�W� L�Ϩp�=ʳ[�r�:*-K&^&lr���ؑ/s���EQ�3�R0���;��"�O�u�U�������]�uן��{��p8�x~Q����iU�H%S�D��DO��t��5"�?��@B���୑N� n`M�I�:�Y�
IaDI��ɬ&��,+8�a���~�r�wy�j�R���|@��\W2�
(BXQ
Ծ_EHȗ���+	K���6en s;T5�� ���9���vy2���^GP�Vҹ",V�Tw5�5�b!N�b]�rnocC�����Z5��5f2[�(����GW�@KoO��`4v��b��7�t�E�Q�l���<u�2V��R���̤��_W�?��o�3ᶴ� ���-Y�r����SI�(d���U�j��DJ����_�ؚ�]�9'jC:I�9�2C�_�����w���Ky&;L)T�Ng`��6��K2�-�fw�5g��M�a�Y�J��R!�L�_>rBoB�)ɸ�:���:��
����{�5O�|���L~r9���#��}��PV�V���}��t�K� %w�c��;���f�+/��X��!C��~4~|��X����~��iظ��q��F��><��эx�w������@JyJ��p�q���������_ށŭ$rE�?��]_�#�׍3�����f����z�a|�m{�!\��[E���e��-��2P������"X��`���RXLzt���칭ؾ3��n���<i��̂����j�j&�#�\6�E���K/B_w�'eSYv�\�l���W\��	���p(D���t&�T&�R9�C���o���v�܅��Z�5k��}��a�V�_7Z���RYR��J� Lw��y%�IKI�jG5 ͠��I0��Bp9�0�����cQXM:�U���G,�i˖�W�Ǿ�~p����Ƚ��A��|�.�m�W�Qp�a1�̳��ɧ-ī�w�WO=���~Ē���d0�i��E���0�4FI��w�at�/8��:
'�F2\��[�~�fx����8����z]b��۹�b�k1�Y8��`�Bx|:�]��=�z��bO�D��is"���Q�B��	.����'��䯝�i�C_��ʫ���B�B����f�d5#�L`��&��a��0e�,��وƁ�~p'�_�1��"W �J��ȴ�_�ʜ��c���էPY�$}��� Ǥ�.�j���4�J��/>�̕�:uQ����}��_�\.[����e|��F����~����|�Z���V�V��@��֣��NA2��բi�2������}�p2F��i=^~�
�*�r)u9V��rVllB�JӼ"ẟ����s-!�?�.p�WZF.���B�>��J�A�T5��r���kQ��8���̚W��~�T����vg%�Y��PP�ňh�a�8$ q<�n��S�do4:��#���g����C�3FE��}����^z������{;�3�m-:��OX��t��Yc�,I�RStEb��	�D��RA��e
��#�I��9���D���p!����Uz�����9��9�i��~�Y�;7g:#AZ�?V �
���~L�X�j3���������^-!m����w��.�B���>[
6��w�F�U�OB��Ȕ`�#}��e@�/��N���=t��d{�L�O����<^A�6��n�&R�����aDU�F*@����4�ע��KH�F�zt:�76�h�!�-���F�V�CCè���V&"z]	��^�3_��E���_�{���NI��~�A�ǅ�g�k�q��IF<�"儍e8�f�������F{k+�����V��_ׄtрp"��R�FA;hN��!I    IDAT�w��˟�̜�7���!�Y�6W �f%��X,��tz�I\slo�1c�D|��'ą&��Ilߺ���3��Q�2�7�� ��9�V�B=0�ʨ��������U����B�=�(��E��z���8ܞ
��S
qbo�-$���Ie��PF��H?�`	u�u|C)�I?��l�U�u�Ȩh��������x{���Άh2��"ς�:�̈́x�v�u�dM�"���ę�ᩪG�`�DF�ҩZN)��n�e5���t
��0�Nh�ζ��K8��q�9���s���?DM�(����P;�E�r���\*�xl����v�Y�=��gcL�x��7��m/��E��[�q��y�F�T�"D��C�߃R1�`p �B3��Á����5k1���dC%$�:�QͳJ[���yx�V�����gn�p �N�*#�m�;Ke�[����#����J�ɹY��y����{쪓4�3��B�o��e�9��i�=~�W>}�ѓz?�;*t��W�5k�]��xjņo���ĤWZ�����g�R�#cЊѣ�1{�!R��!U��T��Վ���W@��Q=�*=[9ԅy��LY*���>%�����oNX�֧�U����X��t�T��r$;�%��
��E�1
�(�X��5� �~~�T
O�
�� Ġ΀�jMcSכ�������צO6˼��P�Uu�&���B{F�nx��˗?y������&~����ڇ��'�n]��WO����zB��7����5��3�7��K�&���,l�y�A.�@kK�����ۃZBX&+�UU�N<V٪���#;*_[Da��.�ݼ��g"�!��B���ِ5�$����ϳf����l�t+�Ѩ0�m��w�Bȕ�(ȁ�J=�<��T��p�_7���b��V��>/z!N2Pp���H�{�"��?s��e�s�\�������%�I������M�uP[W-��E�?�ՂƆ��؛x%�9ᩮC*�V�&�f�_���6+RqX$ ���)�]�[�s���x��/��Չ4�B��T���A"��lF<8�t"�I�ƺ�G�2��j�Fww�#=�8�p��d�IȘy�.��CWH�a��D�<�/ 3�	����:|0�
����@�C �M ��TL"7ԏ���Gb�$�����W�Z_ӈx,#�k:I�v3��^�9�����H[.�M�x�O&Q�^���G5#�����ή\
�10R0�՚i�1��H`��s��X�ի�B9O�ܣ�sq|��8b�?���>P ([,`�������_�1�:ɶL�D�.4�\:*��et����^��6�KxuF������=�39���Y��P�"����ۆA��髐)�2eM�h�8��̠���dV83\'�U^� gb��s�Q�eODU�Ho��S%����dG&���8	e�<.d�?c��)��܋\&!�͵�MHJ�g��@��ˠ�Rix������E��Q�0u��.-�/J�R�-I�#����N��<�x�����_T
��[D�B�L�[(�R�a.�4�Ï��o�������3���-+V\s�����z�����B�yV�ɔ�wET��+�<�9SMX�PgT�n�8�p�s���HJzO�'�L���נL#!`�p%i���Û�r�R�n56'�����vԮ�N�s����fd^.jF�D�5G*��
<.$1USpD��+6�$0�S(�����Z�H���b�d���v����b��jv;�_ñ8��0q��Tg׾�ں��W����/?U��_�ׯ����G��λ7VW�Of��X
v�Ww�<05���V(�H��@�9�ED�Q�X��[�hp �Und�q4�nĔ&�F��\��T�L ���-�����X!4f�D8G���KA�T��=�A�δj�=yn6&���7ϓ{������
��hC��u�!�d˰9�x��a�����%X�q�/@}x�x��4�@yS�2�LJ�De�E"LE%�H"ݘcl�'�S��X���f@�"�j�����q˿�'�huإң�%�&�A�
Ya�S`g������ �N-����&J4_m�ˬz�C�r8]��:m�R���q���8b�i��Er��#bD��d���V����G4�	�\*	S�$�cޜ�2?�e?&�	x|na��uv�5���t��d���J�q�����_nZ�*ѣ������`ӎ=���-е��T&5r�s��5�!�	��P���}����E�.Z��a�����26��TI�Ľj�10؍I[Q[@���鴴Jx?�N�4K��;0��f��x� �Ib��RP1�uȊ��S�e�r!�$g�as�PW-�|�4�bp1�	���8Z��hQ!��`ң���|�D����{�f6TMm���^�C|�y�����kE����b`�>����Eo>�d��@r������j8��m�%Z��-�5�64"M M�^� K�w����@.��fFm�/	'Go��!<N=�ͩ��f:L��h��Lj�!!�\@SC-��a6�D`�������.������
1�1�-,
�D�`(�Em����D�t
�xR<�[Oge�8=>1��I^��s��D	W�}��]#���we;�㵌95/��`I_Ln�Z�O���+�>c�/�;��s�_��rپb�5�]��{^�����o��9���K�,V:�����r���Й,�X*�3l���﷙�:�H�#��D&«ڨ��dg�[�rO�ʃ��vɁ� C�E%��E�2�Sɘ��j�;�V,a�oR���E ������ő+%��*v飃$:�)mr-��F��$�/�C��8�f��h�`Ea���F�h\��~܄��H۾��xeR�.����-7]���f�?���yg����W���{���>�bvX���He��r��Z�+��#l�
ܮb|�L3gL��i��`֗�Xr��3{&vnێ�k֋�O<!�8~F>_�;�8�=����5$CX�F�	�hb8�o�Ǐ�@��1� ����F0$���p�Q�dC������0��y?i^{�ر�C�gI�9BxVA�(j��9��g���8Me<B��ʹF	�)��gOB{��j��!E775)��H����PM�@��P���Y9�g�݂o]x�}�u���_��0$���W]'���W}�Z��d�G�-����iSp����3�j;W�HX��φ	��O�s���>������l��%;�	���^�����nV2��H���z�2�]][���ނ~�(��#ba�p��F������p��1O���3(�3� ��J�����/�W����:1a���u������3�����Npe�?��Z*���1��wa���Mv^aQ`6�q��3q��G���B��?�/�{������a��N�����e,��a8.5��sCG~O&�&9_,V#��$�.'��1��NZ��g ���X˨�hjlFW{'|?�k�?8g���c�"��}_�nk���"��A�+��p�|�Ri��ݍٳg��$�Q��X�lٶ�]��Y�%$b�U0��%�����G,�"rw�M��L*���f�C��'W>��7nAss�\�~mUB�!�}.|�硐K������ol�/�rv���k��-�G��p��P���_>~)/Z�x���a��u�\Gc���j���݃'~�4zz{�HA�*��XPx�|�9pX��PDoo7�Z����?�/PC�u���)�{�E��e|(��Ũ�\5.&L�f��`�
�����!�A�VS9���m�l��w�s�7������n[�b��5k����xZ���]����"�0�B�P��t,[��r��+��V�!�?4�
�޺�B�lo(��e�?[̧�ϥ�2���� a5/��P��֚���3ǁ(�O!Vp���3-*f�n�:���������["K���ɨ��$V<x�CU�3*PAI�/���̝0:�چ�\�I�͈+�qq�m�������'��k����v�'�Rj�d2$���GKO<�ڕ�d�?̵�{��go���7K���]U[*E���L�RY�(��HW�+e,V�x�}	��NG$؋�-�8��y�:����@���N�
��.q��^�a6���vߴ�RI�B7D�I��Ҹ&��������>���$'*D�U��}�%x���a�M�:}�0l�^�!��<�")�m��3ټ�<+ҢNi�S�3�z�2mZ,I@c��B���~�Bg�NKN�g!Ȥ2�`���5+aa�d�bd��Xk+q���S��nWl�DB*/��f�������c�e�P�Ј��$A�7����Gֿ�풃���W^z	8`���1)5[��ޱI*?~v«o��!j���,������̯���OE>���n��P?��g��}'�aT�v����-܏��DP�$N���k0i|���)ek�䉁�6'�	U�,.?���J��+��,��<���&a�՗�\��5�|Q�.���d��\�Qq(�wlk���eW�6l���G?��s'�d-��B��C�fC$�DӘ&|����p��c�7�)
*A��T�3�fs!Oݑ�B"	�Rk!�bB�=_���@���<N� 7DL��a��8�nXMI����aX��V(I��Ő��}1��"U6�����hM�@�B!9GE��T�u���I$Q L^[%�D	ۇCC��IY��!��on�C��d*�X�g��b�"&�3";L(�&�0�9	¶�hAo�F��>��b����|^"�ׅD4��*?���0~L3�0Q�<��L�j��d�����S��� o�Z��`H�xT\ �y���s�D���[�ף��C�p�}�y��}]���'?E$�$��]�2�".��Lƻ�(tlu���T7�6=ؓ�Ll�ݐ����]���E����G@�]s͍S׭����=+�u�V��D�H'�|�����j-�r�r:�)����^�+����\.&�����7i��M�,=�kwO�k��Ϩ��惠8��3b�5�Cu�*��Y	���|wVA��e^a���k��1��y��s� ��_���Ӧ)"��yP�h<x��Y1P�nhxi��u:XE��$#Qu5U�������E�'D�̐�2	/�y!W�����WC�(�P�7o��L���Pv���;`��D���t�!�W���iӥ�y�}��M��ԍ�7�q��g�s���C�ۀΟ?�W,^�ẟD㙩����	���\i�T�T��|V�� �$"X��q�ڲ�#q������O6n��mm8��%X�v-v�ܩ�)�|%[���
��'̮�!0�&���#h�3�SQ(`�I�;Q�nB��Ν��0 Θ=U�u8�s�p��#�c�����-�tG;\�!91�s����H���2}�#a9���p��`�E'��u���P��i��l~�r�9?'?7L^/�]�_g"���%���J��sh�BQ�C�'M�5ŀ�ր/P-A��y���[���7Dʜh0��k�<n��	����.A�Xx�6�'���v`���x�ױz�:�\nD�1yVL�Hf�G�8p������h�+(z��u��h=
� ^|�%̗�J��`��H�c��+_9Z�i�G#���Ԋ6?���`��M�[O� VF
�#���,��K�����\�XB���&,�Q�ڻ��b2i����, ��/��N��w�~9r#�e�U�
_��)J�>��? �KBn0Y�]$��:�|^���=0)&�ˑG
BQ����M	am_�^�E�km6��-�H�k��`5ڑ����&��T�tFF.C�� �vD�qJ�:�	z�V�N&E\[|^l�����x%e�սـt2*/�d&}�|~DA��mj�G�Q�S�Y�D�D0a�ړ|V�Lt�mV�$D�D�@��(]�dg����3I�leJ"�#�Y�QF76�c�@�6[�_Ŀ�h��i�:�"0SWS��� 2�Ƶ4���D�--ryX�s-� )6�H
��u�D��;�w�s&"l��=>�b	$h�ku��4,��D���}2��������SM��s����:�������?�M�ӎt:M�gS�����NW*�J�r���j\�+���r�P,�r��J���������ydd�1���[o��{�y��v�h���{�g aϚ�֢�� �ROT��W��,��� :;���e�=w�����^��\F	<������+LHB�Rɹe3���72�බ��>���\�<_�׊'{\�;y �����V��aȃ��/�is���!F4Ö-[Ѿ�SfR��~�շж����_��008,	�1K�EsS�z�񛧟��6��U2���u�W/{���V�+�9_�Wޜp����h�?I�t��,�t^��I ��(�u�(ƹ�門��q��Xr�|t�ۅ���۶m��O7b�������S��Q�^��N&)�c8Mk'(��I�[�{�=4�7(豿_*�u	�3������,��������?����Hg�vWcTS��}��Hbw{����2�M���VW�I�t�^|8>��CDCCRmp�Nf�M�9��r�(���x��'���Z�8�n�������MǞ����ksܸq�����>���U0T��	���n6�d���}1I}D~x�L%��ۼ��:P2s�D<*�ntC#R����l����zԙ��F��� m$�m�ҩ���>�œ��F��'*^*�2��%9d�h�IXR1A78��q<N���& za1�bQ,V�in��9�ʽkl$���jՂ�`�wE�P�p@bY)�v�T��Y��`�������aU��tR�m=��x�E$��۫&8�"Z~�"z�;`��`�;��@���b����;(�ഛA{�d,(d�Mþ��dR���vz�UI˂�ހO�m.%���Ӈx����������2ii�����"!d��E��@�"�i0a�@Y�̝3��Wָ�2�
��5XWS�|� {I*j��:�	�]��I�TŖN�wV�L.��2!
����C�(��ҁ�~a"R�l�XP�E��,I'��.yn�p�M"����D'��1�����S.�[\UU &�J�9�J<�	�&"�� �����.	��)�K4j��vX��n�"C��.��H0��6'�=}�7�������<�K@���EY3EV��_l�w"Mo�l�������G��������yL��Q��)@W2I� ]�RN ��ٿF
�XE�/�KI?��E�cΌ�d!ǣ
����nf�ғ4(�vnr��za���4+g-����5�Ȍ��
�5׮���'��7�_r�g���r0k�=��:�a�^�Q'߷��S��_U+��=��r��Cq����c�������/�=�ӊB1�q��o�p�w����_��
��۽��=CñSBѴ�@kK�M�1�ѩ�R�R33�4�Y�W����,_v�=6�u�K.��?���WI���D:d�h���D:)����ISS���$���C�+����@'��C�)n>~��$�o��#�0����`�Øh��N���ø	S��Ï��;��	�Ӈ|��ꔋ�\��9�~�hP�G2Nw,2����xs��:�7t��T���B�ȝ�X���~��N�w~�#&9����ُ��ߠ�p����V<�٦"���$ٔ	cgO�T�����z"BAA �is��J���J�?_��=z^'�n"���F���Q��\&/�/��c�qȦSBc 䄄��V�V%1ϓ�F�6�y�ʊ�&OL�X)��F�K��ܫEa73����DQ�&Dr"�<�ʆ���YC�a�C�X�~x�tvt���V<*����_�݂�y�C�A�Ln���&��[OL��;;���. �A�S�n���(�I&_t�#�p¸f�m�[?b +[f�©1�e�&���B�5����Q���R��U6{�D,� 9�n�����0s`��Ą�������d&�$SQ0qb� ,4	�=��*?��D�iykC$�ӥރϗ��\th�$�z��9�@�@,��Z��,�`fT(�HC3Qͦ����A��    IDAT����t����0�MJ�ʜz��ߥMj��sV���3�7[0|��dF�-1N�8o������ry� W��N��s9��,M[v�IP��Â��&}X��&�.�������'-�G���_��¿�{�o����[��|�l�6�ql��\��9�$�e<E�aO[z���D��b��cF*�Ic�J H%�hooGpP�s��#@���E&=l��U�;����
��|kQfC����!��~� 8ߜ/�1<8�ݻ��G2u�cV,�YF&�Fw_�C�Q�ԮohB��]��s�#�E6_@8��7I�WE���O�a�y$����Oo8b���g��ϟu���z�ݏ��-�K:3L6�t!�A����$�pqs��Kp[͘6y"�0��U8����E"6�=����hƯ�kI�x�y�5X�2��;��mh((��I �ۤKW����tf�<��|1�R&���!�Ε��h�F똉2bt���W�s/������{�uW'l��mj�M� uj @翮v����`��q$�H3��J9OT�(,�8eؠ&�A���rQ���@(6D��\;��:�Ð=��F����+�^T?�ʛA9ǃK���Ȕbb�_���a�sz�1q֙��U�C�O���<Dy��g"�������J�љr6�C5�Oi#�r����c�#i��7�UFYa�v�^�d^5I�LT�kb�1
�)H2��KR]W+r��pD��!��'Jq��$�EZ�uau��Ei����K�ߛ��s�oA��U�D�Q%���)/�����/�*[�l�q�l��ۇh(����%��k�ط�
�u���p�qG��G2Bb�l<i%p����,F	\�!�5�m����D�H*�D>��� �+��X\M�����8a�ʐFd�iL��*�����Q��M�<U�L8���Urp��o�Z�m|Nrp���s��|�
\����۫T���W���j$
U������_��9�s{�]�{����\�=�s`��D3������`:��#�4�U�(lÿ3�Ϥ9m�{�v�"][wwbOG'F�k-茺Ho׺��F?|�i�߿��S���T@�/�7�����`�ق�J�O})��P��|*�r���2�Vts
�M�*�_�$E����B��C�d8~���V�i�)�n��l>��!��=�]�C����ϳ��ޓ�*����Cz�9̘9睷\z���y[���߈��aF��z�=���XLF�@�$�<��00�����F:����&'�	~Nf�0���Ȧc��:�+{�晓[�iv�%߽�~��K��m��d���U:'��Ƚ��O9��a��౛�����aޜ����+�Qd���jsү�f|�4< ����� є�P��(�QVRYU�X��pb ��U�FL&L�<Y�7�u�>��]#��!�*c<�Y��3�J0%r��a�S�-/��.��Ǎ�����T�z	��c��ͤ�K^�V��ט�D��`;E#�1)�:RbK�
�߅pI�d%!�:�=�8q��5*k�?�5F��0�ȟ	�/��c	��H��Ϯ���
J�����~���FY�m6��^S�� L�-��R�2PH�,�qU���ʔ���&q�P�~��2�T)���k�J��dR
{�M�g��ׂ����2�k:亰j�~Ir$�Ҝ՞�& ?�`��̨����4��2"٫�k���BZ,���w�����@J��$���2�c��$�y�3V�S��C�Ԍ���n5�b�fK�:'��+�|۷n��@�T���y���+�$���"�Q�HDa%>Z��$�i1F�b�gV�AM�p1��}$��э�n��Ѯ�_�,�`�g[�����C�26�{�����EÄ��-I��2�"�GEX�6�1����>�#�$K�����]�`�mۆu���as����y�u4�N!����$�U��r���HB��PK��}L@�Eā>�o�5.�d�F^5�=��j�y�vރ��[J���_q�+�-;9��U�Q}�\v~���oxo}ۥټ��k��0��	C��B�,���n'IBS�S7<�	*�����+��I �)59n2B,ɈP�6"4�Ϫ�j��׭�|i��)ՠ�P�S���ob5	���^z����uI�_`X�)Y�� !c~�ԩhhT��۷������u�ln 2W��cq��VKB%��<��H'#�����g����V���~�Q�Y��/�.��p"'�iT��1A���>�*��)/���7p�� Ǝk�E睃��=8���`t}֯�@���N_���/����c٠:=&M�$I,-���1P��0#7���[�sV���^�N`ynF
�L�2E6��v��$��uk�����/���2:��[3�!,J��*�M�lY���!XM����*�ʁOkS9 y��zU���I�]&�Z�a`�*t���Ow��GX�C�Ǐ���ە8��=��r_ Y�oM�����i[2��V�v֭��r�)����5hh	��!��x�%�m��=5�I	�yIP2i�Ak&�`l#��D▱\�>;�yV�21#{�^&y��3�*�bQ�ϦH_D�؆���c"M䆯!�1�g�Z�b�H<q��dE� �X���ƷJ�)�`��M�|^^OZ��d�'��0@y����0��/U<Q$޳�={%�;i
n�ѝ����ko���7�@�\�x��#b��s�ګ���c/B��r��"Q��K
�j8I��7ǌLyT��vw�b�2�"��F�2��eZ��M���98��G�	�������E��ȵ�XW/��*�Ӌ.�C׾n�-&�mA����z�޳���Ȃ:�D�d��X�)1��C=T$����ׯG}}�T�E�U*$@C��1K>S"{�+\S��A�~��(jA!Q|_������ƈy�
�R���q8|5��k��X��Hdo.�\y���{��sN�g�9�?*�r���gW|���{�����_��p_(�T��񩨈�ڶ	AF�6p<���*읓)s���+JlL ��/*q>@�sFUEt�b���@�.�_��
������Z`�d�r��MȦY]B�<��4Bg��)�j63���4f7_;���r�ò�x`39b����"�/$���憪�V�|⚙���
��[�Y��g^��l󎍦rR���:�z�]d�����#	E���^�b�f|�����|Д�8��Ӱy�&tt�,���o�����_�=Q�H���h�:ܼ���H8,=7?*L��>nXV�|}�;4�g�?�/�3g�LX�}��R���h3��<���ػo���.�!�hїP�w�m�c�����D����
�ʬF*^�	ټJ�����ƀ�)ש�F&{$�������L��d3u k�9�@Z���w�.U��bh#��x�Z�����7_�����J�{�S�L������a�k)�D"]��|	�H����H@)��u{��Ҋ�]{Dc��"�'�?�KQ�1-Q�c(�}$��,j�Uh=Z`Z^;��:EB�D�����d�$"'�+�qA����س�]֡�*A*C��L�1���z�[2��ѽ��&�e��=m2nF�k'�V�/(�b�D�6�pȣ���͜9S�I��!�U�"Q�)���{��)_�:b�4�tv���ϐ�Ʃ���N;�d6{^����DU�}_�-�!�������s�sOg���Z�?�{��y�{g�^���Ŋ��A�~�݂x"��qP�2�-��t�&�G$ƖcQ
s�/J9c�dДs�B�4�4T��(�J&欖��L¹_(H�qF�OXTѨF#`�߀����?��_YN-
ro�1"���Պ��V �^2k��OT�HT��9N�~r[�NX�Q��pO����#�GSS���zz��o@�z$��	������o�?���z{�l���.�h�r%�3��fNc��z�)%�0�U/Qg��M
Ŭ���*�����Ѡ���p��b]H��aW�i�*nn����j���ܭ�w$͐��*=MO^��*���{21Ȉc���yN�؄VT�T�PU�TA�BQA�Hf���V,II�c���5��JI�|��L���Y����?���N�?��fQ�����e��^{�k���F��՜Ε���M!�~�pB�t���x8��OR�-����]�hh �ݝ8��31al�}�]��yh�رo��\|-��^.7�6k� ΀� FaF����C� �/4n@<���G�)S���L?h� �ׯ�_^{U����⽏?Żk6�[�,�Z�.�C|�k��"��>@��(s�J4������$����*���;~��nk4�Dw6�"�3=��&	B���t	%��H�N��OF��z��\	bTt���E�]}��h!Z][#UNK�(|����X�$Ty��� "=�bN JB�R�� �Í�1�s�nA[4Q&&D�RIz=h����X�o��|>&���m�ā�̙,j��?����OZ`��0y=zv��-ϕ����3ߊ1�{-1��δB���'b��O�8�QP�m;Q_�(S-6�]>���� �M�$t�"��M��4\�ZgN?�>�.mx�����0��y��.>�����
�F5�B�x_=�d,8xV��)��%����5���|���jː�Ă��d^"��N0�ڽk�̡�,�/�:��gL����ɔ�C�k�a����J��u�R�^�t/Ͼh""�<�ĉ���t�>�o�**a'��'Q*�u�3Z�g�52�J��R[McZ����k�_@B�L��['����� R�J+�f;H��,j���_B����\;DFEӂ�Kճ��������9�:��8���vlڻ�u�l�gv���>�`���U�o-��w����[v����#4�f�}:�|2�b�$�(0RԄ�F�@[ܬj��?W�X6���h�-�y��Sd*>8�m�}f�d�vw���Jo^�|lj�Ue�)��r	N��ᐌ-q����u1��
�KQ`�U�$�)����z�|��!�%B�Zd���M&����B*,���5W_���\x�{����vk{�-����O��Zf4;�r%J�-g�ńb�T��I�q9�q�ҩHG.8�}9��`?�|,_~�f�L?p�~�-�z�mp9U���fe����ySf�Ա�x�$��Ơ�{�{M��k����O|�B��H�I�ј��~���ڽG� H�}�9l�k᭮��-m�tW�:V7��h�#�@S�.��;6���
� C31�J���0�#���JVX�oݺ3�ӊȦ�Z5�A�J�-�<!"G2
�Si��=J���s6�`��k)�7EZ��Hd�,�W]C��zy���i�'�lTΜ��A�WL�}h>^-1�L�Cр��V�ص[����$y�>Se�$}Q�Õ����k7�U��Fnd��AH����9j�T�T{�۔r]}���R<HtQ{S��7�wׂB0T��1��Qy��Tc���IV�u h�$����o5�Z�z=l���J��]2�B/��>Xmv�b0��������uk�e|�������x��٘;sV��I�k��[6�X���$I��qlMT;����L��r����TUKR�w�XMʉ�g'+��!	df+'7*J����H�����*@Ʉқ����bQ�f�<Hg8��%#���XPgem�w^/gƹ�8����?�>k��<�f�Y��I(嫵�N9���څ�7���f$���AN��FQ-�>g�~r��������V�S��&FLfd¦��v�ɤȇi�jݮx,-c�J"�y�6T5�!V�a(�7�y�}��~����?s�G����G�r��=÷E��z�����ۍr<�|,����@�Zn0ᾪ`^	,\�����Q�m���.�C�}:up
��d���>�J	T+s�v�J�+�x䆋3�*����-����y���l^�k���d�_���p������Qr���A�O��Q@.��I�����ݳ�Oz�?��ᚚ���Z��;�n���{��Ҽh"宮���40L�F�
<`X�����:	3�s������Ѓ�MEE�2I2w�l��1�~���ካ���գ����А��0�H.�y��)b�~�tB����#���	�'�|��|�;�?>^y�/�ܷO�ٻ�m�Ã�q��W����a����&F�*:̀�iF�ω�}U�2L% 3��ȼ8�D*.	����9:�k㡰w�n��Y�k�&�}�������a��!���D}m��X�{}%xc4
tMȞV��b�4O	S�Jdy�~�mWA���dO&����1��v=�edU��\M�಻1TP?ר:J�G�R�v&f�kj;D����ʤ������s>�{�3D�\�_V�'	NU�����$Ol�+�1�d2�V@em�^��%��!����9nذa�w��aEG�[y~i	��3�`�)o^k94cƠm���H;��p(C���	-���9�l���n&L~��8�83�bwI��JD�8�^aB�$Pc���{.������Ͻ����ĶͩdEG�P­T����2ɉ��!C2�d[�m?~��}�k��0�����*�Y_�q��W�\���ٵk�$�\C|_&�D/�٭ֆ��E��B/���g�p�B�5_�j���؎#׉���������+m�������t���95���k�9J���}tm�CCr��c�Jlp`��������>�k�஫��{{Əm���>����uj�����O>������5����QC�m(���Dhؠ��Q9H /�fX0�
�[��t�@a�z�d���Z �Ե1 �.{�2�Q6(�!Q�Rc8|'pS��zbe����Sa'��i�b���T�c�Rz*A�뒔�ɘr����;+T~]���y�
�R�z�gIe2J!�-կ^��s~��SO��O���c���u��ҫ�oA�25�/���EXB0:�hWI���*y!!Q���X( 90��g���E8D��,��,�(��b�AD(^}��Rq�K�,�,���n6�.R��+s�<��H��A4��"5��D�[�|�	�c����;�`ˮ꾯3���ƞ'�$$u7 `cىQ"%"�r���+!�q%�*���/���*�b�P��Se;W�8�&!FBb���jz��ݯ_���霳������I�R�I�Z������g�����ks{[�:h�Ko~A��?��G�����"0�I������$o������W�_�XxI]�9����t�z��t��|̢J[��?ܶh��z��2 /�k��+��ҟ���îr	(�d��r�`�f��v\�H��1����?�r��$.��q3>?�=.����O*
F���Յ�֒'�9�}(Tm��X{O�	��B~�����|"iP�]�Q8�-�J��j���ڀ�,Wã�2&2�Vib�Dt��X�'c��yx����q��X�o$W#A�����=��������%{�P� �c�����TP�G8���(�R��[r��1-�D���C2m+�G�q��%M#F��u�(/�W�pn%sY����r�`���1���liMy0�|�g���v�M^~�E��׾�ϓV�ȅy�cu�:k�y�+鳞��TM*T�\Tq1�u�l��Z�#�J�a.Œ�x�q�F��>4%U�ZE�3�6J�d��h�������b�8q��_x�[�!o~��Qk���&���}��K�N�:��}�G�����g���a!~����;��ۏ�_���e�8��}S�ܸ|A*�ӯmJ�A'R���K��S͟3��)��AI7ˌ��y!���@����NJ$b9�Z;o�ڐ�S�jd�	k�%���X�L��Pm�g1Ă��A��@���
"���d���jwv7Ny$U�S7a��5)��I�B����:s���������3g��҉8�~瓟�����|cy������g��v����:�Z��)NT"���{�Lh]���y���/�ßW-�M4�[��Mu�    IDATvSS�tB��|�y��~Rst�����bZe�C��(�q��l놔*$��H}�܆Zˉ�����X`��V��h��ܜ,�=,��܃���%��HJ�.N
�!�T�/LI'sr�[ߔ)J�#�����mR�4q�J@+ZS���yC�� Z���N�ǲ6�\zjjZ�UBdޒÇȵ/Iڱj��sB�E&���������k���Ո�1�,�HB�vX��75�5�����J�Օ�K׭:!0�q�����U��*=��j 3�8V88�K����l��q���`̹��(?n��a^[��8�xgLh����q ��bo���7�"���Z��ZǱ:�p-�Fb�Ơ��o�A��b�o�wS�����m��p�-{�{ޖ���ʕ"aKj��	
v*�o���\W��!M��a�������`�ێ�g��pj�H@�g�o< 33�*q��щ��:tô�$����Cmøbй����H����v�5漵�@ I���?��`nG�4n���v_K�ol��S��q$8w�9𔧭�S�=�N�8���]ɞ8��?�����<q+)�k�O�������y���������~��O]��7s
��v#7_�(����[}iJ�5{���P2ͩa̭m'��5�,�䴕�NS�i3����j(�j��I�d"s�a�Cv��PV@�!�WE��q)�kн��8W��9���b�9�!�2�s�*���|S��
K�!�B�R!!P5d4q��&7�����������{�{���N�?z��#������o>y�ݾ��ms�l9~Jn��k�fH�u4B�Wy���:N?�H���-�6���w�;����3]��3=c
U�� �7ƌ�����C,�l����q����
�0
��a�o&�bDD Kj��>Q���|��e�#H��ˈ��o�r�༴�Z�h[^���̷��j:��PIR�^�]�]���L�{D�/\y޴ǛZ|Mι��`D!8G�]#��H�9��@����4�!#�����{����
p�x#�|�Iٟj���5"5U=�j�'q��<m(��cnl�\�+�W�VEG�A�!a.������8��$X� ���R���"S&q��}���	��vD�DpZ�Lx���~i�=���l@zi��H3�-��qb*g�o�kfЍ�����s}lt��C_Q��QW�h-�!Iё��*:���U��9�J���$�X��r���i�rcI;�!�j�,�#�J��N�	d��tj��R:�JE[B-�J�����^�#��ǵ��08[8L\c�1��t&�;�x��K:�ٿ��d���ҧqAO@U0��<�r^Αc�s�_�롁���Yo����W�ȝἹ���i6��A�]�{�ʱ�(����&��k]��ޣ'��篽����/>z��s?X��5�{���/���=��6d�v����CY������T��4�!��L��Z_��dRQ�F�k��8m�����E�}ǋ�,xxf�Ԭc�a��hEtZl����U� ��+�*��U�<�-�`��	�'2��-�����;=%3�=��1��D��ڶRw�e�t�W{֚{A���Te��������ݻ��_�s�V'������?���?��/��Ǟ|ߨ*ι�3;.Y�wP^���+�Л��^�%���AG-�U��2�ZY���)Y_� �7�ц�3uX��5�0u7�Z��Ʊ��O��?FOJ��%.Rq�|'��&6����5�Ĝ�۽�:��䯛J�gZ�C���_囏<$S��D�a�i�kr9�ߣ������O�S�g9���p�� ���d,m<����r��yE"(���bd�s� ��ݢ����B;ۛѼ�����Ҡ��-�[�q\#L��8h �����S]j�ᓰ���Vu���.t=�ֶb�c!�)c��Q���t��P�B�eF#t撊x|�A�AtG^w�u��0F�FN�{�udC>�}!`�/�p1z8�Q������eeuS��6��wў���� �e<Eh4�P�X�\dm冼��U��'����+Խ���,lRs
��#>?�!��]����F����A�H�~��ʞ����B�c^�}`|xdƃ��O����~s�M�q��!�w�<~6Q/F��ii�E�	u�#D���X8����sC�������7�?��\�n�U=1�ёP$-�Z4N��<!g�8'�]��O9�)$��Z��1���o;}������}�}A��������7^�ট{c��E���/]�RS��2�'� �T����jCrS��&����6&q�MәZZ�ߦBe�{P��o� ��
���54�Ù���17�́�<�##s�s�J1��X�x�x��D����נ�
JH��L[U}zA{iʫs�O�v�ؗ��_��O��������������~���3O<~�3�ş�p��{��祥bnT�2��#����-�	�aI 5�a��b4N�h� �y�y7C6�[Z�Ң����5Gh%��"�
�I�J�
U�
��)H�Vk��ۜ����}����Y����Y(p�ZI�9`rՊ
�G�ޞ����E�	q�q��l�-��ɱ���������\��٬{���SX�5�%l�ݹ�D
,���\���9%��1��M���4��6Y`B�3�j�7�t�X��LS����l�u�`�Y\�ƕlJ��nKn�J��Y�̌�h� ܍���;��w~>x���d\�CF73��pR$#��h}�ؼ'-V�Pߧ��/_�h�1D�T�d��Y\�wG���/M�h����~V�;�@���`i2�g�{������W�x������p�F�	��!����>}Z��gΟ�Z���EY�ؔ��uI2�x%�1D�j�U
���f����q_���7��W���Xo{˛Tǜ��v���{��x�HU"8I4��Y�3V�����cc�wR1��Y�.?�\VJ@��}Y�~U�x盵�� �u�T&�M�J��΋fB8�
m�T��VW,*�	��lij�
�-��81��Y��_�M���}��E�ν�"qN`�!�F�="Tс�fL�6eX�EV�s�H4�㷟���_y�֓�~���կ��ɓ'���_���Q����O<�+�r����aS��G��|]
���4d!�BN�z��4cC���L��_�TV��%n��'��5ȩ��$t	��ӼKc������6�l�K�ǈ�V�Id��u�2��Pe�c�ŉȟ�&1���-�:Rl��޻g�+"=~#{d8ڒ�M�DѳW��S�'�������Աc��zݑk�����YVu[�t{�.�G[S矹x��Ͻ�ŗ_���͵;GUs�5yw\g�H[ȟ_[&%�t\]lՈ@�Ay��0Bd�a�+8RKo����LO�#%x����V��W��U�F��֦D��e����C�W���') �7�~8g����
��Em��f2��䝮��*r/�n.����\O����r�W���^�v�����w향
qsr�_��7dvq�6�Q�ܨ��?��E�981�!�e~����ϢC$�"�C�a����4,�Dd�]K�.]�sCKcuˑ[�����v�puhX���^	���$��q#b��q;o�P9�����yH�J�c��D�]�Z_��A�����]�v�Z~U(������lZ�L�f�"'��ͩ�u�%P~ī� 8�8�1O��	5zx��1��C9h6b�<�|�̙3:�WVV5Oޚ���`(+��K����?7muC�h|� V�8eο�Mwʳ�|K{ҟ{�����mhy�pZp��/�z���" �t k��lm3XY���̫9\�}�gN^3\�L�q腁\����t;S2.q̌/D���ı�ED����Ր2������O��Vy�f8:�9�cͼ���w-;F�f�^�v�����t������·<+8r�S��8�w�c��p���I ���)�Y�i�ӷb�/�>q�?�_?�{t}������3��Ǐ�y��?p}��ە����g�Ѐ�$b557���x:�y�9=�Ǻ�J`���Zc)���Z(*�H��+#g]���A<"."ܘ�-F�nQ�=0q��4Kn�]����1Ѣ�l��t�S�<b<cE�#�x���М�'�ۓ�ׯʩ[O����RSӚ��e�✌˾L����n���t�ҁ��K�3S/�I1ʓ,����������������pt����d8b�r�L��bt}M��E��15��+�h�Z|Q�HΘ �gI�S��V�2�^/cA���9��E4 h{�^9�>�h�݋}�W���2ob�X��ތ��էip筶��  ��#u��A 7&��0++7�Mw�^^�V����D�իҌ��ӏ9T�?����M����k<tp��1d
7�4�(d}sKk�EאO�Q¦��d@.螶t�@����c9v���/���������]!LD��������U�u{*��):��$Pm4S+�O�(�Ű���fR{'��J{�#7��uʓSe�kYT]��܂�o�����A���m���S��-�����?��)�jP�Pm��i��#t�C�5�c�Ղ厨���Pr^p�L[���ǈ1g8�hh��m|�h�y� �8���C�-�r*��r��9Y]_���%*]#[��P�A��9�L��gv�'뫫Z�wa^���7K5�#?$���A[��@��g�s@U ]� 5�V9丙��aߓ� i��&F���4b��2�14��5���y��m'����3*���G����gypK�X�����@�����9{V���+Wԑa��<�S���Yu&�����WQ�L�sjN�eRK�C�q��)��5I�M�׀�8Qt�Keq/�]jS!I8<(x���ZՓ7�	��MZ7�~��4:t��H��:yJ����S��8�K���'��{1���9���K�>�{����~�箯�Ni�]��Q��y���f)�N��,<�6�� R�L/ݑ��C?d�{��[��n��,B�@��Qݍ�ߣ1��N� �G����&Qy��q_J�����p�BnPv4d�����,jTy�5�HBA]s?U={��v+���y:L|3N���gE��v�\�9���ȶVp
@H9<���h�E�ݜ�R=P�A�'���8�-i�ɡ#��mߍ�k� CX�C�����a�zB�yƔ�ޫWu�����#̆8dj��Ñ��-��^SJ�M?����R��d喌�7U��H$��a ������4}��Ȱb�P�A�bd�ʔ/-Ggs�Q#!j�>��7dn��v�Z��T�.��(�%�@6�����G�Р���K/i�!�����H�muZJ��e�VJmR�`���k��Y��G�H�����LJ�D�qO�L#{_�4���F#f�NPQ�{*u�M��EL=����PYNW���JP0/�s!���"7�w�
�>�B c#�̙۵�'��} ����p�'@N�*K͡S5�D*�� ���R���w˗���,�\I�-�䶭���g����>�����V;�u��w����ȍ׵��MK9:��ˋ/�9`s�r��,�q����J�UP&
"D��<�on���ix�w�"@�Ք�u�����f[[���0?���u>�����8��C1��g]�HB�)gG
GG�{%\f���&W��,y��@�66� �
Ņ�=�N_�7��z9���\y�\x����ط�O��n�o��c�e��ե�� 1�*[��P-I�֊���b��W<��^\P5�Ǿ��v�\�̵,eρҙ��Wo\�����K��������F �����Ͼ�O|��=z�'WV����nM�y�/���V���Rٿ�^��+����j5�(�9�љ�,���z�H���K����ݧ�s>,:��¯n�kT!���D�]������@�A$!D�!���b��<%�P.ԩ�\���Y����[�(G%h-7O�"0�m>�H�O��Z�-��&+,�Gei[����;�~5���8~*�����Ϯ���Q���,�Ǔ���a�
F�y�r�1����Ӆ�2�MP����x\��^V��<Ӻ�.m_�Z�ҥaQ_�E��!��a�a�2r֌9b����l)�A4o�IM[��	����aX�9��7t!5�j�Ɔ���!'[S1@
 �8����� y�L����E��֛c+	eQMr�nA��E��������o !O�� �07�7D8~�f��'b�w޹^���ɱ��lD��A��d�e��lmm���!A!.�8v$�ahL�]k�+��8T�_��Ź��'�����p�i��S��޽�o����VǍ��}O�v)ּ��G��O?#�}m�A��]���!�2�88������u���Tjǭzƞ�L��&U n���F�[�~4U1��	�RU�Sj�Ky8F�D��;���;N����k�^`���<�~�y��P����I���cj��2���l�=ƙ���
�L�d$�s���y�<��y�"��Z�������7�e}uM�ǅ=��1Ϛ�ĀO���1P�c}[�\���E����f�����S��������b��"t���^���������ñ����{��!d�F8�°ӳB�݌4�Es"t^�8��>�AW�&.�U�o� ��x{b4&���\��پS��@5V>F�& �
88@:j�5��]_1����9�������}%��<��6N��\�u,�w��̐�CX�	kV� ��C"�^�ߊ�݉���e�܂��D�":&��Q'*8P�	c�� ;HF��8�vo�} �=d�R��P㬍{����p�L�pvn^�_x��bX����V�xԮ��S9s��@�~�x����W��|�k!����K2.%W�A=�@�qW9�$��1�X�5�l[���Ѥ$���߉�qF0�8�@��J#;��aZIB,���VU䆸�/��p�:yײ�<�ń�(�g!����"��,nSĐG(CN
�k�`�XD�P" ���g����n�����̧4��}$B�`���Zk�1����8���c�8ƾp�X�c.�����Q��A:Z�bԩ���t�.(�Q��3Cꆹ637��2ה�Hn�1��AS��ć�kG�Q!���ط2m8Ų���>��������j4��Hk1��8M�qC9mtfb�@ ������4Vb(�mՑ�<@�z��<�H������d����Ls�+��ǌ�Ӏ��~_� �G�; �����*"Q�Km܃��⾽2?3��}�t�,d~Ϣ:|8�ڄg0P����0�A�pPT\h<VGzϾE���< O���a�������?m�?��5i��/�������>��3?5�߰��1?�;UY���τ*K�}Q�7>q�rM=v��W�M�F)B-J�rU�(+�7��Υ��I��l�^�N=� ��J�Y��׮����4��4>�)��L��z��#>�AvE%R�������ȥeH2��G.=��o�?4�a!TE1�m�T�V}����U���f^kÓ�����vg'�S�_���$MӤ��P,cW�G�����x���H���;4��!�$�f��S���t�,Ip���v��4�b���o�������{����
r�E�јO��px�Ɛyf��6�Bf�d��`&��$M}���O��g~a��СC�[O>����}R�Y��[�G��u
�:I�������sϥ���4M�fYA*�W�l�)i��-aH�����I曄�����1�3i�i�]4���窦�k��n��L���d��d�c�X5�:Emhĝ��<��|�S$�JX罷�u��z=_�u�el��`���P�����	��=_���s~�]T ��Ѷ��3���X��de�Q�	�z]#�q\��={u?׮]k<�R�G]{���m]1D�p0ޱ[�����;F��+B��'��r�7&o:�V�ҥ�|(S%B�M[R"s��Q�&��ߡ-^w r|��A�4Kڨ�L+���s$}Zl�bwׅ�q����xu�]�u����US��S�  EIDAT��B��$U� ��i��(��9��x��!�j���Xؼ�	jX�&$V��t&��
ٞ��iz�8��0D-�H�%H��T�2pb5�*�@���e1��c��q*"jg0����{fN�ܤQ5�\��O��=�?|�C����ɦ�Y�����/?��oXn�����x�qU���%�ڒ�N�n���,Eu�ŕ��U;W�q����h��q,X̰J��Jj1��4.)��.ɜ��kI��L�&M \�Z�����w94�&�iU��NKH�D�t��ƻL-�-&޻$�I�z�1�b��5�`�\�ڎ��RI�
�5M�j�z��4�i��M��yZՍG]��F��Ƨ]�M+I��V�iS��I�4��`I�|դ���?�7�2�����rh���3n\A�&M�����.%�d� b򤌊���>�����0�D1_5M��#p]���[�s��C²��!��9�{������,���-pS=��o��x:6,K��4���I��]����]L�z����a�q6�
sG�4IH�����+�aѝ����y�����v�ݝ��<��p;/ZN��G����\�""�p�����)ǰb<FWeE���ոl
d=\�ҷ�|���z�W����&N���%k�p��$m�W����+����[U�j��I�gI�����ey^�-�� &veV�.�&�\�a��I���#�!��7z�Z��s-�t6˕;�a�S\�Oo�C�vU�j�Y�U�I��S��o�VZy��,m6��y*f}�E�m�*��|��o%Yޞ��Y!o;��h4?7;�R�UQU��j��ʧY��*�R�G^�-�\ݤiμM�<V��zM[ĒN���I�4�o�̆��'i���֨v>'�H�2�{�%�{xEZ���s&^^�ֆ�%����A��.���G��ZC���?gY���Q��CXWUYM�˝K���Q�"`��3"��)���6�c��
U�#o��	r|�Coz �EҊ|�4��׆F���L���岹�"R�t�:t��b�)%RK������s!�j#!�HHS@�D����@i��Z���)prBZG���ZD�O��,͟.Zş������{�?y��Ø�����������e~�����X����!������R�FҼ�V)e�>�/"�/H�����Rמ���J���2=v2��O���P�o�F�����"�oK~s��w�֜��oԼ���ܶ��h�����lldk+�daO9���Z��s���R>,���a�yʉ��z�瓥n790<ꗺ/Mփá��r{&�$��tZl��jn���әi����ܻ��n���i�}������qϾ�}i����h����B�k���W�>�X��"���7(��+��ߛ�H�J�w �Y�ߑ��d,2ri��I�hCu>rn�sߤ�V��n�ʠ;���lQ�V��ޥ���4񭼓du2�6���|c�5��;D��|��"O�$kr_ʨ�����e�W�ϋV!-I��p�$I��y6�&f�N�N�~E8\�%i�\�e�uP�-4j��Ns���d]d��M�J�,\���@ yu�,�u��aʽ�2��ʖ4�*]�v5����>˲�j�y]�m5�i�nH���HӜ�:�*��"��wS�&��,K����>:HJ���4�Uy��U�)��$^��EC�h�&I��ܦ��wV7�;�zy�Ӭ��zB�N���K��7��8	Q��s8n��d0� ��Ay�x���L��:��wp8��omod�N�y�`��w�s.�m%��v�$�CP��!}�4M㊢(�v[[[I����4�z��<oF��{�]^pپ"X��Q�^2�ۛ��6b{د�{�O�����o�q�/>�����՝�����G����\    IEND�B`�PK   ��6X\�
�@ 6 /   images/56cf4bf5-9c71-4f2a-9d5e-98f1de214099.pngL{eT�]�61t ���HK7!]�0tJ	CIH� �twH" !�H7�����~�]�Ǭ5?�Ϲ���u��H�7
xؔ�HHHx`E9M$$
$$�_����KG��5d�ʇ�o#!�"�夵�M���R�{�η=l�̓�����Y�?�R�� b#y4��8�x�y��L�|��?$4�F��Fɣ��D#[�&e��d7�vpoHwn��1��<R�u6�}�~U}~c����X%�,��,�7������,�ak��n���X]u�[�l�Ծ�e�}����1չ}�^o���Ɓ��10\.Hw��v�bZA�ee��/��Q2��A@x)�$曼�����ꔧ.|�v�̦+�i��Z��cf��6d6<�|4T}�z�e�%��⡼m��Ԥ�)U_�p��&�!!T�?��ʆG�e��G��n{\�EEE��_�/t�d��S��2�ݭ0�2���g{���W�8���<��;t9��nc$����W!ua��D9z���%%�vNN:�!���}���=��x���ݫߏ�b��c�(��Țh>�|�kB���.�Ѥ�)^@�D�*:���7�2Oo��
�W\�������N8��8Fj��k�ު����֢>-ה����=O,+?8?^�Nz��k#.J��hAm6�ʼ�Y����BРg�K�§M���������7��yZjDN�%"����y-bE辪UF;�/.p^h�I5�i�#z���o7��0�9����hb�ZB6�?���Y�)X-G�&�^k(�"=o�v���Fը����ŉ|�y�Q1���t6F�;���u,����Xу���k����o;���m'�S���o�qm�E�EHE��uzGt��B�.˅⬆���8�nS�ˡ�k��5>'�u�ʖ+.������О�����J8t�!�����B�ds�lU����Y%�2;u���֤�Ñ����*U2���n>w y9�B)�-���T̛��d #�"��>��aHRr�V����X53������"���w��S�N�<-A@5-���8�6�2�9��]�'��%E�*㧑\����grc�i�L�ûLljDB7C��[1?�s�T��q0���_}�, 1#6W��Z"���J9���?kYZ��ZS�x����?��"�ߘ[��۝���'K
�B��F`�Q�=�}���%ҊRIZ�(T�6P�$��QѾSr���ȋ�7ʓ� P>C��dg��*М��2de]���QQ�u���-�7���m�.x5�b.Öc�q?F�g]��EJ����W�@LZ4��2m�KÎBKAu+~�o��F7����N��9}�_����wԳ�.Ol���u��3��Ч���;�#�:��`)�����|�-}�V]�[#&֘���U�NX��2<�R�UJ,��+�p)����-͆�j���d�~����^��m�5�8���l�s�JX|E�ɬ�����J<V�{�)q�����j͖7 D��4��w��B��{5+��|�4��h�E�t��igR���|Y��pw���
�e����B� ��oe�|�[A�c3\J 24$��MBzoL����wn0mx7Q䆳9�6����U�Z/��Fy�E�[ڣ� �n�_Ǵ۵��+�q�yo^��x]�x#�0�м��K�,��Y9k��Ȋ�K���������@��c��6@ļ9�~?�ӏ���?no�S�.��D���1(�����ҟ��t-��Z�xp�!xln(][�3��1������n��p]�	��ݤ�ut��C�>�F���҃��2At�w�'��|���F�N�:\���ѥ7����|�B�YUEN�������s�G��7w����k����pN"ĝvZ����n^B.�C)N�>Ke-��%z�Xo�e�D���1���5k���n��U'�S�ɑ5|\_�m��uD�¨�cI��T�[� 9N�u<��sW�e�K+�E�d��ˇ	�ͧrԐMI7�4�%�[�n�X�5uY��ߗ�Sb����J����P���\ܲ����T���j��?,G2gm�/���߅���!M�p��ji%h"��m�&��O��2tK�N�'�,)�Ka�bz�6d�˼v�J��ϳÙ���0Y�+��m��������N}�qy��q��ɋc�E���;j��c_�E??�m���=$�'�@�ȏh��I��k�@x�E�f�uX� u�:~HvM
Y_��GC�v2"{��k��"K.�b��Ԡv���.�{��w�X>Uͬ��᠅f�tk�`����zMT�#J��k�I�yӡ�m�N��qQ�_�1=V�g��Z,����?���k*����l�c������ׯݧ���$ͦ���|���~��4�Wh}�w��i-b�Q��{�w�b��k��X���˗��~v�*3]�hKsϸ$	c��r�ɂ�.�#$����g9[�Oo>֕Ko�J|�L�4nv�3���鋹�l�j��he܃=q�ƧļL<ov��P�{V�u0�j�[��F������T�
QTS�RرQK������e�ވ�-�?v����"�!��ὸq:������|����䥎����Vo�$��YQ��k�:;�g(]���g@�����o�T-Śu�lKj����l��s�8���c���X���٩�M[f�ߗ��hi��،�Q�_o��^�Fs�]��>g���Jx����Nߟ�y����B�&�0���`�kB'i�4�o� �	8���!-�k$��Mr�Z ��p���i��xc����ZB�p3�n�$�|N��$��M���w���w֜d�RD<�i��vV|���]GR�c&A�Fq��nR^?�%�K��<OK�����9�d�+Gt�ɱFo
��_�w�j�J�t���9�I�d���I@[fV��_���~�3�3xl����}�X�P5hܺ;%���(���?G�G�GA&�w�����U ��������%/��1(F�Ág߳[�`�m"��ӒO�R󼜏�+P+�$������t<���1�O�1��'����L���>h�=�[�uY�̫�F�0ᐟE��G:�Z=��"Z�&����S$����RƉ=~�(�����(�~Gok�Q���� 	��ـT�;����������8"ŨM�+\�|�UE���Yn������d>�//�?��z�����b��q�=�"���;.�/l��^g���D���gJ-|{��n�<*_�C�hq@2>\�KW�6�������~�aSѷI��H#K���i�*��1���u\Y�ˋ��ϖa�0ld��L��o�y>"j:��|�ܠu�
�c}��!��'��F�(�M�����?[_�R�y�� �N)��'��8�FB��w��M��r��V����*�(}!�8�2ڬ4!K�X������W��^�A�ԥ��F��X�y�Ƽw�)�m(���r�.�周�>�&���g��p�����0SB���Kl i��k���v����iiS8N������ƱB6����[�7��*h&.r�Fr:5�$����N	>!����6W�um���^i�װ�r�����ZH^�f��m��|l�O5�ښ��/Bg����-��|
�xR�G��׊av��SWY `�^�R�%�ի�	���Y���ZE������s�t�����~�H����)o��<@�yQ�$Ĕ�������"wѦ���C���q��s������	�M�~�!�������~�vm�[�0?��[Q'O;��_
B�տ��9?+����%��bϯ�>�k���pXɾZ�"��*��X��~�4G�D6b�X�Ș#۲�|SRr�w�k#w� ���/̜`���$oBX��)=h�#�)��X-�B��:(��A���-Yٔ��qsU�a�[I[@�V���t�X/�.����{�d.��Z���x�!����%I��9�7ʋ��$��b1d��v�;$���핆��T������������X���ZRj��a��s(��C?F��|Ξ�_���=��c�������E�XsX�4���f�<�F��V�e��[��J�#�� ���:���B�&�����?�`?"�7d�V�pV����^���_ZD��֯;��TE�ޛ���v7ul����`�������I���ǂzS��ѿ�Pp�_QQV�e܈�g�D.����i�9�^>��YCH��z"���L>UO����Ǫ_�:=��Zڈ_�W��!& ��i0P�v��;FKJW�I\0 U�hfr��9T�G����P0�H0D\���X� �5��)78�����Q\={G?�����e*o�2~�ζ�c���o]���Fx/�bgW�X��)��_�`��D����3�ۃ��/���-��Ί���p��h#:d��Jk8����P�L*��Ԙb�~B�h�7)y8:��u={z��<s����7ʼr�A�+�)���?b˯��w}~�P
���e.���6�;�;`���	�����;i�K���G�$%����M����B��o{�{��z��$��nRd0'fQkl��b���FU���u�v�W�y"CgL�:dx^�Oπp
�A_����[�A�i��W�&�j��i��ň������K��__�L��*��� d'!��?�����~���-O;���a_���I�3���9}�H4�6�m��<��A����.)D�5�������F_��G�,6��9�R�Qr��e%>��%l�G��*4�'�6L*)������_���§r���;�I,�j��m����ڍ_���� 6���:�H��"�i��F�W�C�l]��ʹ���L>��Ī@u­P��#��K�9���t�遐�b.�5�쥊�{�c!կ��&˽��$��l�)�t��G�B�lBK����橃��D4l�c;�����e��p����?����&7梫&��U��AQE��ۂ-�?d�C��*�)�yd�	�)G�Ak~��2X�>ʎ�ю!�P,= �pr��!�8ҽG8�}ǁ"���2�T[[_0�C=���o��H=�9,�xj�<�hfg��E����*,>z��I���;N΂͌{ooX��4RF)�$�e+ L�Q�Gk{�W9�7�9#P��I��+g?��f�$�z��X7����G����gҵE��_�h`�N�����q��k����n�?���I`V�/���Y�G�c�(��{����f�*M����a��$>���M��D���*�+����nZ,��/Ӻ���2�\�?��"��	~��������Y�F+��@��C��^��|��Џ�w�@�V�dnC���n��3�S�m��ܕت/�q�y�0ٕ����"w��#���OrŜ���铓�?�z��~��L��ü8	��	);p��c<D�� z⧰0�Bz��D\4:c2��,�K(D�FL��I���($rL�<l����O�0TI�<�����3��K$����	[TVդ��(���QnP���p���l.v���N~O�|0j0��F�ug�������c�����7���'o���#�G��[F~
�]-��SR��`��ت��7c��ʬ�~3"J�\6)ܲ�������(��f��#���}r��9@[��*Q��L (��N�qVċ�5Ɩ�S�Sx�"VM��(�}i*�X,D��m����3u�HI��!�"G���t1����,���m��7iqju��lN���0�@p�ϝ�3�Mc�������Ϸ(�T*
�wܖ(*��:�u��7Ю����6��X���e�D%n�������ۏ�?���p8��(�Ni1w�;��g�A�Rs��g�&�_��r��&m$�O`#�4~c;�j�U��
�BA����bvwh�T�|����w9K��*�9�Ns��@G�S��Y),=pC@���ov���H�.gt8�lQ":��3�YB�~:\��@�z@ڰ��$6P���m��D.m���Hs����:ǳ+���'�I��?��~|}�쳑O4�����`9���Ÿ�o�ks���6=.$[�Ą��#���N�|Xn�``�g{���!A��[��ULY��1��1Ê��
��-���x�te��9�&O+��{�U�x�.Z�o�*,y�o>�Ni|�޸�5�{R�O����z<W�_�ɻ�XC�oo���}ގeIs���Wb2ueb��vN�{�*��K�c$ 2�v D@�nm�8��MD%9�da�&�[5�դ|k�Z�ť�r����Oz�Y8f]����4���Ҋe��y���3�?��\us����4��֬L�+o�\��~�^<�sR�p��^yTs�5�G�#Vъd��ג��Un��^��S�Ѭ���_2V".pX��l���'�.Lx�mgK`1*�����ID���3��}7������%S�t������񻉢{u_��7��{<���π�ʗ&y����'u�^�4��㸏J��rw��v��㣌a�b�����N�F�[E�9JC\ ߇�����Z�������B��)ɐ�+�$��&oȴ�i�%T��4!g'Z����H5�;���X�dt����3��}�L����\��T�Y�x�S�쒘I�{�g����:���Ϛs��o\�͵'�wv�T�/	XrI�<Rl��W�^������H�q���� `�hDψ=TN4�Z@��P�f�g걮��N�h�l��ڵ���<�r�Jm��)�L�N�Q�<�l�J"�-C�>�\�z4<+V�~��M*��+�gBc���b��٬����vSg����w��а�Zu�����k8՗��*�O�Ă�..�NE��)�H�d@<Xb݁�N��x�Nv�ʺH��<=�03.I�)�
�dO4֌�Ѱ�� n%ê"O~�Į3�Z]���+�x����w�вF�u���[л���{}�l��,���r˃�,�[�'!���E���ƹ�c���ǥ<o*���s�mc���^'�X��(�W��n$��5{`��Y�%��x�\(J5����D,]�L��y��]%$�@ϵʶ�A�n���7w2�z���v��VY4�^YNc��U	�����S�5Z�aJ��>5���LjY�ӗ�k�{���E���̟�b/��՛2Æ���xoB��*����B؃#>����C�A�2<�����(��>�Q�#����=,��ҧ-瞤����"�1�G��"2$� �U��_�������[��Tg� F�8�l��j4������vb�O7]qпy¾�s�O�C����s����qAW������S�t���J ����uB���&��İ������`�RSv"�2?�zfd	r�	tq�-Dŗ�2�8��L^1$�[�=�#�&��
���)�r���,�e�xyD�o�~Q˖X�ٜ�3;-`�_{E�F�n~��D�و���jo��%ߥl��dEe3=&�*7�]����9�n���:�(i���*R�¡Q�I�'������d�j�Fۧ�����&.��7i$nx��ԧ)�L���w/@`W�͐�O����U׽�)r�T�A 
�)�a<x�pl^��AJZt�i���N���bw�"��w�=N�\���|���������g�ټY*���7ti��!�I�t�+.�O�r�H&���5*V
�*}��n޺Nu}�f��L
������F$'w2�D�a�� آ��z�j�{\�\K}ٶ���t(�6 �2Ȁ�|!;�Wm�HCK&��)���0�	��GuHs	��7{l�y�����{m7�[H���x��=���t�ٴ>��綳sC*��7��!�Og!s�uu:���b5���7R�&�:U@)+v;�S����>�_�vw��f��VKK��O�,�S�Q�A�5_�j	S
˶��A�;�{
��o����;�z@`�I��C �#}��I�z�e�}�PBA�ˏk�fϞ����9�++�/N̏tn��me����Y ҝs��ê���%&��p�d��-�x4��"F"�� ���{�Z�d���2�9�j�~�O�|
PO�>NK�h9��G_�7��gI�`��='A��dT�O��u[�Q���q���,6����O�nK�2]0��ء��n�R?���.�B��}�����̈�|�E�7�MS���Y�&~��t8�8O9�����s�����p��[s��w=�ޙZ�R;Bl��߿�7����P�l��#�g���
�`���n��L��w<ȉ����#8(r��>�4��k-��s ���c}y�J�e��N?}F֍#�H�w�:ܾ9P��m����ޑ�&4�Ƥ�ὃ����t����^����y
�ʇ2c������⅋��/�.�����b-����s/��L�w�����e�␉����{�����=�Ú�!��]�X<G������
o2�P��D;���m���N��"�ޫ{R0��,^���%��`�:_�0�E�0�V�<{'0����'�X�����S��5���L�����%u*�֦�����c�kl��-�D�V_M�����:?o/}Ƽ}�d�G������m����^������]���j5�.�_%a���\R�˶��G7t b��ѝ�1c
1�� �_����\ʔ�c}���*p�N���9L�T���d�ǝR%L�l�]�p
3gv�ܰj�F�e�����&n����_e�>���|�Ȥ��r��Q���9xc�vXvy��d��ޝ�Q/�޺�L{5�PѶ�Ь�,$v�bmOm��P�F�l���~
�ąZ6�&�g:	����FԳ��83dE ��[�i���f�.̷����F���|vS �{z���'}e�XM��!�w�2���pd�$��0xך�E,X.���"z
�9���`I�EM�O��<0����pc���7W˩ qК�d�e��s(��в]��]����K�����H-��{4mY��-����z���7�w��s�cA�t��I6>��cr�uR���U�X>�e(<�G'�a�_ˉ�������nRю��r��5��p�f�t��]W�#/��(��)>.��#�28�S�o<��X~�E��>�+�;2� �������A/��Z�����EfS}N7�R~��}_;f��;ی����
�`�	n�L z��i��W���@��8!<�Ni�Ų{�׿vv�_�o�v�����/Ihc�JȠ�f°N@��s-	����y|�r��
D��Q��k?ОZN 	�Aā�x(�%>�k��ޱ$A`)u�_��V�?��{�;8$�1gp��FsV��p
 ����8���!��{zp����g#�&c�T�f�JIER�}$�ԝ��c����� �]�U#�FU�A; ւiN'�H�zMp!���/P,	G1�q������5I;M�иp +��0v��X2��@d��/��(JU���7�B�Kg�}$Mʶ�p _e* ���3m��BIiiF�q�Hx�Fegǭa��pS�ӿ��`�%Tv=g�����<���V?&�s,��wzE=�T��֐?a����&��ٸK&�@q���.)�B�k���7�،<�B�?��^A
�8�b����Mq����U����a��a\������UQ�MA9е#��!�:'Þ�l�ڸ�Y�Vo��jധu����-�vpS?5�K,8����Rp���1B��uՌV�$*g'�g���/�d�fl�u A�hɽ�W� "������de	�z�c�e�g�.�a�v�C�s��j�Ù�X��cFi��Z&���̄��Cw�#b���K��^��P۔e#�Ow��N�Q��T)J {�K��S�?
����#� ����ol-�xA(6il2(�2ύ�O��x>�u��S	� !�at�p�i�:clȬz���_�8��s��q?u�u7�m@r>����I�Ά�9.�]vA�S�Aޗ
��I-	�;�r���̭N��������/F	��*f����V�}R	v�ԫ^��݆�ϥ�W� " y4,ǰ���W�B��2�&���@�l���+O�`��xQ��n���pf�����KA��x|�S���k�Ӝ��_)��ߍ�,�":�����1л���ɥ�\����(���X�\1��t��n��I\?M�d�}У�q�w�YE� w�}&��A')٤���n�.,�5=�-�T�,��J��U����e��z)lZ�5!Bz*o���95��U���(%\dy8
�i�`4О�~,��[25a8&!���fjz����	ol�$���M8�}�5��,�6}1�!� �l����볤Qgf��A�4"�kVvu9�*����]�ل�55l>]�?���0T�8N�^H�^fC��@v��_4)���9Lz�Q���̗$=Pt�]l��1h�(F�a�S����K��&���`��U�J��	�%�m�����*qL��:�U�0f�F��QJ}�ѩ',�e?��a��zmQ��B�1"oo_ƄX�?8·�ָ�L����]I?ˀʗ�7�}���f)�o�d��Zv��w�+7RpdF�M��ӉWS�Ge�,���'�U��8����U�_�W�q8#y�9`玠̸�]�x�
ؙj��mmŻ��B��06�z���l��J_NH
'k�M<��˹�0M�y�$H1����ڒM�;:k0�0frPBN�N���l���I���$W�uq��G�4��"��I�YL_��-�������27�~��;�Mo^�����V�:2��i���H��;�jT8�zP���
��<�̺�����|�o��Ґ���̳�hY��Y8l��R�0i�pL`z�Q�
�����g����D}��t��x�x�]��d��`�9�5�̇�Zx��_x}c ���}/=�Te��b��3t6m�]�.��U~�3-�;f����PZ3��KP��)�6/����+	�$��co5FOY�P��'��U�)o��F��&��{�l~  $�������Bb�(J�b�Yu�cz3��F�m&5�x%0W���G��|>m\�v����Ths�����N�JUL��N(3��uMv�w�� �2)��o*]�
H�&�yR���eC7�Klb&Q�/���%�C�1��g�yA�e�����\V=˝�:��E���zOӱ�rx�RQ�M? �}~����OƝc�Nϱx�q����1��
��.������8^q���{�o�����|���(ok;,��n����܉#O!x��t<M��C�<0�>��A�6(J�*�1A���&t�	��}�<?�I]��+�uPzm�{Wh����\?'	�|��#�c�,|���7'�Sl(u�C��D��g��릑:�d ]����6�}7P���z�tm�N*�}[��<���9�[^�ty�����C"e����u�����0�}��Sk�6��[6���}M�G��U�g~<��#{E���~��h��m� �?c����c�������2=�ԄSz�{�܎��IC�]�dE������b.ubl���oKp���4����ت��q�R��l���{t���Dr'�1��9n�΂�J��V�ò#��؃����T�srڨ��h)9xF�F�a!�ޠ�F-����<P���F�d�U�;Pр`c����]տПq%7JJ=�7εn��#�(ûn��$�+b���QA��e�-!S�ζ����>n@רLEg�(Z�.���Ђ�D;���oF��k��C��Uޮ�4q�I�L�B$���z,[M��R5���X����Qk��H��|J�h�heQ:��K^^������a�Y��%F�[\z��/�ݱ�˜�ٯ�F�ʕ�7?'��T`|
܌��V�/���7��P�MZQ&�X�����_��h���ޛgr���
�$1OP^t�q�v���*ʐԦ�
�������RQ��lڛA���FK���޼7,������G��at�i?���Zl_�<��`�}{\�v��Cz�Տ�΀PWE�����b(��ʡFMc�}�;B�	�R�Rp\�`�#M,�[�Cy6r�H��̤��{U�Y�|opY�������u���P��S��jAO���Y8�"7��V���gt�D��-#G���$g�9���	��$�e(��ng?:܅w�^ƋՃ-8�}���_�Ú�?$�������/�F�+�Ǫ�x���S�n�_�ձ�YI�s���?[˾�S�~�y͈*�E���H/��*<�EҚ>I[II�]RG�.�'
D��CG`�o����&9��;(���6�h����b�H]Ձɥ� �f�F^��)�.w���mI��\����o�P ^����ݑ��&8u"v��t
���.�+Ӣ�kn)�Ϛ%�U�8.��{��:E�*~L����O-�۟�������W͍��Kc9,�كO4�o]�����KC	�Ξ�&��"x�4~4�#q߯��n����Nױ-��0~fVBT�L�}�]�D����#ք>Ev��L�΅�~w���`����z�#�Z�5+����~tZ�ē�y+5O`t����4�+�ި��:�mF�n^"�f���@�bU����4��p\6r7N��ySQd;�0�j�F����$Ʈ߂.�Kj_F���ј\�!�_C�DS����+�kt�g��ڵ齵��帴&���:�<3?���ŉ���#����J��1WA�L�J0ZL���%�`^S��h��	%��z���
@��\�:��>L-�� ����6�i��+g�����E��a��@mM�X��[dWa�e����M~�ْ0PH��� �=i�=9"@�'�Ȉe�eﾓ�b��!fK}?��ޢ�:s1��-E޸�W����K�'Xf�M����7��,T�6셇�|�#|�������[5����R��|;V¹Y'X1K������_��2��O�&�(�����0�#>8
A?zn�[��rKd&c*�R���"��횝dK:��Yj�ȓ�1��i�z{�+1�ϗxg�P>D�j?kd�G�U��m��,e��b%3yfƘi�a,��7ĉ���>į���2���#K��3�U�/�A����Ez��m�׽P�B�3Q��KL��w�)��{�3��JSU�q�g�#�I|�g04��-�d}*T��ϐR=7#kGWb���F�f�H�آ��)R(G#�1�RkDho�@��!Lޱ$�n�@���k]��J��{��	t�_E@��H5g�ߒ����t���!F
�x�A�Re��Q����xV�,�C+��#���"t6��TN��f��y�R[�{Q�y��sy�d��`C�F�gǫ0�v���B�y��M�)�7�(�C�����B�F�q9��Zc�MK]q䥨3�@!�{��1{��C ��� O�N	-�h��b�w8~;�/�Li4X0�Xo�l��  QB)����x�[Sp�k!�Ď�m�f	K�"�@ǜs���[�����}:��NB���A��a@svD���=2k��k�G�f� ��*��Obm��d�	���͜��nU��T5횯�C��N�JKt�a3��L����}ʹ��<�̓G���[���fꜸCP��,��� �2��z�7:9��-�L�X6���uw���Sc��3*g<"�~Lt(sI�&�B�"|�_�^��`x��MF�����x��'}G�7�$�8X1$��i�q�*9��:��
�ܙ�M��qV��[)A}�t�P��` ��lW��1�c��h���]�H7��hZyg�B���GkF�ǌ���?�|�/1��'y}�J4�T��<��@��sz�&g�\�^{F�|F�q� ��}�11��wG�$��E���v=em�<T1hw����;���
gj�M��p�tHFo4��d.=Z9Z�h8��i���K|�?oJAD�d�A���R����Gŏ)��u���c�͎'��C,��ʣd	O^~���u��G��4��ΊK�H�����tz��	9�����$��J6�S���+ANaV(�#ᵭ%%��Yo~��u��lZ��vY�oID�`q��إ�>��co���N���)�7	,�Lv8����秼[�]S����؝�Z��y���4�!�]���ἭT�B������x�knz�������U�q�L�B�/&:Re��Ma������6�-�5���ϝ���;}���z��	h��o��s"`.X���#FWl��5���L����1r��iZ�}�)��1c��{���z8����%����R�lCٰ�޿$j�G~\��o)4B�̖]������0\0LJ�$p�ש����@�V���z�����9�WǓ��o�G�Q:3G���͚-
$ME��$ڮ��_T����HG�-�e��4,4|}�����nY��(�4��m�����~���綮X���t���¦�FZɑA"��b�]��R�71�ci�f#�~}��:F>�k�6� "��I��H��x��Ɠ�W����C)?c�/h	a�1I�mw��%���|���]�O$�u����qA.���I�NإAk��4���c�BD�y���a�A ��&a�iC8�0١4����3�e�'i�$�q� �<Ǆ�r�6G������H^���5�Z����)G^���y�aP�NU��V\��6�����m��VSg�@ �*=}�!�0�i�<���yA$�60����"`Ǆ���(�`^���`�|���^�RY8H��huqc)KTn�Sˢ���wtM�K�[�T�z�����-��0���s�&�"�t�=�8 کu�P�=�|ť�0��2y�;�����Y=�?�1�u����V�k�_�8O�Fs���XXKG�7��LB����&��#���6?D�]��S���8&�㝲h ��Nb��@��������f�b�C!-E�?�LP����Yỿ㙯J��<CvШ38��w��Q!=,+}aG�(G�>����?�;8 �����ɇ
R|����^(�)!��d���t�Z	z�6���T�$D�4V,r�v#u��{W^�VR@s��uᖛ.�M��ҥ��+��p���H��1^*Z[	j��w�\`¼L�"[iR1sx_�mgfk��S��ݏyG��P�Ğ���:o��_Ҭ��3H�Af��~߾1dw���nQ5��������Ϻ�T!h?�N���'N��]��oW.wx T����A����oD^��b��NH�ԍl�Hȁ�Y�Td��N86f0������[�0FF"�Ѹ��°܍qY�B�ŊU���;�,i�
�0��|H�'�_�t5�*H��a�b�<�TM
�0W�Ia8��R�2%�}4D��݌���<݂�N��y�AO���r&.%��.�;t��6d��<��Td�L^��(���ײ��<n�T��)�Y�m��:��s��
�d��Y`P�p܌C�W^k;9ź�2��M���kLR�d�ݕ��Hb�Ҽo�ϴm�m��z�y��xF�UNg��lP	�{$]�ыUd���^-Z�T��	R��U��O>�;D�q�w	؁�n�U�����ߵ�� N#Sk.��u�4g�r���1�I��\ǁ�e��P��9:wV��c���5�˅��wZ]�Z/ׯ
>�o~��Dˎf�=���'�z�BpG�TI,�O�_d{�߬�i[j���vq�l��M���{^B��{�#!�����S4��:|̙|�-��3�N�sM�PC�w���s+�@��[e�jQݟ�z:ߵ3\��؜��
?1.�ǲ�6}���C��<���'���u�{K KQ&ۂ��eǗ���X���1q�H��<���Zw��$�:r�gp���;	/6�?1�#��U=��d��̡L�˿�
��YBz^���}J�����LiT��Z#��4����u֐$��a��E׽\`d�J(Ǖ�B#�Ū��a,��2MvAB�c�Xڜ;]s~G��l!»�Dd�q����X]�x�Mܒ��q�$�5ƿ/�:˟���k�LDwW�icE�E�3�չ�L�î$T~w������, �f<��h��<r�\q M��ڱZ-RkAz�!hr���ck8�pl��~�z��?(�P�H�?��.������$�@��\�+�t}$~��j���i6>����lE��dwW����~d�aS�u �~��������ʼnT��L�� �/$/(�����݆��iޯ���r�rz�tD_U��[��{L���H���Y��=Mjl?	,C6��t��ɖ�TG&~�:��W�����q)G$i�`����|$�P��t�mZ~$e�u�o�BR�9
�F�������]�����;�@�%�_ ��Bo�ֲ ��	a�1��i�G� �14*�T�NNǞ��� ��*�J*��B;NA�G�W�� �SE71('�x�8��Sn)����6��O�P�Z�k�{θ�hW�#��7�:�a�?\|Qs4��O��0��I�϶5W3�ӈoʟ��S�W��3���fz�����LFA�qH���z붨��{x`�������A@��CZ��A�[J��NA���������~s]���Yk����y�$}��h�F��2�	O䗺>��fH�����hv`�E�"��1�'��6鱙���"{��7����>�H�W��qr��I9gqON��Y`$^Kmbq.4���P�ØO�����5��@;d�A�1���(:
&�Lr��C���ٖ0�r ��J������x�s�yi��s`�nGH��"F�e/���V�w?�|<Y2��(��Ɯc�?e����co�K�i�qɬ��%�ު(�u����b͏T��'�U�����ݽ�w>bS����� ~�r�u�H|$u�t��V��'�I�q��L�+^�A��`��,�c�]�i��n���93Z�p\�е����	���7�
�m� �{���	�?�������~��%	�#V�$�{H
�|ԭ�R�(��<�[>y�w�ZX�ib��O�E����m����n����� H��G�M͒{{�x\������$|�`���lq��Ub;m,�-1�~S���D`e}����X��!���|^��6�;|sծ��-�('C��%"�����׍|�_��&��,�)�Yyc�K��q@���w�C�J�_j?'K楀����S��q�	͘��_�����}��!KC�O�-b�H$(CE�����E'-5ۅo�К�'9�W%h�`u<����s^�����L��ȿ�|M�v�F0�lo���c5�M�y���O2��-,,r�
>��d�^�5rfP�$ u� $�h�[6��S~չ	U�,��<�΀CQp\�p�st({zZ�(�C��u��B5��w`ߊP͵�-�0�>�7���S��i�D��#�c�d�f�7O��c�͸�<jQP!@�2Z*'gG�^�i;�<WQԷM%|p�5M"�;e�U"���`)�*I"jbB�1.�M^k���'���y���h�U��A
Ofh�������t�w����e�{�*hx��_ϣ�
�YoQ?;���/VRP�!Zz�C�k�|�Ǆ7#4#3���DV�$�q�T�\�iDBYQ�Ѡ�d�Y�:��O� L�( �S�p�K���p�}�1>4=Hgw�W�H��B��V.7��9Z%y����,����Ӊ���<�ٞe(*9�9B�Ƣ-�S����K�|�P�qd�	c��糺�:�9��9:�6�R�j>V�H�/�L���eIOA�b�x4s���ϰm��ݑ�䴾��Z�Cn+^g9?�	��1=6�����t�c�h����lk���l$������k o�\��I������Ya��K�I0Ӄ�K�/0a�Ly����u˖�g3`����T;��r�bF�m�a�,�J�\SFo����%O���K�`��${L�ܽ��E*>��ًW'��^�7�(w���څ�T�}���[ sy,!�h���<c{Z�
��PtzT?X�;QBQm��V������r��?�Ko>�&ƀ����t�VS% -�������Ѓ��h�ر\�r~�{{'vՅ�����hڎ���Jy�\�vJO����n:��d���3��G�߲¨������8��JBK�,��}VDjn�)|�/���h/n�_��__"yX�IR�O���[��Ҡߝ���P���� �m�I<k�z�ѹ'�/D9���e�3K6�n�[�������O�����A��Ŝ�I���pp�����ܽ��0$�Y|`�NX��d�0�Z@��ƤC�������&���\��*NW���.�V��M�s���uz����>1�lB
�a���`��c��v +�~���Ѡc�8oC��ذD�K�k���«%uS�%�.��'����YbE���Z���(�
�@iΕЇ���"=H���5_m���'π`�-�8�B�qr���$3�!8� �$�((
!�ljGD��go�؄���B�O��#A�:�QO3%F�L�� 	����㢷���vԜ[o;Eks�܊�q�ȏ=.-�ӨA�P�L��j2C����R�e�l�����smC�U ��G^@y
�|,
>ƾ�.N�~��bT�r��"��.�>)-��ǽ8�\������xeJ#��1ᜤR%]+j��Ȥ%��QY��Q"f����.֭��M�DYMM�&�����o�h�*�tָ���5.��X֓N�|���W��c)]TB�g!���,E[ri���K�����XZmB�
0�L���B�E����Ƥ�o7�Ѱs�K%��V
�+$��w&��Obw�����_ZfP������pJ�� �+��\3���"�ay�8�H�JQ�(�`�ێ�c�H�7�
U���!�G
ͻ�[_j%"�����$���P<43� �x'G�8%�A-_Z�u��B�N��E!5H�B)��˜Q��1JU�59����^���6�	����Ah��nY���ls����=OL�%Oժ+*4��+�i�AV^h���|��I�kE��V�҈9znfɹ���w#E ���L>߉�Ƙ��(�F��j�$ѵA�'?6q��!��0�}�`��+Ή	`��C1w��Nv�7��y�P&0t�w~���t8�*�bt�!Lj%�)7��(�9`��S.o"=�]����S̅ޣ!B�=���:p�XzO�8F2w<����L	~:��q@Z�:�"Cp�4Sn�����h5��t�IR��^ӗ������u�V��zA��ژ���Je�ϩ9���7�f�ᢿX�қ1�Ci�=��A��J��~����z��4%�`׮��B�6d��T�;Q�?��t�+Q��!� Cl��n����}�#���l���.��=�mt�eQE��e~Tn�y�D���F$�(�~��!Ђ`)��y������� ��M�!
���V`y�ٸX�t����6�J�a�m�g�����S���6-���4�OR0dọ���!9�B1�D���R"��N�|K4[\�+��K�$��rjݑ�����)q��e�������F���̾�����Rg5z,5�� $�/�w=�o;ik�%�ޣ���#�G�s?u����g��A\�3\�^],��a�:�z!m��B��򅑣������a����sA�s�2�MѪq[sg�L��L0&DQ��[w�J�6�����n֛� ���s�O�׼���t'6���3R�E�F9�M�)�1r����>[,�C<�f$B�k���8H.��O�+�V��+k76p�����& 2� � Bˠ�7ğ�E��N�c��//�`�qY�[q�za˫���oB�ӗV��=]���J藝����I}3_����<IrPc7�K�|v�w�:��*i��(�o'87�{�x��{���z�a<@�Y��	V� %R�JÝV@ȃ�1��f�g5NXy?p� �R�cM�ՙ� /W�qΟ��18���ɳL�Zꏧ�m%Z\c].��Cbؠ Nu�̓�8��� �Fƛ_솒&�+d�(�H�#ΘYe!	�p�z[�W"Ʊr��j���cj��F�?<����a��6�-ŉ�.몊^=��״��_�d�����}M3�՝#9�����p�,9�:=�\�|����~��ֈ~���𳲠a�n�R���RYZu+Q8 V�1b���|�
�B�B�l&`��'D5}����h(c�C@NH �d$�h|�"�7=J%���}�/��7����[�[�o^TRk�!p_g��8�`�'��������H��`Y�f���P�7�q����W{h@�ߐd�%�0o��	�h|�hP�b��.�r�|ǁ�Dށ���("�V
u�'=Y�v�)��v��շ����eH��ӊ	DDs���}t=Y�=�pjw`S��ϝ����|��-{�ߵ`�Dٰ�j�0�"�L>VնU��_k�X?�B�f
p��`��ЛҰ"2���e�>�ÜV��O��1b �q̱�ĀT�o_�Qo��l����i�JPl��@ڷfhj���G��Q�,?J\� ��]$8*L����GK&��Ʒ~�e�S���z%ԎɅ��W��ia�ޤj�6N��-T�G+->�m�;d��1�[����:��.c��riҋ�����rE2u�h�b��}"L�D3_� �k����/���?(����S��j�RD�c^}� Q9kY���m^i"f��ϹQ��=!z}�_��Z�K狆��=l��L�:�̒�i��2Y>�c�ͻ1�U���ۭ5kqAF8z�{�9,?�3���(�[M�u��0�1R
[�g����#�bC�F�fQL��Fie�`l�("a�&P�)~�<��#%K���eE���_��t9�.ɊU��O�)\:����V(#���%!^�9�R!�/�����$ju���\�@�vq"�"��\D"�1�� �pI�;�[n��|F_B��C7&���Z�r�zB��_���vG�I�42�͉ ��o'���`2�u�!̖ᕨX�4���W@5D5W���xJ�<��D�j�{vB%.�/�/.�$b �6q�f��$0��m�B4��k-����r+.�θ�)�R-\��^�o�Ѧ;)� ,�a]����w9Ǔ8�L�� �{cl�.��U��7�T)����`�m����]���.��ASc�`�4������H�Q��z,��Z?=�u��W`#�=gU�f��D���Z?�i{px����+n�.C��o9-7kZ������ku���p�~������?[�
&G�SZDI
��!f;�T9!�c&�,�U�������%
���aP.ݦ���@$�6u=���!�ś^�*O6e-�I$�i@
�3� �t/�9p5���r���gW�t�ݐ�]hd&*���6
椎����ݠL#x��!�Ť�H�MR6���|@R�ow��7�X8�Ey�gʩ+cF?��_�)N��?�_D�J	�1O�\�+)��A�	�q�`�Kp���S�����?�.�^2U8d��w䵈����%�w����*G?�w��Do;�=O	�MV�oe�`Z.׷ԋ�ɐC �|�_�q�}8#@��q��d���N��k隶���:2C��>D�hF�x��im��@��U�ϟO��`Y�w��"�u@g���ux��Ð�tP������%�{Ggi�u� }�L{!��쳽�p��S����@���[������t˸��N����F���ܢ3L��0Œ^x��U�F��@�[n|��X��?���[��e3�(:�o�A�ATn0�Ӣ�_�n��犱�ͦ����4>W�C��k_}dh� $H��BN:����⁝Xee���Dg�\Hp5.0̿e�NQ����z	��\$�2�f�Ơ;ۂ��<R��Mx#���5�p�)]��)[ 똻!���P�nT!o�]�z�e�'K�����f.�O���Pj��-�e�G�4�W���|�q=3��#Qn�4��$���'�û�����3�n�~�֌8�c1L�ؙ�z6a�F�Mw�h��� ��Y�����A��5�|�%���<Ά��"�ލ>T8����g�M~���ޔ
����E��:�Չ�4��H�۩����`+yٜ�Ue�edmE�D���
�ze`���"!$�Vۥ�qF�KOr�-���Z��Ħ[�XG��c�c����̓�I!���?p�%��6�'�#���:�j�w�J5����(�T��Fӱ��S�R=�B��9�w�wFݿ��S�	i0��o�R�U)|���� ��y6��d8A���(�^�%.����GK���5~�����>}!�9��5�G]����D�X���m�0	�����e�2�@�b?	��C^V�m�Iw�Y9��d�7��ʢƴ��7�[�^�g�9ڟ½j3��{�\E3�Zj��_��V��3���"`�v��5Jk��\�J	rM��"Ŝ	9=��h2jQ��<.U���Uq���b��U+�E�A:
>Y� �7�#�yѻ��7q6�/DƏ����K�ZԄ-Π��{y�3�<ň���B-3\㭂�Z&��r�ȣH�?�����e�r��P�x]�,�/p��|�c?�d�i�1�4�3�ݺ������$7��)̸�>�y�N�� <��}�<*���,0�~]��F0 �KG}��@��I��[�6���Ӻ?� Σ�
�܅N���!�}��o���r��m�ux��4�ޥ����M(�~�Ρ�w`zu�HB�oB�>��6`?g�'� ���"ܽ>�cDLʉ�w����C�1hM�s |ZBr�/ԝ���4N�f����s���!�x��_IPS�����/�,���s��#������x�u��۰�v���Q:�/�b�:ڐ�i�T���俘?��qyH��=���q�nV#k0�U��s)��7�zq�<�}@�-g�Ʃ�QkhA�O���	�o��>��/sVg�M+ᆵ��2YZ�[�ܒ3�� ��Ȑ[��|�H!����X�3&����e���w�9#�tu>�)�e)�ޘ�IⰠ�n�$ϵC�X�ǫ����:��	?������7�hUו�j�c.����47�j��*3��#�n�1k&q�<(Ύ!���*/e���$QJ��NJ�=����7v���I�x�en<��(W�oyzO)��";>\�HZ�8�F�����@�` @�meFi)�/�D������?Uh��q����� �Z,�
΍����i"i��\W��og4E�>*�Y�3"�&b6g�����͊��& �V���$Zf�HLP�Q/:z��?��Jd���e���<`���kd��+8&�'	�K��I��i���DD'#>C>��T2��>���j�叶�	�c�_#Iiz�[��2��j���xԾ�/�@���=Ĥ��Y~���i��}�f+�O�R�v��"�y��o�٬wɼշ�=���Lf��^�S��_�U�bB�	 3*
T��'�ϴF��~V����؏����U0���(d��e�ьs�^����&��=a���מkώb�g&����T��V+z+6��LiW���:j�~�	�|![�?pbb�0m�*-f�`��?��җ�+5[E�����8N������KI�o�*� � <J��ja�j�Ӳm�@���"m� A���s�mU�"�pX�C	F�@�<ii�t���[/���Su��v�_Q��X}�/b�����`��>Z���e���!w� g3c�~�������B;��+<(��*�B�Ď�M2���*h�Nkc�l�+E�ٌ_A�Er�P{���Tfxa�t&u�IО~s��_���&>n��Ո��dg�B�_�A�Ҧ�����'`�S���g�E:y��R�l':!��L�@ـ&~�UH�p��'�G0g�D���i"��"��f`A
Q�F�
��b�
�mr������5/_ϓ������)/���D�kT���H�R���H`L:�M����l�0����5��<�s������9��s��v�Ls�Yj�UIQ��T�������q̊�#�}/�[��d\&f�t�bF�|{+���������Y��Ht����Q:�g�M�y<��́�T�����c���*؄�D�iS�ሉl��gFlC �o݉��g)w�9A�d���m����1C|�$'��b�-#r���6�q>YT{� �:5p浪�tC�&m�\� ��-�<��k���yT���h�GP@��)S�2/��ܿ�t9?�M�e�����!ԑ���1 <g��;_�R�;�D�z�4�}��d���_����s_��E����^䆒��e�V_�C��+�D�8S��E���@в���TL�b�z�c"�C��5�Z����q$���Y}��4���B��A���`�͞2-\Rg
��i�!N�H���t��$�&���M�]���F�[W�.ܤ���t��kò�HW}v^��Rk�%b t�_��Lu_���LLG���rz,}�}5�M�}�h�.��u簹Q�O���<��و=��MumͪØG-V������L�oaר�o˙��R?�8w��~u]��4x��'�k��Dn��2��t���Rnu�=��_�5W��A���T����'��K��WX�Y��d���_�C	Fe��Q�OJ��>ʎ���N$ �M,�y] 7hg�-��
~���I?%��'<S�Ko��װ��k�8�׆��Oz<�qC���=j�p-�1�簘yI>ʡ���o��*�.8���)�oY/b����Y �bR�WYְ������X}�A����~e�]����T67�-Sl9YE�$�ry���Z��)�lB;��r	=���>��yjK�c���#�������s}��o<&�sXՒ��9�-���Q
���1"2�"��@���E<r7y�^�&���2����Ю~c��B1����^^�/�4�)�5�i��v;7�����+�������o����Fdv&%qt̚�g�w6��U�,����
��Vj3'��d��Ҍ$��rU������.Ӎx��BȂ���4�f�fD4���n�>s�"���3���Ӫ�E�*� hV��o������!�thZ�8 �#�Ӥ?a��x"q�+)�mª�]����G�ƙ���@�̄��ѐ
[��s��dl��J��"��#:Sng�����Ջ-?�(�~���ؔG;� D���Qs�Q&e|d��������C��}o*�T�R-r\f\�ԇm�o�D �@,�8[=݃����]-�84�d����*Mx���N�M����~��=b����;��|��n�ݏ�X�]�n�-���{������Y�'����O=v��.wk���4�?	����`����,�t�(�DX&$캹��ei�)�aKf��ű>�Y ��'-��қ��U��'�+vʙ�$�u�r�]��7��	�!�P�I�@� �+�ǵ	m�������'Hc#�ӨM����AR΁B����[�Ŵ��AM�q�qw�ݺ�6�x�16���U:w~1���(��1ə�Cѹ�.��̢�K�FI����c�5�x/g���h~6���yYЇ���Z#3��� �K�'��c�������8Z��vG����xE��i�q��x���4����σ�۟�(q��u߻�*������(���'�f|NV�3��{�G�7���z+�X��!Vȧ��0�U� �x���< ���A4:U�����s����g�JK�,=#�Wi�`��C
9,�ib�L�N��1SB٠�"��2�����4�8��ױ�8�����Ku�
)��~}��e�S���,�����pW�J����(�x�t��л��U��&)�`1�{�D��0�Xe>���1Cgk樚�
9%�v � �)���M{�y�T:�223���b�[�pW�q�z���hۥ;�oɌh$������-�5�F͇���)u�!��S:�\�mS�%�w�~����Z◿4�������>�H�/a�����8��1�-�/rj�)���:��܂�ш�M-T��t�x��K�g���+�ޙ��?eʬ�e ��if�v��T@N����q��A:���Ε>�c�t�g����-�B��f�K^�ß�L@'��K2�iaTК�z��SԶ���1&�Q<��y��_�b(΃��}9s��7F��C{���j��p�:\Wd�,�J�p�uƲ�"9J���e��CrƔC~��%�3� r��'A��d	h��aV�X1dor8-�](��{�;h��zq�B� VuT
�}�s���*�G�'�4w�K���x����g��'�z�N?�%�~!�mij�>_�����K�:��� D:(8��٘�(E��,Z�糧���W�V�4�dD1�\;z:��5a���4 ��z�����i,jŮ`qM�ȴ�=�_�m�13,�2�TZ��������}Q3Bk6l��-��c�	R�;���Dft��TC'�+�z�V���p!������)3����H� ���w�F}�?�[3i�z]�>f3�$��4��U���R�B� �@b(��
���u�t�`3�n�g��P�4��SA-��R�j��a�xH���4�B�t��_0����5�/ٞo�QpL�M�������սư�}:�������h6�i����oY�S37M�V��uP)to2Db�2�ò�=K�j#?ނ�{k���
ܼ1��		��A�]���+>Q���f���-HV�~o�� g���p�}�2bF����؃����]
@=�\a"�둄	���D�1=7�ZF�{�ڃ8��j(9��h;�q.�"O��sE�IɉS��E�aaa�30��� ��F�o��ũ�p��\��.\�l\��\���js��u��e�C�k�*h�J[c1�x^��P�lr�1X�,G�2fkw�_Ј��*]s�%A��TU����i-"�Pa�c6Qm��&tX˙6;77�|^S�v���Q��f��]8�Zֵٻ��u-�#-���;���!��6�L>'Z<�=͠Ypƒk�o��E�O�ި���Qa:�raq#�V���X�\����1 �I���h|��,j�d�о^=|�`JLYχ}��t��=@�BD�����	]C�D1$ꀐt4�!Om�ִ<hh�r*U��������s2lei���(�%����`�`\����0�s���x�\�@�u���H���T�A�AFM!>���rW�a��P�$���r:�SIfDnQ�gq��o�l�LwcU�[��\��*�K�B-�Uz��	}q���l8Jze,��Xr}f+��}9�c�͚򣶗�������N��+�)���[xj@!��ñ���69���F�=\�_��.rA6��Q�M?�v�V�ۣ�Z/�8�# �5cs��Y�	�� ���p�1u�j�Z��L�]o��N�ES��\�{8����kq�0���Π�s��*���R��:�zT�9���G��r�Ĵt�}���_n�u̵��:�+9��͆h���а3\���kZ���w�,@���=~�9�L;�;�^j"�,�(���E^�����W�25AZ��)oa|P �4�S�@�
��J4?*�T��"3���P l �yN�����F>x?�p~�'�k{
���m74x���,R��jZ����|�ohv�c��r�A�rw�2�j�OȰ�ɓ�����>ٗ���ȡ�,6æ�{M�z~�l����}q�Eu^��7��y���>��Q5�����g�S�/К-�*�����<�AȘY�0 ?R.�,X�r�{�肉���$�"!����'ɷv���b��<�"
NH��*�'݆���v�J�d��B�ϟ&�uZY ۀG,�M� N�� d�)��V]��e��2�f��h�uC�W��*@q�}!?#ڨ���m��i�9�c�����xZ��}$�<j��ESd�&�A�hg�/��*����Fo�!;�RDIAl#�ַ��MM�כ���B$h~(�����{h��x3��m���N��M!���L:�x/�mӵ�����$������ݼ|U":���3yT>����u5C�Բ�z��DXާ�D��[�7��	Ͳ"�X[�)��o�hz�6�����*��"������2�������]��!�3N�\�z��R�sYPv�W~���������>��DW+��_5r���esm����d��4픩�P9��&�*�fE���S��;�y���Z��$��se���ˁ^U�X�������'e|g8��������&�H���ȿmu&�)��pD�S`��!���u�NQ��y�l[���-=���|�!���ß�ꖍ���+����%�����:f�uX@����gu>�ܗ�<����]��z����[��nvSt�x�����;����h������}�	e�X�?��ȽtB1��4oi
�󇦨b�!��՜N��$��_=��*|^�#�H��p�-��C��+pGz�W!d���h�(	H4oÐ#�g�ɳ�t	����@������Ud���8I'ğ+8E7&���W?L>�l�T�1�VY��ܦ��ŋ���n�q,L�-�L�!�U����{k��U��x�[��F�ѱ���'qJ`��@�[�~��52��{V�G�f
�jq�!Q)37��g���7iqOE�'�>g�������ٙ���pt��K���m���*�|^&<ЩIo���2lrX�f'���wX�{��o*�v`<���r\������o3�f$w���9g*v�ҁ�83s���o�%�ң�|4�w
M�J�ohk�0� ���k���SމP��1R����%���#�ғ&؇��Z��߭'=��~{kS-���'���5�>hAp��gb\r�r�r��BG�3'�W� n�/w����`���Q��K`(�+�p�V*��qz�ힸ��Z�a����,��7�F67g���H0ě�����l�9�f��z��|6[���Nz�!�R�s��gb��e&�30�H)���-�F�Ӥ#��m
[�-����+�{�;����7��u�8b���b�coYt�O���K���%/�s����m��n� �m�A���	���N�~u@L�A��U/����(�/^k��MUX��Y~W��ή����p�i�8���ɹ��0���a)K��p���ŭr�w��3�����p�P��Q�U�a���Ҩ�F�=[�&1�G]�^�-0W���7���;�(�7QK��s9=-(S0�IjA>�!$10�����k>{[��y���E�Vƣ\�����-�˄���+k��w��̛B�k��b,r�3���ُ-���_�Y�� ���?�?.Ċ���Տ��we&��:���tX�*]�V���ϡRҬ1�p�P˄r=�XC��n�(�(�8�$)�#TSO`0F`2?��bDG/��[Kk�� (f$-���e��������M��rb.��F?�|��3޹S-<b�u�87x�u����@�4�O�����P�����؂�+޵�6z�R~a%V�^;�����ʡh�N�p^��ߔ��z�S8��L-�-MEeLT�e��2^�gg��55�gP�]g�^w��\��:��R5��s�D/F1nx���X-���"��k	��ؾ�`^�V�jSn�?h�s0ǟ��S����b�"`������,"-��Z����4�h��U�X)l�z�3yG ��J��}�\�knyc�\dޱ?Z�\�7�=!��O�����1��?�ny��I�	���PQ>�E�x5~�c\��$�w����F��&g����v���fz����@0)��)boƪ��"�d&�ׯ��M�)�����G�g EO�I����:�5��6��V�#z���q߲En��B��-�����"��_ �Ҳ�*.~���E)��)�n�f��Y��P�or�r$�h��d��������][��H�F�?z�F&nH�K�]4�H�U�0�ﺕ��-eIH�	�O��@�^�Z�94,�U��IPR�s;V�7�@�;7j�1�X���ч Sy�~x�M�m�՟��VT�v���+�"J%$b���4��S[�d�5!T��Qz��]G>C�O�]D(�e��dB���8�᲌#	����U<��i�S�˙�5� C��8�������Ħl�
�
����Z��H�gjW&)�<��{z�偳Z��:&�#��QX_�N!���y<����]蘾�탍���Y�gy���� a����*sӅu]���zpabK�jrX�jL��'�$#I��-����a��۶ֺ�U#O(�Q�)�w����0Keh��U��X��q�{q@�Rs��s�����sc�x-2=] ������#K���MM�ݬ����\���Y�����/�a0�h���O3�^v�#S�_�L��[�6�����T9��6���ج�H���}^�d=�6�p���ףQ�!?�QC�C}�G=~���Aw�`uj��X5�{ؕ�!a6&0K}g�;q#��3KV��'�*(<2GbE�XEJ���Ob���@
��"w�v\��搭�D�q�aÑH�ӟrrT$ԓ����N롬�.3�8%�L�پ�|��5jQ�d���2̠q��Ե�������"Z�����5ct���m��4;=B���a�`���Y� �	���pY^����>�f(���i��,p�~��ل�n��h�qA�����tݐ8Gȃ��|�4��d�cαy��;�ɧ	�e�5��i�;h�Rg�_�d��:]�K�@\�RhcCH�0��}�Yr�#
�`һHU��L�������;kZ}^y-�S|���a����XO�s��8�V""��d��98$�Ѿ"�<,̇����#c+�e_l��.H垿;��G����q�VX��
�(��?��D3~��D�Ud��Ft��l�vJ�Kfu.A�L�I�:͙�� B�o�ds����:(�#n���G�� uj����}KI@ ���WmZ�Mi��kŃ�,�w����D�5��'�`	/c�����)F�9�H0 Zq=`^k�/�ʌ�)g	��D����2~֫�x����
����d p�g�=��+g�o`�=��8n���1�<�nW:��La��Wq8�An}O_�PA�������4�����ʛ�*�/$Y��Oe�����.C��W�ſ�j_�A
�&�k5~��u��Z�T}=�jLDCN�ǚ��S�.�^>ީ华� ����y�J�m��R��aq����i��(�=��l�|/'T�e�Lt����gp��fg4ѯ$˰�A��9�H5�~����ʭiF.�Y����W���>����[s�z�vf�Ҏ�3��y�!���ff?z�'���֞�hP��Ȍ2��R��Gօ]�>%lQ0J�F�K��M����|�w�pv�Z�p"J뒽�L�O%��s���+�CH�T̬�~����fc�Kv�p%�'C�+�[!����f3��ǜ��bl,���n�?[$џ�m�"N�]GFFR��B���##}��W���Z����"P��^D�B0���
a͍,Jy�T�8��O��M�s"�@j���FI��EfHK˺�(qV�>=^�ˉٽ|T�[w����f	�3@i.�u�7��1�[���/�mOBA i>Rm,�S\/�v���#Т������pi�+1ek7���*�_����%ʙ��G'D�r�S<P!J�`^̏;q6]�[<���S�_��9|������^B*�p ��H��'�=j��H"=���/rJ�4�My0b,�T�_f�������h� ��x
��5���Y�`,��!������=�d$�i��,\d�yr�5�N�Ψ0������㎩.���~,��",����O����R`Q�]�S_��)��R�/J$tu�^$��x���o�?�8t8��k0�3dd�wP����d"��48����r�kF2�w�[L�P�7,G$RC�d�p�*l��8.R	4Nf������A�$j�v��UU;Ev�w�������Y��D7�����͢p�Y�e������.?l�����_U�sO�$����=���;��Y�~u�D��7���3�u�|,]���|:��%�]���Z�v���ř����/ō�g��w"�nWIS������1a���q*�����e�`v��D�73[��V�V��6Jq��.��zΜ��)mIF�'�L)���w����ç6++��a���&��e���o��v��{��Şڻ,��t_v��{�Ղ�|���n��O�%�AMi�T7ș=<ɖ����_0��C�ik�iY�w˾�1a\�i��ð����Q����٨�|��>A�uV߃�
c�0������ϯ4��������YQ����h��j뗇Y��iEv����h�����ˑ��[����F�2i`D�� ��*L��j�k�0l$]�{���$]p�Uװ	T��b�5솧�� �nСs��S�c����u���0*&J�3�d�M��{�D�$�����I�WӿCm�˓l���]��}fӿ��y����ՠS��D%�9��:�ptE����@�^�R�]���ϒg�Z��mRɵ��a�s��x:g�Y*�R�^�U���xhh�������$��h��'Jl�P5��X�L!5�&���'��D
�2�,������Y�.�n��ҧBs� �!"��X�O��Igi����g��o�r����Һ�����y�ƻ[	>�^
�8�z�&p!�煮/����K�w�������@��>�Յ�*~��'@#H�Jq�T���؀I8����|<kmy�;���@G�a�DX���|9�PqZͱL~�}Z���_��ȱ��	��.7�Y3���؆��2+++׳���Mc���\*u�{XO��`�Xq��{U��!��A\X�i6'ػ�ޱ��(�Y_��Xr߃`�U������fo�����0u�m�d�N6'��S�5�dL�9a�m۶&s2�����w]���^룵W�A��[̨��#�!��8m��,z>�{S�t:�-��#�qߩ#H4+ђ K��k��J���T�N�E���j�S�'�˙�&��ƒѣ��V�����.��8b0H�(�)�d,ݝP�$LZҙ\l�3�!!���
`>�@Sj_$��h`x�
s�e����dqBE�r���< �іQ]!!�G�r)�z�P~�cg�?8>B+^/�]:���A��x��Um�
��a~�ၐ���:q��`e>!�9Ů�n3K
�&���JnP���{*�ҩz9��8��MUF���*��wC�0I�P�꠺E�MW���&����r[�Mel��:2FlP���Z���H�|c�W���Ĩ��A)�gU�
���1�L��q)����SP�0�X��!�,���~�R�T<��t�db���毕hQ ٥'4�p�Q6 �RR�/��ܝu½��K��D)�|�:��D��M�Z̒�H��JVi���ºKu��A<�̬�Ve�{�۸���3�r�ۍ���&+�����l@ߢ�v�p˧��p���"ez��+����'�j�� �-�>g�jE��u�#�_B6��k�q�$��R�2�גe`В>��o��R�M�h�0��.K��S�28&s�?�F���s-}x<ȶ��ܔJ��Z��[}Zl��� a��6-v�\o��'�0�[.L�� ������f��%�x뢟7 ڈ �h�*���A0b(� �d)V|r��K,�f�j�m�&�玔��*���N-ϕ�WM�����є�3�#�(���$����F28>���b�8��Hc6�w����:jR����v�]�|���f��t����	'~��\���?T�j�|r�y/�������ڕ��-b�ye?��'?����O���+�M&����JlV�辏�q*�^l�
�)���[.�����A7N���I���;����B�9�^���FH'�#&YNw����%< ]�b������Z�x���tL�D�a  �z��0E�WĪ��9�Y8�p,
���5ܕ	H�w�=��=7��j�]MYS@�ْ h�l�p�)�N�6�,��P�S'�|<�3;m�^�����*M(D�-g��)O�O����PL�X�Ɂ9����ĭ
�;e�)hݴX�iR�"CsX{�J��qJ��%��^.yl�����h(?~���u@v�,K�*�����zc��z�n�"�m)��99�Ws� �H8z�/�EE)Ξ�H(6�/��C��5m]�2O�i�~=��	�#��:ɫ5���u��c���F���>H���h+&�ƪ�.����<�ɹ�p�w:�_WV��IY�"֕����vm��$(��p5!e<Ñ2�9����i�~o���_9�J�Ն!��eK�d�v��td*<ǽ�´�SX���8�!tJ�\�x2�/{Z�ܛ��nhp�d������ �hd͆��f�pŧE�B���=}�|��|3�ݐy"𥟫ߧDVp�vmI��|�3��\BNk'-O[���&��!��)�0>MТZ���l�2��4��6���r+kݮ��:�ylqo��$�~}hw'��g.�JE;rh������{�| ���3�a)C�h1�z��q0��!��/��m�e��|�%w��;�����
SIɵ��Ն�,I�@c`8�F�Ӱ���gP��-5-=bP+4wZ�N��_���TG-����:_�W�j/�F�cQ�wT5}H(ĢU��o����-{��M�h���ŕwQi/��6,⢧S�/Y/������)}���&ߒ[�FO��Q�7�Roݧ�(S&�M�|�%�P���NW�[
~���q%,u9YH�C���mC�Ҳ��s๓��S@��X��p`5�mQ��z�y���!�\�.�:5��A��5��"��?W�v-l�\f�-(VU�\�}���r�5����`/So��H~��dt����W]u`F�E\�$`�`�!����\�I�$T"كViܟ%osX��?�R���x�Z��(u��F�]�P˳��8�J�K���7u4�w�r�m�!�6AGg�78�Z�X{dR���X&�T�6�VE��d��^15F�o�=HU&�/
n�o-�iSǢ�xҢ�Y��7��ǡɊ�w��|�v�=t��{�t/]��I)V!.4�I ���(����3zM�>�]�}�r�HD`����xc�6C������0[�����Ϗ��WB^�S-�c[�tMo/�0�L"�՘������q|0�R4 �	(-����~�*�H��KN�q���� ��i�����0�aQ~Bz�Cj��o��y���*��/��K��ս�)�_GΡ�v���"��u8��8O���#%�TP��D����fy������ ��aLC�]������ސ��k�N�F�>�]>�C�㞊����,��'�V�6۹�i��l�G��?�,�1�>��{-¾#0�	�2CQ�5�y*�(�']��w苮���������f:�r$A�p0&l�����{��X�r�ٛ�a*aE!β</��i�(�K*�79��C`�F�
uɡ��`3��=��-�
���
����m���/�� J�n���yH�D��?F%�l��e`��+���e=��-��jB��0fT�A*$�D(�J{O:\B�gҳ ��!�޾�V�&�D�A^����~�K�n��=T�n��� �0׏���d�N��ih�m�y�4�
�G���w��������������%!���(}^�[���I�� K��`T��|����(s�	GZ�m�z_� �|jJ� =�)�c�2����NX���A����Q!b� k)�V�p�P�iFj3�
���W���'s����k��hey>~st��~�oM�UCi���)p�g�I�;������J��b9E��l��g��6��
M�Z��`���@��ϙ��j���n���)�)�Ը?"@<��:��g��󾰲�:U�<��x��H|w*"�^�[��XT�^�^�p�C���^a�pd�ס�~��a쩇qwd��e{�'�	+k�U��{[�����g҆=;�%͙p<�[�}���Ks�h��?x���E*wr�W����+230�&��[��i���;��0�8Zk�JgJ���6]B�~~}��P�E4͌�6�K�]�8�ǁb2x��c���o`G)���Ҹ���0c����	�x�HT�*R.��ͅ3��7�@����|�w������ƹ�VE��J��6�����7Z�,�� ��7E2U?�C�{���鞕B�i
9?���[��'�5*�)C
��gh}�`oYH�w�3��k����g��hY�Z"��̝:���?��k��k��OK��`Kz @�T�I�e �����[1�ZLDĠ�~,�������P�R�?HcH��q��^�(�-=-w�o���H�)SC�W�P�hsq'ȮX�B�F�p�t���4mQH�K:�g�O�$&�Y��jS�Xߵ�A����(�q��a����B
������dA��i>."<��b��h�H�}�w��f.|���ˏq�K���L�ކ��|Y,#z�9Ö�p���F�>C@wL��Uro9��a��|�����Gl�Z(6� s�&�kM� 9Jy6TԶ�����;�`�Rه����n�T:��gr3݁uX���o ��Z�[�Q�F���wS���FX9�.�o�k?/��]��xp�� �!�:����4���_�$��K��y��`���v{4+%.��$�����i�6L���O�E���\��k+l.u���r�ў�qN�����z���v'-�\?�_�@b�ϯ���uV�.g:��II7��\�;�'���˟tcRm�Զ��~8��	4=�s.��6�뿽:֔�6B��"
�d�����3���f������(���Q���!�h����*n-dotQ������j��RN<H
�^�F���V������'k�K�3_R���<��L���%m�h�1��|�i�E�Akq<�K���5<\�x'[𙎔t�D虓�咈�P^ZT�P^�I0I��j��H4��}"e��ٷv5�:~znɶ�[�h'*��Q�c{N���=W �`���[#QF���dC&9F�#mr�,��r�:d[���WX���]B��o^�e<��"����NKe���	�Ow�Q7�L(C7��Ip'b�R�],�X�GABh�\vHi��?OcA�54�L��.��%a�V`�e��(�V>�
�D|���c)�����W;���=®6�t5���$B����
&S��?ɥ�L�m�(�v%uԻ�D����ﾵ���M� J3��q9A2�m�ՌѸ�|� W8l��n�������4�N�4�^≇~�������x3�E;�w�@�00-���w��=�JiM��	�"��r��0����6d&Ȕ-`�����ZZFf���5�������סV�(z�u?Oe�ˡ�$�B�I�^0��F���ݟ�"��Ȗ����Y 3+�z�����Ua�)���7����g����|�Jdr�
��d�vQNڋK�&�
�ƨ��V7�����W��͋�x�KJ)�#��Y)s�mr��j�b���Ԥ;}W��rE�T����3%_q�1|�q� ��s�T鸬��Z�c�~:&��>��f'9�ln�Дq�а3�aQ�fh�u
�-��肂�"��׹��{c}��F1�X��_�#�/�]�4�?���0��Ƣ�/*!C)�Uwy���9Y<zP������yZ,Fd`ڸǜ}��D,s<�l&0±��8V��j� ���{�>�A�0�5���>�4#��Y�:+ݣ'|~6����|-B�÷j��'*ƮN��'�&�_�n�E:
���7�|�'4c��g��Z��f|�[���X<qYDreyc���aR��
��8Y����#*�SX��F {�9M�I:(v�B����=[O�-��$�[^mJP�tZM%]������!c!j2��y8`�b�F���p����<�qs�RhM%~:iZ��x�Ư��
���)�� �F)f��\�ˇM@l�އ���|$.G��vA4^�֣��I�2�@��s�{\�8��]�ǩ�Կ��-��^�NZ��*�r��,�j5�5F��~b��k�[��h��������������}V�@�V׳ԣ[�XR��u�S���݌K>k?�	��ڇ��1|j�%��'���z*��jItzK�L��ɋ����|�h����'A��v�>R�'ti9�&�ic�=V8!�> ǜx�O�;�@��-����x�Asn�]�M�$�%ξW���H��Ѣ5a49]�Qw^�e0�����ֶqՏ��6S�,�S���M8�N�iHz|�r�T���l������O�>{�h���Āoő�� OBE2��B��(V���!���J���� ˶Z�q�+�5pO��/� r�&�����Z�*0��ù������Y`�u7di�!��Vɹ�<�w��ӧ"�M��A����]��;.Y߾�#�H�3<��L?M���m��	���rlX|�il�H/����a���Vi��ZR�t��Ȧd�]����4%�Y,�\�{*��r̀�=���1X�~����Xs����tL��mz�O�	̹���L8�/��rpt��Xk1�p%��m �i@��:s��j�R�Ob�jY
v�9w��%%	����ƻ�
���k�p`�zx:��fW��e~���*w!��p'$�mۅ��P-�S��i�����=a����$掇ɥ��<��� ��h�3�(,�%J�Qi���p`��r<���sZiq�2{3W,�r�x����B���|8���.�b�\�U����ȩ��R$��P�?�C��TYb���@Ɇ?����T'��'@�x������j��n��Ϊk-MS�=n�5֟�Y�g�g�6D��v��R���XWWW�����'�f���Ax��֩��D$#'��%��uDnF�U}2�(ZS##�.y��a�tf�~��A � �@&r\	�3a��|\6*nP�Ƀ��)�Rs�Ĭ�����t�0��{U�"š�SMEf��QJ� )��t��y�ӽ�/vu���]�Ke<�WUUrl�k����s��dL̹����]��c�Nh��	G迆����vOɆ�w�EL�6�5�_U}R�l�����h�Yu�sE���w����ňq��R'D���f���~���m�BI|D0qp�E������k���9�}f�Ѫ!A[(��>����ɭ��~.����^�#CQ�h�>曨�[[K0�Vq�{U��L�Ok*�
�ޥF�^��

R���	�����x~1v��/Oz�;�>��v�z!5�j~��j�M.t� +�qƗyE٘|B�b��Ԇz�Ó� �b����Y�7ܞ��ҝ��8�G�4��}�Y�l�{$,����o�^lv6Nj����͔�����_V9���c�V!��q�8��cg_��R��+}_K��n	�ͳ�����č�&����-�7�9�N'���������)]��~��GuY����a�hv\�br��4�B/�"z�R���	���9��~� oJ�g�*��'[�3!��ZQQ�g�mcx"���V���N�NE�y�n��gkqj�ňV;e����1�	�l�X��{���R�u!�������6��C�R$�7�ss?j���4�뵉�|:\[{����l�m�,\z��x��j�?@��e�lP����Z��X�Lԉ�њ��.��G,�T���>M�Z��|WLU�+s�m��3�n6D��
�[ٗ%_�vjF�0R4�⌧�yB�^�5�H\�7��Mϩ�XD5�����O�:X���޼x���s<��1����⟫�����5T�����`�*����S�C�Ƕr9$(qEv36h"�J<P�E�t���Ls��jC9!��s��_��[� �'MK�N}��mKA���0پo�f��D�b��V��8P,:�EX�����-���L"�q�g�z>���˧���`���)1�3!Ͼ�����7��Dz_��Ֆ���>tc�����<E���G�\0�T�t���Dn|zLу_�q�V+��!��ܗ*7���7ha__�KXR���H���ѓ�,/�ּ���'�S�~��"�����yX��n��x��D�/����ޭ�t����D��I�0�Q����.��sO���E8�6�?m��n8ߟ�����niѫ�ʮLB��6��n�MLL�P�yo��%�y'� �}�~�����SXx�&�?�wp�G��OM�����|<����4t���1��Z��p����L��5Go ��7���Pw��0(�9�C,Y6��n��ў<�ӯˣ�V^TblM^�12�m��n�Ԇ�(��[�ܛm�����J����C"6�����J�����t+�]l||D�3P���kL�-6�.q7�?�8WVy�5�����.��v�Y�S}�Ӻˢ����\&$��B�u��t�2�º:���K���^�3/�lI\�]��;r2���Ҋ#7�݁�}��� ������(Bލ�&frr�F��Q6�:�nl�6��}�[�/��u*�(M� 9�
�W˙�
��|�`��蜞�����rH�lD'��6� �|���*RXιf�W��@ҏ0.a�[-��1H��}[SF+�~�`��Va�'D�x�2��}�A�ߓ�Qi�7�Y)���e�f*�h�wZ�����p�-����Q���lq�l}q��*��˓���L�a�������ϗu�YMk�L�Ǌ[߹�<��|�z1�����h��8�c�Ǽ�op�d�ݶ弜-z���ߚ����� �K(1��~��������L�v�Jd'M}�MvR:ۈ�����$LG;�Ɩo������f0�O���UhĜ�"TA,`o�#��
�Z�
���K�'s�����)1�.�t�'9�] i\-F�����@|�4�Y���|�����עL��U�K������p|��`����%l48��w���k��4��:M�C���آ���J��Bn�|��f������o��޹ڵ˞m�����c��U�����+�nM��6�$X����m�^�Y$�朆��6�9�-!���jC&�,o^��I9���J�I��n���Ug�8*�UՏd�4�!�e��E
��k�f�����(��"B[��3����a~4m�f���8e��_|�Vsƕ�솘A�َ(�UG�e��h@����\�'豱*��?d`Q���.��^���~qߋ��G���E8�ъm�KL	RZ~�,.�u��Rs�E���eg,�(�-�?�M
�ϵ�	N�#	҂٬x�א�~�d@�XP��:^�v算��5  �?K�}�c���I�~��\��%?����~��iRb"���[뺂��4Xd�
g��`F�D�fx�r���T��kD�]x3M݁M���gSӝ�0r..�vV��r=:�g1�;�T�,�Ram_�[���C1��7y����~�����}3o^���hi��S23�Ŋ8���Na*0"\��H�xڂ��g����-��O��Z��qڶ�_N��>�4�X�(e��~,<{�M>�!�����.�(:��OT��IE�s��U���+]��̾E���Zkv�.*(k��+�ϟ�/Y<aQ�P�S�e��������@B"�y��/���U�Օ�,h�(���~��?�W�q�\��}ޞ��LZ�=:v�S,��J���&r��?�&��h������Wl�z�l���꯮g+��z�-�t��Zk�p&�]9d���q3d�C�#*�:n�	�W+ZZ�o�<_�#%)h�?LC��U�j��y�`c�յYm��,(裧�خ������'>s�M�{������Ĥ�a����O��ޖ����+��A!Z1���@U��d��5OPљ5��K�YIq)".+92�ʮ�$��i���''���J��h�X��Uon�&����9f�,>?��:�q/��ie_���W%�`?Vb����S�,��ÒIZ���G����>[m|=}�=�h���mŗ���0�C?����<O��]�]3%W��i�����+�����Խ��Z�ۮV[�U��r;�LH�ˋ��8���������6�j�w3�qY�3V=��BBP�L��Tv���(:'SC�ӭ�斫�<��dn��-�z}ў�k�Cկ�Ϗ?*�^�]�7y�9�X+!/�M[,3��g��i�Zpa�M�����f������J�]��yݤ�|�7<���NP�̛i�M�?�?/����B�(�/��/��<N��E<�:�i3�b )�AX%e�֒i�<�`�B��W���ޣ$'�a�T�:������3��c�ܐ�9��#S#��2~V��{��x^�s���و���8� s�\��Q��Nl�&��<DL��4�t#_�1�Zo��y��sPz-#�~�]�"��-"VɔEPݟ��NlW~8�����O,a�a�T_5l���Q�����q��!P�_T������􂜅g�e������54�Z�V�g�v�^�`�t���DV�!���zH�@��~�0b/.)�jhL�Ԃ�.T|��i��lT/Ո��$�wS�x'�."���$	f�`�v2eVT���8��g��(����q�@�T��QՐS�������"|�	�o��ئ�@6t�݀�e��vm�	���ÿ�h���N�檪�󶶗KA��b��{(+�z8�5-�����W�l��<��é�^���a\��:Jq����}���o����b�
Ȁ���a^��\S�=�����d��������o0a[��D���rl�q��?�2e�Un&B3��ģ��0��;��YI��u��M
	(�	�,Ӻ5�
s�ruu%������)�⎍S~���6AL����ȇ��;M�~��j�^�	P��<�hʗk�]�-F����6k-�)M?�9�6:kPw�A�2� ������zu^)�[ľ���6LT�����2�%�z��B���
�����C �o�ْmEY�T�,x.�M�Z!��o䚴�F���qn߉���3��ت�n���j�P�!��hcUR_9�o���� �U@�}*Ol���Y�=*Ѭ�"�ΗB��!{����jq9�f1��XJ�������[�ճrv/������¬Fd־�2D��Ze�Ƭ"	���~:�޸�tS7�#Ytk����u�������Q���<�F�HHrt��oő���"ɶ�s'k	��JJu��{�(lS�6��N��\@(=�u�M����A R]��>;���r$��H�����V MюNI9d>�8 Ν�#xuϝO"�m@�"&d"���ǭ7|�|'敋�+�wT�k��'��I5KM��}}}�D|u�������ճ��N��ܮ���}��ȥ���h���� �+��g���
p��cR�6�fL"���I+�]�af������Y?s�1n��S�x�.TH7��U�zf����nx�\���r��wu��*�F���R����ߚ$O�Z���$w\5��d��1�d���㒓���Ґ���:��M�y+)�:�: ܬ<(��i�1!���؊�">j�>��<C�p3e���}���8*�g��@��SBD���8 \���m��l˩����vѭo��j���*^  �:��������`��%F�Y���|xp'�&%�M5�E� Ď���%f��XmR�+�)A��R�����#��B^K7ǥv��oG��4P �]d��ceI��3��"�M&������z��)�]��n�y8~�
,��x�T�W�B����Z�H�b}Б�f`�=(�pn�Ť�*ԟ����*a�WFEK(�b
����C��Y$�TNuU��3� �8��z�߉�����O.̴֛��0�E�
��^�[|1�

(�y��G{qY�D^���\�{��}AI��}|��a+�����g���U�����s�
;'=���l`V�h()Ca�����fiWA��fff���0���l���P_�'������]�8�+�J�������k���oʦlI��DC:}��=�ꘘ{_�>��
O���p�^���!�8�E��1((�]�ז`���z��l����l
�͔����������f���q9V3�+M� �kwݝUvX�_4H/���|3ՆJw��ׂ�@���v4v������S����1K���,�"y�5fr�9"P���T�Y2�}'�1�^��c�V�^�~���WaA&���?��C|,�����o<#�	�VUM!�At��R�Z�z�*��\������M(��-��$w1v:��7Z�f��"���~x��*S�l��ﵙp!���v��M�Lȶq�qʒ�4wXd�˵ ~U���*�"�p|J[��u��J�J�}`P�1/��GaA����|l��߉_� ���m͵�ޏ�1|A8���r�?*O�!A:dg�B�CʟZ,�I�&ox^d����1�@��9�jf�(�LY���e7���]EG�{��)G{�E��e��l�,����+L��X�E����ϗ�ʎ'�[�l������Xs��R@u��߯�U�M�-KH�� U�!���h8���ڈ�"�+A���f��l^}C"�k�f���?��>�~���ܯv���L��ͩ�f��˚���go`Ё,��(�X���+���4��^���T��S�Rg!i�yV_�4~<�R���|E���<�0�Z)����Q�XK��p��R0�><<���|G��ͭ�6��|���J��;�Ü�3m٦��B����{f*��=�o$ܪ����پ��CF{{{3���߾}?[���-T�����q�	�/��/�aaW�+�3�NL'�Ō�c>��M��8��Gqyָ����������{O#�M:���?O��V�m�Ս��!oK����e�<_9����w��ۼ>�Q��W��� 8H0����uh?i��hj�x�]Otq6�v��rr�����#��&���^l�+i`�Y�~�mȯ���?�!���M��c�f���c$laj`��9,����ۓa"f�gB"~g�ǳ�w�S�2���d9��O��Ӎ/�]{��RY<��ek��^:yj^�oQ2���C������钽�Iؽ��CSƋ�n�s���0.�X��JL�+˩�W�wz�|�Ȭ�d�e[�,�f�OAt8��c$��ڴ���FD`FQ�2Ej�e
�6�z�'��$6l7$C�X!>������Bnz�럮�u<w̛ed;�,���`^ط /�֋L��~����I(ff������A�<V�����"r��w�d���v����drQm��OC�J��@�Kf�v�$�2|q�cHr`<������b�Wh1�N��Ìy��܁{�%��lQt�tsR)Eğ0aJ��%@@�@��)�����ÊM��?���8���N1^��.:8xǶul��6�F��z�ԨH8ل��������\ �?� �fi`�u��6w���X6�h�9��|ٵz�8�k�������8%��^o5ޯZonn���L�l���*�u�PH��l5���a+��_4)e�9����0QR,���PB��x�u�D(��VF&���r
�E!$$B��X�Ǘ�TC���۸)��Ǹ7���� o������\�����~PPP ��u)Q��n��X:e���4Sᬬ,�4��Q�΋������e(y\j����N�!��b0��[�-�v#�]R��ᓝj�' ���Åʎ�� �6�C��a��l9K��R��U)r�og�̵�4	i2���re�w�[
��ζ=c)�;9�����c4�uNZ������'k���RN5�~n[T,���epBf����u���4{�^����G$iw�����>��[���ʶ�n����m���w��.<0��
��W�4R�c�ɋ���_!�M�Gd�Lc��Y��Y��c`s�=�X��qle)���wZIII��%ㆲ����'��M�q.5��4}{�����Jl�F��u��D���I "x�oaf̌�wseʇ���sX�������%��ag�:�rџ���l�����o:iv_���k��r���IԽޠRɄOPEezai)E>S1ۢv99����c����X�"��|��e,�2c0�f���e����Yx�?�@sBRH��J��e8� `P}��q�(�om���Pc�覥�CSQ��hv;�Z�wӗT��>�3���wo({y9U�`����Qf���A2�l��Y�G�o�*���Fi�����UK��M7åX2������mo����� MFTX� &F{���*>�mFfFF���NßP��x0k?�q���Y���m��%3�h�Gp������@]�.xL�x��7�v�R$��.��=�ϡn�I�ώN3�#"�����k�	Y�� ��Kg����AӖ�d�>���>d���=R�%�~j~F����!Z]�Ɉ�6����Tk1L�5yun&���՗XL�G���yTID`�V�8�rC�������������`�� ��g�ڄ���Q�(F�6���B�D1�ֽ\��lt����?sp����m���TB�5���#gj�a�F�0e�֚�*�.4 ��ڏ�Δ����0ܢ-�ۨ���.c���b��~����Cu>�͍�`�~���oopE�P���Ў���k���R�h���D�����:5���Ҫ�?op7�KKM�t�ɽ������:�!���~���.����r�ˉr����������.�ZD��[i?�xH�O;6)�U�_��Y���9��Q?�-�&d^��Z�m��k�oSs���S��mT�	�&�����
ƴƗ��/�C1�_n���<~�����W5= �n��ƅ^ofkj�z�82���v���K�N�C���QhR�`���j������rΣ�9�2�I,�~��V�b�_��eJa��8�mL���g�:�J������%�F�'y%^�Q�C`I���������E'(���u�;�2�F)�B
9��Xdh��<�ߪ��� q�?��7����J,��'���dI��.6B-��]�$J��ĥ�U�"��r����l�
��>�z>�bN�8*�2_�R�<�l�\��6ȴy�����$'&�4�B�q"�I��P�'�P&��<Qa#%�:O���B��G\��>Q��M���Z������!:�(9;�jS ��S��uꚚq���S1��ⱋ8���b�:��'���5��98dͺ��ͅ|iI������� ��H�2�۹8'.#� ʹ󘱷��{�l���"=�׻d�d�m���R+7�Y׹���)n��}�d=1d@�_E
��n<��xmt�@J2�E&�"@`v#�i�D��x����ţ��5�4���jVr2&JJ*��ϔ�MM�0X88k/:Ұ>v,��s�-��v�:�+;��<�&���zM����?�UNDM�ָ�լ���?2fVl�d!���B@�'�RiEyV���s��v����
g����:��߿5�O��DCCwiU�!�`Pa'8�P���*�=�2e�/�I��y̖)�̭�#���/�^������ ��б�-����������H,֛�F
vzpv�nXJ]v455eW4��+	�.5�����+ϐ�^��U������»�!''�΋Ծ�Y�1L��}�{�J�*
�~�y72���#ǈηe�����Q.�ui��1�>���-���N��ѣ�q}�����p���c�݀��("�"|�����aN���������Huo���E�6zA�C�U ��ZQQS������&*���і��1���\��7�|FN���';R���~K4��nP�O=� c1)&~��>R�9�<��|��/��e��?��(���L~�~��I����C���;����ȓO� �fhH>8jd���p~mC�@JSݷ,�'(�2Jh���_��e'������>�qf�������.�jA����������������=6S��a����D%.�喉[z�E����൚�o�:�@�`��b�o��)#<ƻU趞3��+w�w��%4H�e�^�֮��^Bp9>Y���k�y.�.�U˗SUU]�Z�����L�D��J@0��&�g��7�aH���+U%�ix
B�a3�Τ��"Z����o���|�{��(;�{�*#��H�o����$v*�.f(�jE`����+Ld1P��y-�7_:t�t�sE>������x�5��X#Sr��nq��J�gy p|6�_�7^9����Eƍʓ���o?U"�D��(x�M�A��]{���,�5y� �̕X����g����_|f�I-Ų?}��I��<���C2�#>�ߑm���C;�uw7�7=5�d��5 �޸��x��/�L-E��KĠ%
��C�W��NDD��X#�p��[�u�8�W��]��E��\~�c~t 9���ę��U�|��W�ٵ55�����i����4��01��j�i{(�o:��O��n�q�o6]�n��o�3�e��2�J�Ėt�� ht��]�3R�?ݹ3HmI������$eI�#0K�؝�����9�q�(c	;J��NM����,Bk%rc	J\F���w�顐 ?����w�m2-�X>|I��귝8�����F]~_��k��%%��#����I?�m7�2H��)c�O�b���1�gpb����v�2�wRq��
$�y�dr'&�$����6�N�L>�}�С�v�"|����$s���S7�6rûy�J�H h���B�)S=)�q��`��\� g!$4�	q#�%/�KA�L���2��t�RI(��$��Fde�=���Ϟ��m���k�U(bX_d��j�b����^9"�>U��x�'����_@>���e��UI��=����u�����W��p�_�դp��Eֹ�����r���Ŧp�B�kd^�n_,�T(0��Ј��i����zYQ$]WQ����F.�U���Sd�����e�0����i��Fœ�jM�Z�4F,b���C��ܨj@لy��yj��PJ�ş�j8��G-s�*b{6�6�m/;�{�/��*�I"�T1�e32��j"W�9��u�īM)��?P�J��޵  ���]���<�&Y�꯯&Oh�#dR���NwEi{�X|�(��}�]$��mQ,:[�����bR43�/�>a������C�%<\���}ˢ;��_L����0%��i|���G��&�̓iy]&�5�U�xAwy��S�>bP�q�ɖ�i���bcH(t�~�3��`4N3��W���_Pq�ڸz$1���%m��a�k��]�25�e���z��Q���umWŶm�Êm۶:NǶ�a;�ضm����Η}���_�����c�k�k]�7c�̑ݰ��ݷ�ʗ�������Wwx���	/�a���+@m�a�>Pʵ[j��������:��~>���򽉘� ����G���@�Bg`��p����A|��b�a��E�J��s�� 3�B+>�0>�� �,�n�=ۭ<��Т���VHPz�B�����y��Üi�À�A��9��aO9Uɱ�d����N�d��dOo1�E�YiH�Ť'EI�U��� mR�ƅ��M�����V���j�Φ�R�Ő�����ۥ�u;�((���������i7��I�NW�/Q܁}��J�FC0S)��J��#b߻����;��U����x��V�XdŒtm"cb�P�w+œ,&C,1����`���pV�
q�6��mr� �8��^`}��y����ܜ��oԲ���}��]�j��Ь������3S�MAk��`��dY��n2��O`��w7s���,Q>s��D<����VctXI��oȕ+��`
��@�����ɫ��2�Xf"�����\8�/|�H=�����+۬��s�c��^>-�Y��&i�����3U��8��}�h/��J�?e��M_7_�z�@GG?_-��7�:m����l����p E�e��3���r����6Z��!2�G`�i/P��z����?�%D�5�O{D�(�� �����IX-�ԓ%�'�,�O�C!��_��]K��\`���!��y�Ō�n���-,h���B��FUd@p,��"\�u-k���������=P���	���an�d��������H����d:G�����������=��vi!��4�����^����p߼2�f�K�Jb�J�v_U�����aIP�?
����::��W�����<4	�����"j(_����U!�@2^�d�����]RLk ���i��P�w}�)���9�x�:U�>m����Pz��D��3+���0�����"!�;%e�Ib�@��y�2��K��tOW��I�Z2o��DI��B���]��Z�a�:�a7��a���y�;	��n�`��!����k1ssh�_tex]���>���9==mx�h�E���m�<�O��^�?��lF���=#�8S����a[4�a�s�T���;�{�b���͎��_���� K�J4@B�@<:5��G��K��#&�s�����wVh�/"�gl����o<i��rL95
@[0R�H��8�	�v���Q��Ixs2����:|�ج�Q㩌�����Dp/$]3rpI$I����?P��98���:��4������C�A�NON��`�@��6ғ����欭�ك�����Л�@����%���d����n��U��Ϸj��PAZ�w!�Q$)&��N�&@Iz �S�Z2�z����*���u���犱�lZBR�K"aHB�k�B3�+WWHH��[�9m��1t�Q��j ���&T����e���(.���_��������76dP�{X�[��^�}/���C��F/ˢ>���v'4Tz���/}�����g�aA�K3-6c�=�j�-4	`�ט��Y��Ƚ/�WH���HG�H��Wт�ğ}M�K�;��"!@������D��R��y��q!�}ZP*54(�C(�o	A$���>6氲*�sd&
�%�t��U5'^Ġ'�q�g>�R��./e���q�W�����@(B��T�Tv��'D�w20�0j�T�y�p�/�#��dq��LO�Aq\t�^ϟnf�[)-�k�H��_��,��<h�BМc��ї6��\�s-4#10��:�V�HAWv�A��b��r`�Y�B3�{.�9�øz<�%��� ��L��M��®x������q#S�u;ո>�Ə���*�ܮ��<�'�D����C�Fez��
�%j����}'O$x^�L�4�=P/��|���¿}%�*%-m}�]����GM4!�6drF�ʩ�@�\Ǜ�����C�gTo�dxw�˙^'��"��گ5�"�s�����CGZ�(�~	���:�*X@�Jb��@⛇�
sj�I�������Αe�sx0� ��(���������z�6��pF̮� \��a�u�����β9;!�\6�H���(�饀�TV���&��RL��d�y�p�*�Ȋꮌ��O����у��"�v7�(|��,� ��h�������.>�!i��V�Ek������W�݋������$�~1-�
��:7��Ō �>ݾ�������|�i���X��O��	`�K��=!�����ɜ6�����jr��VN;<N������/N�Hh"E���F��a�Z�"6�;����&hIg aᄰw��nURY>T#��H[V��/*N�����%��ȴ�1W8ް���hS�0�n�W����F/�l|6�+���e�����6��]W���Ӥ=y3
��3��O�-]i��?�LH �iC�(���%���trF��t�ʉ��4��ᆌ��D����|�	~$�!�geb���wY����dn��e9S���:����ƌ'G��)�l�LU�ͅ
������xi�Y̸�H~L���Џ���6��b��YfR[,A^��&��A�
C NՋ3��b��q5�8���ZsO���z5���I�9	3��ʕ�R�>���֞�ͦ��C��Ś3�X���UIp�1��Ǥ��q���=_�$i��R�:��)���(���I(:�WR,>ZjO�g�:�n��P�P�z��)�v��ؔ%:'.�bi{H1p�c�������>��/�;�?�C�f��oq��kw��>Ul�ypp�x�LH2��%X�x'�">2�Lx�z�B����7�g�e\�vt�Y���#�j?)M|H*M��&A�l0!�t���w�D�y�r�J�������'��RŶxX�5f� i���#t�n�B!��
*�(]*Q�g�	�^��1t3'���h���Pɳ��)�K콈+/}��P{�l>��swI2�~�VbV�� ���q�2�3����H�i�#��#o��X���bmQѲ���G�*�r����(�fl{&�]���m��Y�w� ��*�Ė��y6�;$�߫)2����x*�;q1`IT�'�|md��wȟ����	�6�)��	�R�.��B()HiunjM�cS(oD�¦u��0-�У��^<�{����/�"��UH����|!6�-ꘗG�a���o��z_�����'hF��6u���cE��m�\
���k��ll�ww�s<v~��P�����"f~�}��`�?f��0?@O�:�=�)Iӧ�phw?h����������I��lY�g��� ��������q�y>����S^���3x��ﴰl�O;9<44%��"��'�I�ŕD�
�.2ң��~aDN{̜�+�bh��S犊�Cģ)�e��8
e��CA�d����B�.Uz����b�2N�6.�x�f�
.�/�xcj�=ҵ�[�F����*���
��p+�@��!�h��2��kF����¶|M�a�)�"���+9��)�z;�����Fz�/�� ��Ƒ��Y�J�n������Й�$��c{o�ʹ�K
HY_��2�K�һ4d0`�U�mQ)����L@�B�7��6�uWc3��\��UpaDJ����5�����`ƍAQo�uU��=藔��B�G�$d�zl�V����� �kN{�!v�Ie,R^{Ҡ-짟�	+XmPȿaN{li�w|=��Q�*�Javh��D�ە���ء��4v��icX<���������s2�IJBŕ`KKs�n�=���N)*,�p^x�B���
_����/0-+N8��B��s���ĐSv ��&U'k ��t4V�YR)%ˁ��.�j��=�)ɭ��M��Ii?�\��!���zb|`�Zɿ0KC,x}���'��� 2�1w+B�AٰY(�C�0Kf2"�u��E&	�S�N�p�x�|�+��H�"���6d��4C
28((?׍3��jFB̒`(����4܇��
�*	$$"�		@ ���aX��hT�|�ڵ0� �An+b!�*�`E�f.$����3�};U�D�15n6�/pيaޭ�29�&�B���;���T��d��9{�>�'�����r����I����m��X���I���mI��1�f���w�l}�y}w���`����S�6��j8+i�'?-��L^�����������rсI�r&&{R���@��>����_�xX��@aj"ңh���@<2B6�'Rǽ��k'��-������B������O���s\F�5��!��5�
�J��-��<H$�ߨ�]�ZLUFIhi����J�5X��;p�&��h�g�w���D�5�n\��=�񝷀�򶵏�N9S�c�dTq�3�H����ځ��o�g��j(�4*J'p*ayS,,�K]����ho�~?_�n'&:K�:�Z-;���u��{*�_�A����	�m89#Aђ{e�s��b�K�d�^k]i]��;����N�:	��X߮^JLՉ����'�	��R���{q��	zI���!�Q������V��
���N��ߖ�hf�Geuuu��p�h�FEz2Ի��֊f �N}ۡ�[��9*B�W�2T��mc4$IJ��*]l۞  ���;(�O͍�.��3��tB�ҥ7�>�l$�A���]�C9B�Q�v b�ڠu��7�ť?�k�%�����
�x���lAZ#��n��F����<xo�_�:`��~��G6��\7��|��s�~�d��qi*��*뜳��s�c��w��<�4/�O� ��7��A���nW;�K��fE��&c�U2y苁Q��H�d��VO���<'Q���nD7�8G��������`�_�����r8��U`
i��C@Y�Ґ�P6}��Ju*a��л�f����8o�)�
�ñ�y��,�<A�c�X�L�d���D9&�4�i��ΐ�
v��M��V���K`�{�H��.��l���g;~!�#`�_�)Cњ���{F��jz���V��Xk�g̊RjQk ��Tdj}������{�V�Z��y�;l���揚Κȡ9��R����$`U[�����~�<��P�!�F3�v����5Y��#s�h,Ivvv��*m�[�W��TDtϼ/�;å�Su��.�'3�+�����d�Z�^��x�I��k�}�����7FǹȒ.�x��]'#��G| �2���g0
sI�ؗb���*���Α�U,�AkIgF��,���ow���Hh������Կ��'(�ܻ�?�]�!���B+e~C�Qt������K%O�E��#�9��\lQh�h>f�CO��[/�:ꢭ���;�a���ir������a+A��V�2�s?�k1��^�����a*�9AO�کO�G�� �(�*��H����}���������l����<�A�*Uk[����4�l:hC�e]yq��ӥG�w��L��^��Ǧ��}l������� ����?������klll��(�-}I_��q�VK���D$7���r����I�����'����a
�x���XJ§n�ZZC�l�=�|�̧=#�v:H�E��  8@0��}&@��E����M�miب8�^�K3���J��\���HEN'��w0�_	���1�I�LN��W�Ww{*���G��&�O0|�pz�dn��+�Z�p �#]�yI��0ɺ\�_�й���tH��� ��]]���cl�Y��d0�sV@�E�{{�jE�|�*�����&�����7�4.�q�2m�I����+�����S�j��{���b?�u���k{��I�)�7ۿaC7��I[�@�@�(���&�x�8���"�k̈�>�sN�[���4�E6��s�H4TH��gA�ɖ�\_	0� =�sP�	���\_��W[�J	���Dg0�Q@�E�L�iǅ�1�U�x�6��u9����B�<�XZ��}�@WZ͐�r���u�A`)�]�h�zEW]~�1���u����i����rU{�-J��k �N |�W��b��$��5�6�A��R���ۢ��/W���~ش	����ˌH,����(#-�3�Y;<)��Z}��˸/���F��M���"�28����m(y�Uhg!�A���!H����~��Z�8]�O�J��0�ǌ���v�JP��B��7�9.��b����̨TR{��-������i�e�o,�o!��$K�_��o#L��S�%� �7����\Wcn=W� cmW/�&��v��`S�9Zn�zV\rSM����//b�8ѮZ������%�.C��ĮJ\ջɴ��o��9�^��V�s��'�� R#�W�NZ[e��L�.���Mxb�7��Qꜷ��܏�p�
�r�/�5����78n�~ &��@���vM���Swt��K�\֬��^�7>�d[kr���D^M]�J��y�~q�(%%��Q#�}��xF� 7M���Y��k�+�/�iր�:q-�ڈ�H*YʍoYJ�<G�"��� \F��r��}-
���洂��@��v82�y[I��Y�!��ROR��Y5���u�98Vǧ�(�KnF�<���,�����Jj鯺*�E ��m�ȵJ���4� �^����(��^��hc�e'��<��N�G���az�V�e����P�B�(�e�"T��P��`�߀Z��K];��1�\�2��1tZZ��2�?M�{Aw��<��_��6�~w���v u����:�X6*j`24�S��ss�?��O���gma�773��4�(.��.U��\S*�s�(��"g���(�[����S��\�F#�����\A�2��|��ZgǍ���*��;I���*9b�|�P**j���f\�c�1��}���2O�$tKv%-��8�E��F\��xI'g�QV`.>!�L��HQ�|gE<H �r�)D��+`�ͽU�j�_WRcQ���nź�
?W��/�&������
���l�]uv�6�ZO�����SQ�wz�D(��@�I��P��0~�2Omq
���k��Kɛ?S���c��X�
#���%��G� �E�����y�t�,^�Q�@�j9���d�U��Ӫ���4o�g�Ĕ���⳪��9u�XLz+{K����mn��'��L^��%аdZ�u"A��H�!�І��#��6rR��(�IO��Ȗ�:%��!�۝�"#z6{N���dK�ZU���I�ŧ>���q���(1U�bܮ�Z-�����J�&�>�FТ��3�/z�n���C�V
�f.�sz�_P}�Is�֧-9����9vo��cR��<_k��S����]yX�h!Ȓ�(n͒H�J���/4��p[�?�Y��0K�e����Z�HVv�0�L�QS*��t�`�2��Oǧ3wo<d���D���.�A���^^ �i���_���*�M�!�$p�=�~v����$��Fx�[mjg����������B;0����{f�)W�F Ifp��X|����^��`�B-���s&��u�ad��:B�$\ˎG |��Tۚ�( m�ԨD[���J���}�h���Ny�[� Rg��.����a��ꮏ��tC
��Ť�̈́��9���,�
喫�}e?o�n G�i��x�^��⽍Ξj����z�i%������D ��'�2���U"h,Έ #d������_��v�)�������p�[����n�ؾ3
 lN� gAN������7��Iޠ�!x={�eS�P[��8**�>%E�������cK�+��n�<� ���&V�� v��=H�d�&'��u�ب�{�2�g��t�s�2��nK�����)���Rw�A�+>~f\�qOd��Ī%��_��kB�#sE��'\�ar 1KR{Uϲ�d5ږ���hTX���2̉�w9i��}�BI��D�%S�?]�Vc��N��7�G
������(�	WH��������ݙ����$����v��㛊���4�lڬ�#{5[Nwe~�M����ڷ-ϒM�eyO��ġ����f���t�x���H�%���������y6�aQU��v+-�#��؈�C���1�'�,B�P�V�͍�]M/���vv1^�D��ʉ��N���b}�[w��舨	����-,'!1� s���i���aŦ4�G�E������������`������ό6�m~i����B~���}y�/߆����܅Q���v����n��X ���m�KQ�C$0�;=��;E�W�����~�K�Y-�Ԅ��Ic7Qʬ~�T�s$]��c?.�����������X�Yeuұ8���U!Ɲ���X'+��z�0=Y�զ6�u���f���`"���kdB�;h{(��/�ۭF�%I ]��!�8��}DKj�*����YC]�>^�<)���({��K	�(�h����������	��N�4M�,�A[��s���9L�� �̈[���qX<���qU���wg���wׁ*��$E�����{��Z^�����,p�O�d�&U�ϟ��8�g	;hn�_��S���VTw}��EE�B�&R�pQ�\ig��WN�J�)���|�&B3(�!̖r��ȸ�]�"��s:����Ee/4�/��ؓsb�+����H1 ̞��䢱Y�>�٤�J>uq�-Y�/�S硑���-G��ۨ��xI��]i��[~�����ޅ����$��ӎqA�5�8{�A�$v�6�f](�j];��M~saɵ��Ġ����]�V?<�Z����+#��d�[Ǻ�
$Ϡ[k��wQ����-��/�իJ:I��]dל�~AU��LzH��j�Μ>�'�<qm?��p�vZ����.��oJ����qD}��C�����5=5>��_o{�YtK1�����鮄cHzKFE��!�#G���.u��Q8���:Au�JW�X�=��t�����\��$S�]��-��������̌����T���Ӵwnf��m f�"�U���������k��<.��.�!"�;{�x~�]A��7R�S�$�oC��TEyD9 �p��<]�BI7����	���d�Y�X�/��Jd�	�{s���"2
�̹�p��!`�`TT4�frڣ)�K3㦨�d.�q#f���9�FPl��U��Z�v��i(EIQz��6a�{]�U��xW���(���/���x5�{y׶��Mt���/�m�$��8G!|�Y:	_Y[�(ڊY�ęV���8%���OJ��L�]��͈B�0v�0ՁM�@��\�
ڝ�boy�"��L���	'n�X
��u��gfT<x�Y=��=ШVLpT:�jJ�*:����7,x����a"�c����idI�-]���ھ#Q���]�����c�jkz�P:Ba���ET��i[h�J�_� ���pW¹�/ �b$R�vkz��ʊ&VWL+�
-
�����ʨ���X6�����_�#�wÉu�S�B��ՙii1���*.W�׿�|��d�%���+z�Z;����?󴀁��e�g�I��!BP�x0��d�:���N��{u��� y�j�K�2�n_��]�Z���>U�o�@�5h�'�B��v��9�r�զ��s7�#�Ďڀc���8p�q!���Ʌ�!� �3�S���qnͪG�󝹜�>��}�$~���X��*�����W�����_=�R�,��5���x��؋UJ��D�&��]�v����Mt��4ƌ�φ����5IԢ�Gƴ.��h&K��śu�T�l���H$��ث9wZD�	�QB��~��Ѭ7Y������ ��ǀ���ݏO�����ž����~��lA?7]�w#�A�@�����|���i��3Tw89@��d�_,�;P+��ǌ��ӻ���	�d+(aƓ���0wz�~Y��|�q=N�	�'�w9_���s�Do���5x޼u�D�c�7[��r;�XI�l'���ɨ����{f��yD(�.IƼI���d ��뢔������>�wYL�+��J#>]�#+n�8�
5���@��WT|�S�� !�;�B�4�����W.�l|�����~ր3�@�_����A� ��;`$H���b ]�����߇��`���늏"F�����)��k�q�XgS����X�a���� #+[��g�x9s�=���r�����w�
|i�S.����{���� �F�y�Q�頼9��j���K��/Uq�`.��l=F���ɵt��,쎗 �7�׬k��T��3����v��ܼ_�����������*/?���^
�AdHJ1|�y9���*.|�,�H�c��i�G~��N�Ҁ�(�e�Cs8�ݏ��y����`R�Ӂ��Ә/o����+*Nsj	�Aq"N�u
*b�a#�uG2��T��iֲ�f���֚LQ�r�Ր!��%"��$�ĥ*�
+��'w�ҭ��C$aO"
�Н2"����è�ϙ����ZNvp�ԧ�����5�e(k,�����k�TwF<�Zgl�ŧ}��"�k�"��xى���?��������3��B!�	�v�`��>_�&��J�������:A�eف�Uŀ��j�J	���F�I�G?c�a��6�����n����-�H����-���9�J)"�#��YFsԹd����B�EY�``����~���Gz\6�'aU�ðMep����}{��d��&�u΁�,��f�h
�D��
^���&�s��&{��6Ҍx�k��Par�� �J�+�"��&�Q�S����rBZ�(��S	e��J�]2�\}�;		̈R�JO�,]� ��!��J���2�Y�S��&��@�'VT}�nR��)��H�tܸ��aC���!����	i��5�w{ƆyP����n�<S$�I��C������w.���`}dΎ���ktŭ��E��2�Q���i�j�8�z���t�T63e�����g�;Λ��m��?�ҭJ���Z�[�ah�Ǖ����5�Ai�qXP��*��#�|i6�z�BǴ�"�
<�qm�ԯ�uO^4���.9�n��ޞ� CD�F����Շ�B<@���2/M���|�=ҍu�7aS�-�3��l���ކ7B"�'*������C����e�+SG��5�nL���Ku`>f^Ɛ�9 �.m�9����Ɓ�q�'�P�_�<�<@��
�=>((w�}�����|TS��d��ŝb�u����̬e4�L[p4�jV>}t�io�ʒ�𭌊J�AY'�(��ҳFXG��b��z�)%�Y��J��X�w��e�q�ʰz �ĭ��|�ˢI��g�]�ϟp�[��_X��/NR\x�Q+RM�O�8z��U��Yk�JJH��jL�,�#��qݶ���ކg�D,+������7��L��GlC����L�P�<$`Nw��r#�� 8�Z�Wj�/┃��pcB��B4���� ���$\'�
�9�D(��()��5�w�_�Q��wr�a� d8��pGV�Ě����V�%���&�Z@�����U ���L &-���	���F!/�3�@���\6y �jl����+t��P;���[��?��?��,�c.=
�2����n�@�$��&�ݾu^�������$�\@l�<~Q����Cʜ���J��DPLbu֨�S�:�� r�k[�P����Y�8 ʕW�������ɉ�������b��࠽���{952�2���FY�B\DY�>��8�]���wy�h*��M��W�Ca�̆����������/�k�:ݯ����?���V����5��\82f��"����#���Z�~)H2Y��LIeOZ&@���E���'&#�SFK��+<h��Nd�O�>(b����"	���<�rBR�ӱ�1��P�>�I��$F���#*9g6�414w|-��s�P<c3�n'j9��l��r~�#��H�0�EQ2+TԀ�m�/(�Z5��m|���|<��	��-�>v̪��EIK��l��k������t��ZN��� ��
0�MD�����|a�2T�D S1���!�@x�H�e2��&���R��X�o����ç���<�S΢B�����w��e)�f� �B��zG�]��ίyy~����m��O7ۿ�pɛu>ny�oy_Dc�z����Gz wo_�t�&���@�����Ci��;j����|a�p���J9����J2�8 P���ykd�N <� �6�DT�k���bج(OZ�,{xdT!C��e���Aw^��]�i��3Pa<��|H[oaN���	�����<�T��Y��PS[��EG�7�[~G��!"��*}Y�����=���8����Ӡ�	pE�����1(�v���f�.�m���FUu�ي%j_R�2H�����lW5E+�{�Li�"�Z7��g�P�"6/�CA�,>�� �E�_�<L��>��}q�A[��:N_�q\eĲ2_W	'�c�lىqj�1��"�\�e�58N�j1F��L�O�?���7�⎭�}�n@<�~D���ǴL�P2_qB$�
�`�|���a'���L�`�(˪iPNn"#%��A��Dw��*�ܨ�� @��*S�n� d�/�����S���~���+\� �/�y��y����$H�H����!�>��=� y�D<j:��ｺc�=g�B�ţ k�$���l��b�|�@��P������@��1Hk������a@IX_Qs�����k��x�7;�ҷu0���lh�я��ڿ��;Rl��J;�΄jM��"7�5�2��L&�����2N5���K�+�Q}۠v9d��T���II��L@��[�`�E�����o�����������ҞV,��V/R���F����
C�k&<\N�U�����~�Ǐg�1�K��8m��)�5|Z��XW�����4�cX- �)-C|N5�#?�_>�
c�ĝt6��1ë�)~����B�tf �7����W��OX��V�輼~���J�NP��=.�0x.���Y
�	�)����.�;6`�-�4���*M�����&�Q9R!|ܞ[��$N6��b0TC\��8� Y�O�4��`,���-j���-X�E�p��c7%7�Y���NY���<��������Q�����k���|��6��C��S�{�r��W��8=���	p��4{����L�$�R*���B@595%�jg{����,0��V�Ӆ�O=�	�@���1��P�R]�5T
x��@�{*��b(�<qd��y�������EH���u|���Ů�'�ˑ� 2ю�QI7�r�*y���;�� 8��f�"�����#Q����"��=�����ޏ���L��O��xxk�8����A�p�9�op�se�b� ���n)����t:z�n�l\"y �XN���<� <��nr�Ӕv	��Y��w��E��e����f�j{y���{��0[)�'v�%{ޗ���%��q(����vU�IL}o'��6ۊ���H��M����;40��?�U�Ŷ�0��:�B�ЄRtT��kl��|�v�e�B�00)�)����)��bb��7�`Fp�+�	�c.M��*�	�f���~K��-o7��oM���#Y��,�I���M�nfY� 	�D���M����Zy'��5;�vJʩ�	;�Mr�2e�	2㦺�����<�n�U�C��r0��Gb�b��1ųZ�U��<��;�e���B*�&a��Q�v��f�u��&G�����E�p��,��S���_�#j�^����e!�>��U�9_bL_~��Z�jF����ӡ���Oтf��Oc$nw��VKSڋ�:I��"]y�u�$�o7���lW��yJ�;3�G��n�zx/;�/R3�kdӘ$������U���(�S�[���h�T�Tz��٘,hv�����$���X �~ �c��|�e���x��j��!�!B��e^!B�_2pTLo�{�'���!����������w�����q��`ݭ���k���׉��[-��4)��H�������J��Z��5]��Ҫz��#�]	Ԟ !Z*eDX�.�6t���)	9�j�s� ��Úɒ��}#�8Zet1Yv��{�_z��8+JB��'�}���t4�N�7�?����>i�Q�d�$}a�D]��e�'�G�Ig��[�������(���ǎZ��t�r�X=^l�}@�~���Ӳ���ɟ?x@�3��n�W4�J�_'\
�O[��\�Ո�~[�_���� �x5'����*Y��#?2�
j��2LOb-+�^�~�Bz��D�mMvm���G5h�y8���1�
�b"=1i|JQtG��3�v�"Bz�����|3-�*�K =U�?,iC�-nZ;r���qQ��w�	A�0�q?�=�b�CC@�=b���G ~��� ��h�S!�uˑ�Q�OȸlOp畴锁2��3����a!�5 �\���ġ-g.w�T��X�0�DJ�Fw�k@��J�`���`"�+z>9��� ?T�� k$on�܍�g���t� ��^|�2�z4\S'�H�-�����ҁ,jk���>������yz���$�CF�����6��'�t�S~����0�	� *+դr��y�ۮ�f%�}KKk�H�%�j���٢�^�������L��:�q����肯�m��$Vr��f�rpdHG-��_sV��jwfwTn(;%���� #�P#xHm2Mw���d�y��v�,��w��F�)SC�{�+�%���MMX*;���/��4��^?ݵ�?t�͠��v�F�(��b��[�^:tb⯀����X+����~&)���3���sq���}����w�#����RO��q���h���W���W$��e0� J �1��#��X{cr0�Uõ�����J��&��
6B�@���4&;��ݯ5�<��&:��7IywFz+�Kw�
"j%ns=���GVxo����g�~��m�e�&V�Rj'b)Z���d�4c�8LFn���}C�e������+�?�0̬�p���ʅ�V����֦,�Rr��!��?���g34�	6c @�lh�סi�Y�|SR!#��R.Xݫ�F���GJ�dsޏ�|6����ý������9	�?�γ�
���A�%�tttT���R��Ș��S�A��b����t��U7��X�!����0γi֖Յ���?�ONwц�G |F���R�ޮ�_	۪' ��V��z�V�*��N~�$:]Vڢ��k��(������[�����A둈'��ݑ  1@���`'�E��C�;-� ��q!FA�8q�f����￯q?�<o��8���4�8�&F���Zu��WI�p��[�j�C!�\7�:��~��2�7�"���b�7`X�}{�����]2YP�=  xߎe�/)�,R$�%����f�b�mN��J��uiP��dYSc��U�/�}0PtP��B!���'�82�̟��
���t�/.�&!G����|��(u�Nc��ޠ,RT��>���x���`�#4��v��M
d�F���3�]�24$,^�3�nmees�J��X\�>F��J�sc$�I�[%2�q����㙼솶a� �_�w1�R��dkݙ�gb�6M�^cV�����4��f�*dhz����Sd�\绂�g��0i��W���?`�v������D*|���W��*�15�<'���B_Y�bǻNb�K�#��+�NLU�*�&�r>��|����ُ�+���zF�s�T}}ߋ�y��H�������\��M>s��� ��\�iRF`��E%\OM)}���m�~7_eϱ��
�����_��� ~;��2=��n��x
�0�ġ1?7�7is��s��F08(�m[�&�x��KB��%����b�T����G�W͠�b����d?��pЄ?��C�w��哺4��^�{��]�0���Eb{�V]���o���ib�E� vX�G�"M�/�ռL"9z$�.���=�;�n
,?IXL�:>2�e���p;��^��6 ���<|��C����hj��y�!�d���.�0�L���U	����ψ�"Y���333�d�_��.�%�|��p�{�oɻ��p����8�ˑ�����@�tv���*>�E*�=4W"��0߈NH��B��BԼ�9�#�3&E[F\H��S��M囁�ق�"o �㚹!Rg�GR>�Fz�q���	��}��k�o�V���M�D7�%l�i
�������ƪG�h�M�"�����"���t"��9tT2�t���w������/���J8��L}ePM���{p�`�����9�!������݂���=�sy������[5�=���L�*�87C�rR�s���IDb�\,iY��J�&�9���ŋ���+�Q/��y=UV�'B����^�?�e'�?3���q�n������C�jjXQk�����%q��d���Inv�۟�=m;>ֻ��u?�}�ny_�e񸾀uȧ�K�d�O�/UjV���ג��/՝�q�U�B��gi������-�ms�����
-��� �՟\�W]��# Bb�
�����y�u9��hY���Qj��j��2�p�H7�h �ܽ,׭�fu;���Y�̔�'C�J|�����`K{ޟ.�1�jx�\��0b����K�]��2�?����Tm	t���v�/Fl�O�w���ސ�)���A\[��n�&*�6<ޜ����*�8�Ñ��&���(Jaٜ���f�~�L=�W���Q5�+�4�b���!>*�˓WpV�DU@���8�QA���Bi�#�����YA}2�^2::K�A�X�8s-��H��|��y(���rO��a����~���cr���\�y�������x� �_ �C]Ex\�������"�,4��D�_q\�<�A"�z�����w�K��M�SH/���^�ρ���` {�qXb5�Q�VD������#V�*��5K�:�Lrj�|���Y�P�)�3�8RdN�r�/���-O�kc���c��OFcZE��O0�m�;!%��L����5.����;�Gko�=ޱ�J<A9�B%!�iVw^�^�b���l�֫E|�Y�$/y�/�+j'�9xQ�!��W�(�Gs�[�)YgN��[]U�É�d* fD��5[�.��I]:~�f�=��A��Dbl������lWSG���@��ȫo-rB�>�`��]@7�'������o'�L"f��`"���#�x�㦂�uLR�l�!�0T �����~����R��/
.X%��6�Y��7���0֛�W�=R?�K��W�Q�Ĝ��j���K��#��PCB�iK�7��u��J�S��<�%�d�7;;_���BC�)�C\��%��8��rr�4ʔ7{y5z���a0�Z�q��{E;��}��C�$v���{����1���#���{������:�r�E0�"̏^1䏰�A���1�GF�"yˆf����![��>�i��Y�ƥ��c
��Tj5T�'��:��2qq�=W���`&a,�W�"������ā���[����U��U�?�@'3y]��/�4/]�μ��M�]]a �*P(�iw$O��u�DZk�^t��y����~]�C�j>�?�\=>�b����oE��;c�7B��������g���AH��Ǘ����Le*���b�������w���Ï9��ΣlO"ǎN�Z�?��;��І;�TJCL�?���c���+
e_Hm�B*e���y� ��w�Le0 _����GR`�x�Pcs�`}:��U1�|�a)G�`���,���,(��9�c��Y�O'��-��Ԉ���!��(�.��)I��=�uS
Wl.��xx���Ef��UT�ᆻ��	|�]T��@���S����B��/7-'�֊m?����aYZE^]hZY��ͩ�j��h+ދ���ם>���,s����%�)�d�r��:C�DI��,���)���愆�:�x��.o;,Wq|\�P$����xn���dL�����2�{K��J�}�v�n��^��/��<���>&0S�����'��y�����W����Y���9!�U2m�\MS�j���|k��%2�>＊ �Tf8��C��UJ��?"U�2T�ϕ�W9y�S�4��`7���L�a�$�f���l>f�����
\�l�(�G�G�_X iqk���+ɱ��DD��K���l��"���=��-W�?{k^�8�DT׋9)d��Ɩ���O�Dd6�thT�0ӛ��tg�y2�Q�סbW�ry �f�z�0.Hc1�Sw�U55�@|�����Kw�xRK���L0[I��켔K��@�R�@e\� LJ_����&�J[{�9�+��.#�����צO��0dL�������r��"����Oߺӥ�E����Z��-'N�o+���ޡ�V�\�.���V�+�?�^5�}Vy�B��ۓ��nX��f�B��q9���ج�32g��|���[/�J�unn�p$:kp�� @�d�N�.�"����k���C��LC�� r�:f�Y(J��n&���d��ʩ��=��D_-Խ��	��h�j��:Ć�H �'˯� �$$����_��gG���I��A2t<�Ѹ�+j�~hNj��ġ\屘�N��<5rQ��&+�8�F�B�v2'i���b���R����ل�"���6�B�t:�a�^��T�	`�(� b�2C�g�Ht�[e����I��u0�:< �4=-��2Ī$1�zy6.9�����(����F�2��d���
?�M v��h�IrJ�/��M2��J̾1S�gr^$(�� �c!2I�`Hpo�+7����s�Z�^'��֏X��P���R�xO
��,k������x���)��er>�8�ڜ����rl�p�s?=?O���z5��e�h�4Ň�7U쩬RVxÞYuA
��g䨊8>ee�;F@�PZ�8�q��"��A!7�Դ����J��s��#��$Dɟ��9U||�8�)��@(�R}h�$��x�S콝����#�2]_ҳi��j�b���X�)�
�����JN��0�ʄ��$'���
ؼ̟�ZNkRn rh�3���j�Q(_���ʋˎ*=��9{�$�|���d8u���:n�s��&555S_� f�(e&(=�M����h51n�C�B�LV�q�q)��X���]�`��{���n�B
�TF��|1腥�D
�I��*������{D���*����������|���*���!,��/���0��L�JI9��U���q����½�����9���r���㺥�r�kB�7Y�}t+�^"��?��A<�ҁ��զ z��F�0�����$5�s�D�������^����֯o��!�0����"o#��a]A^&�.I�-��h��ZT����ɛK^6|�L�?�[����5��� ��G��*�I�<ʲ\������o���~��ݥ}^�$Y��U�|�!E�C�O�;�����7��|a�(c�`��ݝӭm��8��Jh�j?��n�%"�g�󭖫ö�<)�,-é!�����Z	�Ƴ��)�Qx�����J�w�$�}�B	�8�e'�ښ�]X����lE�(�Z���v����O���U�f�L�����,�O{y�X�B0N�Ó��?v�8�b�>췻\����9�	�%6��@L�/O���~��SQS#�v�����l���T	Z��� E��I��������f"y׾����u�B��ꋔ�S��r|�'�x]���|�����k�t롷yj<��_"��
���y���c��%)vLZ5�^=��@�|�R�`�\)_��CO�;Vq,�l�Y2���`4�<�z9���ɴ�Sm��0)\d�d��G�E�>]�6�PYd~�W!"K �Z*�V5�������(\,��8�^��Sr�X��>�U����	��AaSC���nL��Cˋ'Snê�
_ִכqt��4,쫩���-T[l��ƒ�l��̙NЧ�{�Z�w{Kp��I���촟ɐ�f⡲�/��*���Dڼ�4���\3Jv8�ʵ�v�����a���jE
���cUyy����p(����$�F_�`�a5��dh��y�zᚲB2�Z���ϳ�f@IҼ��a |�wc�ر�P9���p�F��p5��.ߍ�sVղ6��w�����������Pq��� �[l�/��!z؈M���½:����zo����_�����WO���k�D6��̆n���9��)W��^���T��"�������G(~G2=�? W�w�T�k���1���[���]�|�q�<1c�����F���*ܢ��ۚ�E1ؒr����� ���~��R�Lf��'��',U��閛°��?��e"&��{ PjE���V��ʐ��o4��P)I)� �(T(ґ����ۓ10r��~�ϙ>�'������ThT�F�b�ҵ~�a�;��|�--ۆ%����MAZdgs�%m�8�d�>12n���#�HFb}�s���h�S����|��9�{�vg��/q�3�ž��[���~�.Ot�&��C &�OT�����
�������-�~������Ƿ�q��j[�-��qp@��w��R��u+2��}�?o����n3L�kL|G�xQ�
I�`9�����Le����t�N�O�,��NXd���&�����<;�q\5@6���t���� �b0ğm���Ǔ�v[�"N]r��H�O\X ��w{Q�8������=>��C+ �B�;��.���R�m��Be\˗ st�CI(�s�w/~�p���<��0�R���8��&MS�pT߀}8*c��VG˴��3y�� �u�^�q����;	n�l��h�ܼ�!���o:�W�_����KS;yED���_��'t�����1j@�D�j�S8k�gi�W}8�=ݸ�Qِy���׺u\�H4:;��\T�iQ�ﭮ��_(��z���,�7�k~Z���m�I��t�_af��Y��Hm�w�b��o���ܓ��W���~3���e�N(S�����|����g"��g�f("E����Wrb\���j�3�i���� 2~!}�/���H�<=���=1}�MM��!�D��p���5&���ɈC=~F�3�X˯M���e/�/�_I�Q�R&ډ+�$�}0�ϊ�BaY��<'!{fߐ��+�_���C
4f��5�5wCX5��T2��Ƙ�_(�T�cyU�#��sƈ�9���͢i�����O�AEb��*�7��G
M���:�K���>�g׊�)�pR�jW{:���'^9�fS���c]��5���OE�$JW�z&p��0���uD�u�7�������C����ǎ����0��U�~��ؐ���u��#�x�2���ؼ��=Ϗ����V`UY��*U�@�4�M��FS(����C%�0A�N��[\���-��*���&7�L��O�f%�3��o���M#?{!&���77;��#�σ,�7S�K<j�ƃ[��N�+|��Wj�7��,C�� �ï���gvsNE!\Mg���A��BE5���Hn��,��{>�Ւk�Z꿝H�K(��+�O s@����U�
	F�1�6��A����?67������k��.�*�a<[���������h�Q�AAe�	��]��ZJ��,ߏ��NK�3��}ˌY���7�㖰������%��lT�)��***�/a)	˛E>P��e1\N4��˘�clF���� ��y�����o���(�9U���B���dY� �1.�?^���o�.M�2,���.잝�7М2�0��:���?,a;[����pR���l�i���nc6��7a#������t�9����Q�����v��}�h�C��f%ߢӍ������h��<K���(�"4|���5�[~�Be{݌}L|��455�j�h@@ 9p8��_����6W�P�FK���oyU��N�H>�ᐈAv�L��U��ro�e�J��\uF�v������"_�\Aw���E��Ze-E�hNc,Px����."���H���6c(������#��?Eha-|+,����' ��5�Qh9/6 Z�"��Pw�C�-<�����S ~*�4�d��0���bt.�a��sÓ�����6=�ou'�a�U�7�5�-aX��T�s��� Hd]6����b������j����3���y;���|A�O�6�h�DrU,��"����׽`*�c�6%��M�*P���!��݄�Z����I q�Oɼ��n�a����[Z�0�����d��X�,����l����$vPW��A���2W�xpc�:��������J_ �]���V�����m��w<�{���Z=�[-�w �=4Lq[M=����<��gHf`Xo5y��iF����c��uQ�zu��A8R{�22N�	��cfV�""Ϝ7}������C?LjD���?k<�q�d"��{��=��W93j6��<�a��HEy��K�=:�WN��F��H5��~�����<j�H>���;O�dY/�/��_�:�Eߙ�Ԍ)%ev�$Y9���{�t�Y�`s���a`T������~ȸ�L&-��j#zTO�]N�_-�ɤ�i���ϿS�f�Hx�+�CCbպ>��mF�_)//_2?_oJ#5m�]J
~�G�_jl��>\8^4���͏�yI�P0ɇ�py�P6o����aɉO�~xb�����.<!��e�:���9gK�#ʴc�h;�����K����wc�J�"�!��wi�ˇ�����2�س����`x��&Â������,0r���+����c��Jd�����������mdp̷�]����{��y׶�T���o:b�ْw���ߌ���Y�����E�tQ��8Rp����ec]5��ڐ�X�.�T�uKrf��pHj��ã�ɰ�!�N25�,l�����p����ȿw��^4�ځ{�っ�;���(	mT
���tU�[o���k�G���8�L(�)G��A���e��W�]n���r�ݗ����\��X5���m�,JF�䴏nL���HGh=�;2զu��:��f�X��eϕ��75�	0�S=��}HJ��k��gjj�$�B�E��0c��՟gεv�� ��m&y������� 95����q/�E�9T��L�lB�4�	k2�/���\�|���n�7��<�K�����+�ɚ�M��=������ik�����~��v�k�����:Ǧ�m����������.)qR����T����m/�S"���~���_����ښV=7/�o~ff����.d�(f���r��07i�"k�?�k�`jvy4]=�_u�@��F�PF���~C$�OF{8�ƒ,:�[��-�Z��B�Wp@�^Z[79 �b��ۻ��].��D�SJ���BvSj}�	���d�{�^D�q��+�(䱏r�+�����[W�$~�V���+����r�Mca(q ��vL�U�p�oTU�a'��󒴈�"^��L^�.�լ�	�6���̕�{V�g��-�J���X�K��r�4$��~�*�¼'�b�hM��O08E� ��~������α+y��F�P�  ;B�PفQ���.�� �9`���1�2R�9�1G�cs�������T���uu݆GS��?���w�*�$�ݦ?��h�p$��������x!L�g;��:l ���	����Ҧ��>�����	�`��'ׂ%,�\v\���L�,��e�l��j�t�`�����.��J��j�{m9_\�w��v��/H�@��[L��2��2>�qqqɛ>�������ia�D`�0�4h�^܁��n6���J�F�(9��8�����R2�!Y��e���μ��G��sZd���EQQ�������@�_".��S"��#k����^t^�����W<<<�=����ݖ�����>=���0A�����z�)]��P�b� ��,�����~����T�-2M���ӟ�ӵi�����8ts�$EX��&Y���ssr.{A�a�;&�y*�¤o	
�G�X�QQ��>���;�(]���c�7Y���<1�W�H�5#�@J��>o۸q���2�>~����4���倌|nhd�[�貚��fR �qq��"JDˑkǪ��B���f�8A ��Ph7F@�� }�(9���A��b�xw������ v|>�f�[X���9U15r�Y�� <�z{�� R�w�o#���.�� H���f1En����.���Ѳ��+xѱ%c�W&�4�".��/M�4�ǲ�۬7v��(	?R�u��4u}��>^�[l�ڋ����tw��mu�S��ص�/*a͈<��F|�&��al��7S�Lx�G�#�xw�W���f�o����JW��iqS�N��ml[6�t�k>�?�c̐�n=\�q��E0��� c�xeR�mo�37�7���`t�A�����l��ܖ ��޿t�R�rv�����j�磞�� Z�Pu�ݸ@y�~�m����7�� �$i�N}����&�&��e���Ɛv���&�ev�"e(999���{r666��`EF�(̅�%LvV���;s�?�Y�>H!���+7��ϗ�5��
N������'����)#6mY�<)WĂ��ť�/7Y�9~�? �3�{Ǩ��B�L%�[ �e�<;i<�a���Hy(mi���yޞt'�6A^X3�E�iԻ�;�״$�J=gi�P�9����}iH�����汩����������͙k�f�N)�x_z��q�F�bT�
��T��<��nU�afz�B�}�H�t
�v�~E��HV���~H#��G�K}`EK�Zޱ@����H
�;�^㶚X�s|�I�����z����΅Ldbeǽ��$|�Y�Lo#���+9�89 ى����HF�(CQ�.�r�ә�����:P��� ����wu�y9���8�c�I�"��$��l�L����	�?2�5������H"O�Ct���������N rO��l�O�=����2�����{��9yD�ӅK�Eϲ�^�Ǵ3 �+�݊T�n��_��Z#�!��C�&����>Qf}���~+�L����4��Y0��8���o�)�?pѨ�NSZ��2���q�(Φ*�0u)*6_ae��%��e� �3QTAejo�=u�`��5 o\;��U�ЗLl~L���!��g �VSS�cI�u��~�|����O�X���m ����p��yZ&q�}Fx��~�����5������T�<H?�{>�/̦r>3%���8{̦���ɶ*�l�v���T��5Y�?�u�ƌ�o�̚7������t��i+���L�O���XZZz��՜`"J&ܘV&n8����>	Q$�^�-\����Qi���9ľ�U"d�~J�\@%�ӥ�����p�q�X�T>�x̹EZ�^�k��vrbt��?ӽEY���� �y�K���-W��Y����s��Eٕ0\��;zj\�@\�8[&�F�e�'x���^�i�C`ڳ�, ������Z9.NX}���I�-A-I�%W9�P]�z�ߊ�-z�b��N��sQ-'�y��LLXT�[
 &����!�"��zǬH�*n�ssܩ�q��$��8�y����ݱ���Z�r��bb�KSYM�?0���>���ߓ����FG"-p9j��ö%�2��B��ie8���c�x&����e�(+S��3��V��W�q�R�"�Q�?�i?��s2�b�u+~���t��W�5Es�
���)-+�eN�����-�g�ǯ�(c�5�Eh/9��\�〽�S�Q@��T߂���l�o���z�#;4��*�w�]���n{�-a�I]̶d$C���wcњ4��I"��wN��=YnY3f��]7�-�ׇ��IW��H��EW�c|�&^[K}^ n:��ƅ�-w,=�H_�>�x[^6CF���X��+5Û�U�k*�Wv�b�@.5ZmD<\��d�R��8��s�g���̯��1� �</������	9�vX(�������/���|ۏ�y�f+�G����*��"||vk�?.����˜;�Ql׫7�)s�
�VK�m;?��>ߎ8.e�U��;���b�_F��#Q1�dR~g�>�P&�u�k/`�9�͗(l��yf}���󟞝���w^��N��&�u�R)+�I��� E����:"����M� e����#9�!F*GnM�"c\���)Z6gΊ)�`�+��#�c�Dv�Ȟ�2R�\Ǘ�̒�@L�ǵ�I�@���z�Sv�×@s�a�?.̺��w]�R�5�A�����Aj���5�O|���Nl������p��O�S[�i���Z����!������_i��f����F�#��_<��ݴ2��\���"m�D���Ҡ�^�d�h/vFݾ��٧J}�,��眑�D�9��]`4q���E���Y�☦�J.M`� �T�ӟ/�2Kg~�Ōx���c�'��S����/�E��̈́�	��g2�6����=������iO/S�{h莑���Io��0�)����t�v�MK�Ҿ�~'��E�U̲ܪ�Z�ÌL��M�%$,���'�Z�J)N��2u�ѽ�����:��
�\�l��{]���t�WȻ�F��U�Q�!f�e����>$�2�
�=b>*8�%ꖬ��{ޒ��t�s%�j)��ts�^�A��FX��6�<�7��S��r�,�,����>�����v��ؽ��R�Uo>=��|ZE&��Ϩ`z��m!�����B ��>4���Gp���?��D���S�m�T8KH�������[��rѲ��H㣅D�s,�&��Wԅ��[0b�Eݫ��ժ�Ai>gWW�զ�tXo{
5Z()�j�<�'�O_�y
E}��3���㨨+sh%;@q�t�H���2��e���D �|��<+.���~�b��zp���YeXO��ٰۡ�����%6���b�¶�Ht�|�y}$u��C[�����x~�\n�Q���2�4/(1<<�35�����L��� o�>rZ\^��G
!ˠ�GQ�v��U�r�>�-z��=l�D	�k�y12�I�/]���|0G��OT���!Z��@L� M� g� �;U8O�=*��$_�y�:�%]ć���9�k�K�2r���&�|�8R����d�/&^s�F��y��jK>�� �h�qU����=��a��Va�i��6�*!�QF�8Rv1�c/�7KF�����{�Rz�	-o��ǎ9'��r�Hq5�|kk���J�]�܏��U,�:�&Nf�Z��hŠ#�nn�x���D�]�E�>��,n5H�a��kkG&�kC��PKf�$-n��c��)�rOb���4U�t��#Xt���z�C��J��Q���n�~yAQhF�����3�ψ= G��ci:**"H?,�)�a����G����Y��7�V���$E�Ң&Q�v�*E��y���*z�P��V���q@�r:�������L�F�Sj[�m�>�]�[W�/�v�P�Ľ<Q%$�����a���ڣ���\<�<VD��v-f��#Aq�}����T��^#��-E� �.mﲹ�.0]u�^�Y-U�F �`յE.��`���b�8�o��*M��4���8�=�� ���:Ler�peM��ˌ����`'��rD��|7�"
�ȅ�}��.����1I_���M����(F�^b$����ˈ4O���f�k�M�N�Z0l:a,h���w�����b`��Pl�Q��Y26���U�D��K$˰ ^��8�)���Zs���������?2��w�����Hs�+��?r�_�.\7|N+����n"^}��Sa�#Y��|�'A�m^O���E��"n�:׹sEQ��v;�ǻD��Q��k�7�؂�t�5�k�^	8����w�?[l�1�8ao�(b�+Nr0
������1bhK�v?Z4�)��A�voΩ�,C�goA�fI&*?��A��NKs!��	�䙧�H���3Y���!2�P�LOr֊���Ĳ�"�-9��A������1a�*Rʫ:�~�4�-���8� i,Q�$��/���/�N"�Qse��q;N����?p��.�{�O��*��9e7�_�p��<{uY���U�ܐCUXɋp�B��bUE�*����L��`]�q%��,��n��0���J�X���\}���I!��N���T��Γ��mG-v�$��d���:�lCE�7�P�(�#uu��̯��t�ЇF)ngƿc����C�����FSO�W>%�SŌ�,dǣ�[�i���7�A�g��i'�M�[��=�4��O�e�RB5���Vl<�����y��7T��PJ#x[Q3�~dJ��_0O3d����]?��L�1�(BI�]�kT��]��Jx����Q���C���%:[vk��B��ai��6p�����^9��⁔�s�%��MW�wS��e62 ̾V�5'0Z:}�&W�P3<�0���$��H:�ڄ�of�\�eca���Z���L>�bD�iC���}y8s=�@�����Q&�˻�Q{5V���	�K+*��}�4h�yu�5�J�>�
A���(���tg�K����(�A����gL�54�eL��C�6Z7��z����'f�,8�A�u���F�$㓺���1۾�7Z�o���|;�i�|�H��=��b6�2t;-��U�v���@漽s�~2�w5����f9���r��; �>�e
�������#T��e<G�-�Y��F"�Y$��9�{ݎ'�s'���<�L�GF;�<)ir�PQ�>y�r}�v
���ޗ�Y�E��W�@\�ւ٬���T�4w<\Ҡ�/i)jD��40[�I����5��k׾�*)�$A�1I�2� �-Hqq]�"�3�/����e�A0��_X�k������a�Ģ��76i<)�q�������5�l*�s`T�V��e�ej'�W0��i�l �e��W��ғN�d�ӽG�H�X���+	�4���Λ����T=���c�4�/BY� &c��x�P�:��D�^3�3�A��ppm:�P�B�P(T��4 l!����ו6�
�|����8�6Q�y^�����ru�2�<��%�TXj��^��0�r҃"�]_��� ‷�l�R{L	�<i=U4q9S������'������ݞbݳ�fw�yN��f�wmt\68&mT���u� G�3�<ۥ@�_����J�
|���v�����b�XZ�&�.����g6�۲5�  ����B�|�I�T{fgT�办T61���E��i����1�Պ���������p���9\��&���lb��xrc���b ��r�*��}��l�u1��I�Ȯ���5���?��'b�k�|_��*�_���6��̲^�D����F�F4�u���ہ 2���A����J��Fx-���r��!UB���BF��Ńgcc5���M�4������t-"��ۮ�����{_�9$�ź������a��,��VΝ8o��d:�k�e9\M��l8��<��lj�T{�d B'�� z��z�������'�-p�F�~:��ö�2�F	�5���� �;s���w��C1П��y��V2W�Ư85y���v*@�<��G~*�iC���D�Lu&=�s��ɜ���#�<��J��f@H�����-ϫ���IN���h��ƿ��28�̟a);}�O?�O�0������M���v� �.�_m5[~[�}�,�4kҲ�_݅l(��C��7!s_�*�m]*46��n�w9 <}?��/�[__C��%$�����_^^����x��WV4�E�ENC�\:U����rEs���Yr?��,���co�Ji��"���!e��.�p�\a�ԡ�͌�����6k�<m�=�m��������X���G�I.8�GG��+�B��(BݻS�_��Y��
����&#d��cB�������G�!�˛!d���3��7��^1ګ������qua%m�b�
ހ��0��.���ު���c<���^���zWU�q��O�~�\]l�C�O�G_1{|��N�>v�b�i���q^.���Cf����X
��@�2}֠���H��|�-)w��J��l>�-���3��$f0��󮗡�M�#uw$����Tg���,���M��z21u�X&F��k���.w��Oo��q ��0«�kzP5�ZZx�Q� lmb~J8s�z��`5]r��Q���QI��[�q���˜��ﻮϻ-�<�!���[����}*Ͷ�ɷG�+SL��8��96� DkU�>���O��x^���<���,����x�Y��-"���/Н�1Ƙ4Lf�D�uO%�F�e������/|^/8��!q�??��u�����ܓK��{)x5;�Qg� �ya��|���ַ>E�%�;�A�����p >�����
���+�&,L%e<�l��I��l�!M���0De��p�ѳ�na�(G���Kˈ9�X�Ia��ǥ�ۘ0y�9ї�=�[9�b:*#��<�7���dZ�o:݁#��-�3�\�16�q���TVG�ru����v�Ru�<:t,�����&�W}����7����嫄$9�Rڢ���������{A>0hX%�R&XFlB� H�U��鞜7O\ȟ�����g����j��`Z3��ׄ�0�ǆ�eX/�/4�*"��>� b� w�v&�@��6#6�ܐCv����֜vP���a��[#����+nj(��)���;:�|�ߊ���,�����f(H�P���+>Z���h���\�Ξ��+֥�L�/�v�v�-��Z}���<���xR���r�$|�U}��7�,0,˓7Q��Fw8���.��t�ZiAm���Q��%!p�TY��l'�ڶ��AS�e6x��Qa��2��nrf\�Qz�t��p�ә��lM���Ɵ�+C�s��(���=B�e�z�Hwot_���e��<v��r6h�ԗ�H3G~B���a����f�D�4#&nS p		���l�G���G�e��e���er��嘘�nT���k�Ă�3��j)�He�/�3}�k�����BC� ������χӕ2�};i+@�;��V�"�(�J#R�Õ�χ�[~��}�.����2u]fn���Һ:�b;^n|���_(b*'ش�o6^ٓp��sB��ΣMϕb`c�,����^\��! )`��z9v�n��A.,^qVy�^Ƿ����2t�'NYQV9MU�me�TD��*81�G�,��~��Qg}� s�V��Ia�6G>-R��Z��$�E%Y����(�
:P(�����b~7|W��[��	�L u?]�~s���e����|�hf�}�dG�?�p����Mߓd�<%�WIAj���Nv@qR��O%��������}ā���JKG���y�Bᆺ �a��X�r�/'���]�*�(���!��H4�2��Rc��L_��5�^2O"�tё�~��~�x�������V`�O0@�5�Gv&��^�Z2��(#a!�Is����Z����0٠ �Ag�Պ<	)��Ve��3���n�E��b��2��_�Xl?��K�[����j��Lt\΢[�G�H}�Щ#�ԣ�bK7���
e�!�����p�hD=���J��U�;��¨�XШ ƈ�C4��I���c-2#��f�}�d�?�Y ���i2`���i�Ƭґ249$(�D���/ҍ!2��=?;k�m�/��F�)��?ކɹ&p���y���c��L�pt�v����2����%D�Ss��jCf��JDB^�{"x�cɱ�N����7`x>�������y|�I�q�O�x��6���N��p���&,�+�,w�y�� T`���g��u[e�é�a�)�}�8!���vr��ۙ5M#���g��`��W��p6���I�F/OnyV�����jK���}u}�.�=4�</)�dp�(���Е�y��M0F������V�	�����	B}�0C�uZĺ�C��L��S��|�4J����BM�<���D0�u=�jb����Mj�p�F���f[�%�A ���lP�:mJ�\�J�����l��5�u��N�J՛ſ�d�2 �D�Dv�>����/�Nr��Eǐ��25u~i,m��h��V!�i�cL0S����-�Ae-�����B�~�TXmW��.-zߠ��Y��e(����tu��B�%���w�d��?LZm�* '���U�BٻH��; �v{��f�W�ᨨI؀��E��]��U�>EP�PJqp���=]������@���ռf�1d��d�W�Vp�����b������w��X0�M�i��)H����$���&:�Inp�QFE6)?ȑx=�JK��bO�m�&#7�A���I]��Րn4����xbV-l����~x�;'��7�53~�9���Td�xTޡ9r�Q�#=jew�G�KY?��=RH\+ŋ�)l�TÌV�Y�G�#����zx�Z����^#O�(Jd�]�:;D	[E��LOX���q�L�٬��R���n��f	,䇞?�@��dC͐��m���Ċ�c@�F��b��%C�2J��4"p�R���B��n�6���>�m��~�
&mJF�7��'+��,&��-�����|��ӤQ�#��D@�����?���GV�#n<7�s�`̝;ߞݶ�4�,��G�X��.���^��פ�}�ݗپu���CC����9cڔ�L&�X�V�
�|5�(��yK&	�K���,�pF�(U���j���D��+�L�ZMU�<�J�t<��\�V��J)K�&K�+�3�ؤ��E�\�l-��#w�s�V�=��deT\��mlEqI�1�D��`	���Nd �~�@xa�XH�$r�уx�����kAV�Ae�5\YxZ�,u�	����`��rZ��OzeA뺜׷}[4<0hE_j��T,{���bKx��H�%-��M�V���)�ɖ�����w)'ц�|<�\8�7�ֆD��sow�B�e&A�@���x��P�Ld�qm���(ݕ�s���&�הZ 2��W��*C�9<O�� �u��7X��C�]WJ�>ҵm����m�~�`�1ߕ�(@ӡ���ݭ����''�.���N�3'Ė�L�LL����Pٙ?�Us���N�:��\�"C(���z��b>�NY��]�9¼c��&ܰ~�����x��H�*k�{b��i7�18�����,V��Y�X�\����K����j�y"X����Z�����!�4�&�F̆�R�fUc����ѽ�W�N�ʗ�X��$�'<����P��Z(�3H*�q�Q���7k
�j(?Š(��*��*����i�݈oz��c )Ì�����hc��ڸF+�a����D�u����^���dr{GG��?��O^r�Ǯ��������^{�;�<������g�<n�T��3V�j�2��hi��|;�ܶx��ξ��O���h���\p܏���׬yv��|�����6���@�Z<S25�6?��s?z�QG�vAG[��G>��~��66<83��d[zH��n졶�n5����l���r�9>|ɂ$�bL��B�~�Z�YEV�䈺TݏF�y�/<�EI�Uƕw!�"��,$	)YYL(����6��FB�LX��y,��\���6���|��,��#�������LD�1,�u4N��F�����5Ȑ�6�v�3E<6f@VGa�R�d��#a�8�i�r�����	. T.w���pM1��3tWȒ�У!k$��=�̞mm�����\j,Rzq���X�7 �8ĩ�R6V�$K�����`��A���@�����|� ��n&B �3 �cYna&�ÅVݕ�ݎ ��0T(�ͼC�YU­d�8��x!`'�|��pZ�ڊ�)xI�	�MTj�e
h���q>֢ ���	����缳#|vE�������n�C�'����z�tc�u�z�f(�B=��<,x:+̖��]m@���.���!� ���=Tx$�u�e�a.��%!��9��x�p6��,��wp奶��B��o
���XS�h�>�Ok�]��>�EcY4�d��S	���O����5����M�g�<�kĴ�Έ^�%�����s����-���L ��� s7 )j�q<��{�Ⱦcl��QB���%K�.{��N�{����+��k�o�uǯ�4y���߼���W�~��?p�	�F�2���J{'��y�!����=�d���ϟ��K.���Z�/⋛o�y�W���_�j�U�$���r�a����?n1?�+[�h��]����ne c�ƍ�o��U)Q����5z�_���S\(5|���~k��B�;��B+G �A"��;3Y�R�l�\,y��ŗ~3��o� 1��rC���9O�`P28��� �K��T��I�5�֤ѵ䯗eC�2!m��R� Kq�`�	�������(����L������}���li��"�F�����\$�6�,H�MC�ٙ��/Γ�5�DlX���R �-�bѢ���"������9^�B>T���6�"�M�4�|R�cHǆkL$Hi�	��P�H��{���S�Ł��%}�ϥ�5.���o��3��1;�w;[�aN>߁�Ĳړ�	?���6�
��Ϭ��9�;sO�ya�-o��a���IO5������`eHp!�אE�[L헂�5m`���D�F�v��q����>ge�����w�$��BKdx �6m�ʒ(%�#�pZp��E� zjJ��b������㼲5������Cv,�1��hr�N��i��@�TT.zIm�K�&a!K+ �O�Vp�q�7&e0�(q��$T<CE�_e���c�3ӐE��K�����_F��,��y��1�\W�� ��
r�#wPȨ!c��"���k���Q���U/��۰� �b��Iމ����8��Rd���4���x�g?��O<��뮻n׋/��[�|�w���M�.��q���W7�=|�������lj�!��������/O�֡�>������[o{�E��.z�$�nB��uR:j�h���w���'.�m91��*���kN��o���996<by�=�-Pk ���-h�TI�`(�~L�:�d��k#N�7���U@Ȭ�T"*Sf7��吡�����lW�B!����%��(� ���b�b�3�W�WJ��H{��E׆q���uM&4� �� a�] ��У�e��B���dE��R��J�7@
�B4q�T��^�B
S����B�	�88�>2�y!Y�����v��\���z�٧p�d�)hU�E��8F�Pћ �]<�ߐ���\�&2�D�e��Ȫ�:�:F���bA�.������>=�~>�
�)��w������������ޝ����"�)�5y�$T�%��:F��)3>1(}�3}�P���h��/&��B2��V���Je�Z�$��p2��d��R�X�76�45wtu���c��֖}6nܸ�;�kB�|�9���@M�Z��)��[���a���UsiP4�g�z���G
)B��N�#	�#��ì�a/�$:<Cp^��W�����@��U����k}�[�c�ю���O�K�������NZ�?,��j�����}&bW����O�(sE�nf(Z��\S��@��%X_��u��GfI6غ���Be���c�����'e���Rc!0ó�������y�8�L�c�#15���I`'��dhd���nʔ����|�!�s�:�:���o\��%K���b�(:�~�]�9/�HE����۱�ߞ��U�Z�0/����H��)������?�|����y���9���֭[���3fڳ �q��X�"�{3��|n�U����~���;�s�d���|dp��ӧN��FG�]�ω�8㌨Z.�hQ�hhk�"���J��c��p0��G��w!Ȉ����	�X���&lwC���@F1:����R9��qMȗ�T+���BNQ�N�r��-�NR��и�%VאxPT�Ѯ��MV����mv/ ����L�d��/�1�W����.f��{W��-a��Yh�P�
6�����i`7I�^�	_�Y]i�9��V4������N����h'm�ri
�s�y�/�EV�E�����S�x	 Yi&����o�B��������&��3@0Y�K���� ` �I;wR����	����L�6jLCp�k��SB��c�g�w7��'�ɱl6;�N��Qu�%F��:�J�G�#m-m=M-M���;�7�����ڶ����L�6�0u���S�����&���u�?8����p����?��H�[� 5?,�l�8�D�3��/��Ր�=N կ�=��
`�^��6l��$z�	�&��h��|�c-��!X�AD#��ِ�PB���7 �����S9�X���T)�]0|��q��L���E�+�%@H?(�A���uƩ}��??�0Ͻ���^k�b�u!�y -Z��E��ǲ�b��yi�4�5ZW�-����}�xq���!H�nW����9�#�"��N0/<@�*&[��6�7��Y7��\��K �\�1P��޳�!�p�����|���P��_��������-����T*��a�-1�#�ĀE�y�*<�@�͵\ƞ�\.���'��oy׻����R�/�/|�G\��}���w6s���= 2�1�d)nٲ���c���v[��|�۵��~'�x�9�����qx{ks��d���fG�s�����x4Za,油&���c5�M���rD�P��g�%�Pڗ�u� 4���� 80�Dі�=ѻ�uN4R��-�	�Q���)Ċ[�ࠈ� �Z#����곔��-�d��g1��,<~�~�%��X1�e
.]������B��k�$s��0Z���+ȷ���uV��j���Z R�*�%�2��|����o�����ch!K�	 H��8���8�1Ƅ6mڰq�"a!a%�$�����ٙ��w$R�R�j�x�E�\ C²6��쇝)�}����\�!l�ͫ���-��_ֿ��u��n*���es뒩�p5J��t!ߘI%��[��NY��Ҳ~֬�[[�����;�M�]�F����lv|ٲe�__��K���;�w��M�J�s3�>�E�m����y��;�v9 c�y�@nn��ƙ9�y���6?�CL�Q�Io�v��nI����,�&��a������Ĕ >Xg(�[)S�g�G#����"C���}�o�h�G����n���a�/��ӸRqXkDl"�B� ���'AaE+�řOg�m�����/�Ř�R�.1��O#9"&�1H�|�/��������C��4�3�����s�_,�g_l����.ne��\-�;{���l�?c���L�Ĉ�;���N��l�:88������ꫯ�P'���O~�ӧ<����388x�����g�q<6n�زbn�p�(�U��gm�_�1ܷ���G�����w<��Z�O����~p������%�n����F��gk�>sw�=v�o��N;�Z��j�Qg����.�s�%�4�s�3�Yg�=ںus\ˠ�)��V��	6�E�B(7DH���N�s��U(ᄬ�c ���ڳ-����s�Ic2x�J��"�>>�+	4橇���a��\���ڧ���P&m�#K�I �B�?��p_,,����en����a��H
]@ŭ\
@U��|br�P=������!��W���[1R��������S�F2��ey��P���YN6z��>�w�ж`c��YIh�.;jF	τ�?�{ɋZԶ�+���P��Ki��?T����5^Ȃ�ٵ��vv���A�kxl���h��]��wn��ᜐ�Pf�=s���\����~��W-[�,�{�B���?��[o�s��?=��[o?������y����`�c#=v�g
��ոHTM�0g�JU��Rr��K0��uμ9$8�x�M�6���}��^-�+���g]�M׫e���E�r�X���ce�Ŝ�f�߸ق�P�blĸ��(b�X�%C�1������h�1�M�-�=#���Ͻֈ�1�������ݙ3��JY&xQ�2dh=��X,14�:̽�2/p(���%WS���s+�ƻb�(�%���&�8�L*i�BL�2ڸ'�lt}�2[�bf��tbUgGǯ���|������iE��䷾u��o��?�C�(�!`����a*6���EB?)A��Pjm����)S��|�Iǟ��'o�}W�'>�W��.ٸq�b����-&�����r��c�� c���u`�҃O���?}�iC������~�=�������Jw'�1-&4384���"�̊�SXt|kKK-V���"�S{��FΕ�E�{[Zf���J�mں�����ef�����!IE���J�a%ES��z����S��W�YRR&�cT�E-j�gb`ZZ[�ѱa˾�oVV�'�C%����ajK���(Y�b:�w��|��W����6�AV�O\�Q|�����r�$� �EA�z�c:���D2G���	t,����S:m���L�5����,�R)���q^��z(�U#,;�+E���2ꯝ)�X�X�2j@1�]-je�c��Q;B�*}g�\xq�" Kܓ��P�J�)���	��ٌ ����/s����cMQ~�� ���X��2�H>���~T7��    IDAT���;p�ś�ϟ�{��N(�B�������^{�>����7=�fݡ�ju~�u� ��ܲ��^�F8��E_��:|����,U���uW�8��`�z`�h������݇#X�._X/nI0<ս&���6�'��6�jw��e�	���R�'cŘA���Ɇ�����1�X�q����]b@8+�?�|k��F4j�ش5:��4�jU��x��}-����-�f���Z_<2�~S�)ǋ��M\�@S�*P-�##��	׳J�3�qf�y�jq�����XW���0r�M ����VĆ��\�2Ɗ��-�{�����ξ��3N�����_��߽��GYuj�PX����b����XX�m޲(GFH�wYO��c��`�ZrWw�ڮ��O|�[�|������ξ(��yo[�f��6m�2��3��G@,k�祢'�=r����i�ϻ�ҋ?�|��+Wf�>�{J��~,�J�͝5�6]����ˣg֭5?%�rd�7�I�2vtU�^Ԉ�(q��y����*�%*�=��
�sgy�J�9&�� 7��x�Z�9��+�|#���	^���Cj�a����*)���:����Z��oRR���`[޷p�Q�j�,T-�
���H~��	J>{0�oP��Q฿��9D�Q����P���-:(^v��L?�[�V7 �V��k�"�%%� �l���0���R����
��sE	;�IG�x\C+Fּ[;N�K�j����w��{�+Yz��e݄�t�#C�'0�6L5b��_���l>$|<��t4�X+fѧ��+��;��Dq�_=����ƦMЈ��^��D"�֖ۢj��E��db�T(���^+����[^��~� �;Ｓ��˯��_��3564O����▵���<�˜3�;Qŀ`�x�`%���ZV�T�j*UVc�]�uF�Է~�Z[l<��&��c#`G�tx�׶�-c�����%�[[��ł(�kr�Q���`.<.Ak2���=ϥy�ZP�&
��U,$�d
�T,��6�����'W2,���ܔ" �~���������k�F*ώ�el��[�Of-a�M�� .�Cj��˳S`� \�.�l�1|'v
y&i�0r�>2R��r����s?�O�~�𥉉���K�����L������7��0�5*��L���G�k�f#��-�����������>���k`�*���yᯏzݺ�o۴is3�����l>����2N�	�tt����s����m|����pν�Ry?A�/����2�8�Љ����w���y����E��Z!Z{>�{3X��J9�1m�Ł��hll��pO^�w�)�X-�i�Q֎�)^�R�`]),u��k�](k�+����cB-N��'�:ߨ��P�\u��ФRD���e��<�ҥd���xcS*,"�W�9/�]��9�ܹ.��@Yl��9>����B��L��.�1�>;H�W���k�`��5���5��
dU���� ����{�lY�r9	:��f�2�@$E� �I� \�w�t���|g�q�{�����_sQ��ΰ��H�h� B��z2F�z����g\�F�!�,#��ռ	�l��j<�u�U�x��޿\.����ON�6���-��zj��Y�/Z�h�w	<
�}�[��ӟް��'�<zlllI*�J�6�r^�W�e�p]r��9!e�8ᚴ��Q\i2�`
�sP�Rb�;�.����:�9���> �cx8b#<�b.+ 7E}}�k��>�Kڀ�d��+]q]�̩�KƊ㑭�H�q�p�d	s>�g4�'N+�@�[��)@���ڗ�@Q3�3�6>^c�47k "p;��B�L�PYk
2�����Xj�3��h�� =m�� ��arqgn�J1���k�!��AN1&�D�h�i����:P! �]v#���)��3)d3镯}����o\t����?�{�Ϳ���[o?qKO�!�Ba�����6�g|y1����˵T������d ��[Hu�Z)Μ1�;'�~���-�_*�������ꪫ?�z��'��\�fm� .ȜdsC\$*� ��������ǿ��3�|Q��	�cO}�[348��B�P0���)���X(=��ݒ����P��*�TI�L���K��l��F�)]���U���oΔ�0�������Q��N��UըXq�l���n���F5��z$ȵ�B���,�*��'�3�����[����T2jK<3&���:�迩lp}+�}�zn�z�>�
�,�!�wL�yR�1B �e�r~m��ؒN%�=*\PK�A�*I��C���Wʷ�B�K�{e<��(vG1'܃bGs�po����<�@�-�:xյP�r�B��Rh<��`-�r�P�$�J*�����*���M:��g��V�J��҆iT��!X�m��<a��؍���у��8��1D�˰ߎWT`��}P'
����i�����uc;R��/��]�@���	?2X뢙e
HKIp�g[l&����}�Y|��^u���{��P ~��;�?��́�������:��)����YG,�F������A?55c�57z ��D)�3�Y�����2G�h��������u�cz���>Ykb�$Kh'm�2��P�^�J�׷���>��a<,8�W0���^��?c��h̎g������֑�o����p�L�d�e�1s���	���B\H��hm3P�U�}�]����`,p�9�s���?��(���$d81�S�:���X�z�������sz�2�w�,�Ƕ�:�[/���wu�Q�_��W����_����AJ�7������Θ���-��.c�&�x��Vg؝i��&&��jii����������89륀�������馛>322��鹘1$U� O�E�NV�Zi}��esݴ�6�uԫ���G>rϋ��'�ȝz�[�<�\�j���n7�=s�Mh����,H�ֆ5�ސE�`�V���:��M���ζ�Z���a��X�<aY-�#�Ԓ�Zx�o�5\L��LU��J�k�!��
�W��q���w�5�?]�x�3K �
Q�Ъ�Y�M,�,�h�G�΀�P=��]Fc�������1.�î�Pb�0�=����\J��a<�J~_S`�U �U
N�K)c0T�<~),�in��&C�Z���'�����5i���G�A섁�,� � �LV(�L&����P.�L�Ӄ�tj$�Ύdҩ�\6���Ը���ms�)?�I$�S�T!�L�3��T
��K�"݌]e����H��)����J�|�<�444�P,�w�JӋ�Bw�T�*WJ�b��R�t���r��V(Ӟ)���gg�{�[���0L�R�������\x���d�M��,�T���_J��0�cB
J{;p-����!+1�˭�m���Y���[6�[�~뭷۷c��a�*�t����k�57aJg�䎐�l�$X�� fڗ�T��ܼ 3"Di;�|\�a�w���� ���ˊ�f�*�\,��_��嘐��{�?�=X+0NʊP}�3����A�.T/g4�\�~7�o<GL@��IF'bP!9Ļb"}��� T\:A`U`K.��|yڤ˵P�r���F�[�2���K;gB�<8ݍ`���Q���%��rg�(/Y��o~�>��>mÍ7���o�������g���42v���2�sW�oةy�Ջ�h�����'=;����R�x����Ǿ�׿o��u�]7������}晵oo��y���`�0�ڶ�'�J��e��.��k�y� �ƒ�Zz�]#ÃKY��o+N�):c�t����>40��TQ�
�yl�B\�Y���X�,�&�ts>���b9�$Z
RcT(��L6oR��#櫥=����&V�4�,4(�R��Z�
A��g�l�8�@@Ȑj�^�YBG@@\�.T!�Q޻o��Ϣ��~�P��}��Pr��&���Cv+ �=U�EL��0-t6�������Gq�}LɝB�"�9V��I�2��BĢ�� (<�Ǝ������R>z��r�L&ݗ�dwd2�T&��ؐ����|z�)��:u�S�fM�5k�X{{��A4S�R�K=�k�I��D����SOmʏ�l�޶�o��������bql��BqJ�P�^/w
��b������,��0d\���`�R���kUw��m� ��Y�)]��l���v����b��hh�PK�����.����4�

�[�.�9������ȑ[��V�)�� ӳx)�9�s	aO� �� \pM����t+]L��u�5����ẖ)`i�d����bW���so��[��r>���
���4�\����8+�B���p>�O�^�8m8��7�̑R�Ș�"j���5y���1@} &����b"%�4�u���I�h���M-{n����Ii3.r۪�����X$�N�4���8b6X��o�RKK������xW2�j�R�>�˵Z}���f���-�W�X<�G�7 ~.�g�E���h���>���|��'ox������ˎ��;>��߿?�o��,��h�}��m��Uiv�mi~[Fg[�뮻|���z���ZOA|��s�	����g�9�J2���vjjZ�$S��@؄L�-�_�H��HTZ��۬P6�g#����G� *m�ii�6l�mڲ�@�-���	wL�N����m2O�������z��WA�x�<|�B�:&�ey� K���)F���>&*n͋~��X&��J�H��F��ps1��\��z@Q�-8&W����Bգ�t����Aຆ��a�H�A����6چ"�����d��E&���>�_.��8RC�t�7���hmm���Һ�����ٳg�6kּ���M���~��E��?ڡ�\sM�U�wl�������m��ch``�����RyZ�Z��Je�����es���&L�mEW,���6ݚ\�ք�-Iᄛ���c8�1U !Ǹ���F���i���>bdmKɅkN
G� Y���X�r�(>G�6�gn�l�����3�}�ow K �X3 M��m���4h=���3��}���dSkCu#d��(������TH�*�QǱ~4>a�\�n8�ix�W�A C��l|/&�7�T>�A���<)q��rV�73֌��>����6����|xƎ^f@<MWL����D_w�L��H�v��a�L���T@�X��W�V�r�1�\���c�j5O��\WH��}�|nP1�K���b�x��OPo����m#�l���,����7-[���F~����ӟ��|�I$� /V���=jeӵ'� ��50��G �rт�v���eG�{�i��/�%�L"�y�;/�����C�9S�z�5{FT'>�;�5s�u����iYg�ŚRlԃ��j�J��e�|&+e�L5���}F ORxQ2��vl�(�d�&�./��rMQ&��|`E��ѕ�F��]:��zi���^4����@�.��o�1�����ѩq�1![�yL6���L�p1i2�d)���~��m������G[3yӧϴ &̓>h�@�����B�RY��E�r]��ϟk��W�Aln���ea�~�C�t`��d�0E��,g��	ɳ�L銎<�H�~x�R)?����Lgw��,�y���,����ٳfΜ黺�/y}���e��jyr����Ϭ��v�}������6V�U�]R�T#n@���=�������ɀ�6���u%UOKd.1���bN=��c67��,e�5�XiN�E��b����`�������5�Pň(c`���K����`-uW,�'��-~ 댭���S=����� �7�s���֊�hs�9��:`�ɂ�Mu�ͷ���1?a܉��(��{���'1f@)�l!R�ώ���Ğ�|Js�貨�r�\����1��g���H^JAìk^s�� J��&7c9N�E���>�Q(w�Xx/X�L�\pO�G8�܇ߛ��j������SB�u�n���j�4����v�?�sG��_�����.�`�[n����>��_��g�9X�S�L�uK�ُ��\\��n����v[��o>�M�-[��ww?_�d\r�7�p��W~�*ו�Q>��N9�d�(?2��`-@�����H�<HHU--���0�g)\À�!�[��a崩&�o@�I���&7�r���(8&a.�=���/u[D�.s�=�~2Ӱ3�N&L�`B !H�
�1CNJ���r�pd�S��C0
(�.V�������e
�G�{eh�h1��#�5Ǆ"�����7��vП�B�*W�s�"�"XqJ���c(+� ��W�d�h�_S���Y$��m���=��E
8���`�̃�����N��R6G���������t��w���'���I����[n�%}�}�ι��[�<�����8/Ƨ&�ɶ����Y&޳AV�}�\�+59��_��G�t����p�mpu!3�hP@�,j�� F���H��������L΋o�&D�� ˽��#�&T���5a1�g���5�HK�[(��Q����7g�ʥ2#�A<�[��O����'A{,���Ş�v�q	�D����C��D�K�	�������o�k����aqC��3�2����O@U�R�0�e;k��Lx��I��W`z"��L�dx���#�Z6�c&+�v�T�?9�碧��d܆���f�<;K��>W���;�:��u?|�q˿x��>��Ȱ�����x��~��7��gHM�=�Ǻ�;� ����T� ���W����X���,_~�����l��y�}{}��tS6��5:4%S��oN;=�w�E�@ߎh`p{���ʬ�x�9�P�5�k=�T�:M4�Ы���Q�.�`B]ͱ(��}CQ�R�V?�TtۭwZ�,uR�MNM*-��RҤ�&��M�T�-b���d�1"�f������ �@P*�]���%<�nY�Z$j�~��\ks0�:����p��~���<�Þ���KOOO2��	���,y�Q���_��|��C+�v�p�YgE�w\t�o��P^���Z�7�}�Y�P?#e e�U� V_e�K����ن����rq�_���8�/]������?��S�����佲m=�&K�Z"B�朂Q��1g�xP��֔c������.�cC�T��&�����B*ǩ�d�\(=�^5�a���A��L�X�֘��ɫxz��N� k32Z�����Β�F����du�dM��vjMs,��a��}��C�B���� ��������7��=�Ʌx#6ſPK��(��j���2�$%C���r�LC!f�����<h5����1�����W����@� ��R}��� 1Ib�􊋍s]�n0]���u��u \�gkl�Mڶ456]��W��s�9g�K]�w�yg�7ܰ���o��m۶�n```���g�O�:Â�K��a� -֐{{��ǫ@$L�>c���s?�勾x�Km���j;�����سu�I�B1�F���Ï�]�
�@fk�Fc1�[<�+k�B'���&^�F����AQ���5�a�DƂS�nF�J4>V�֬]���ۣ�1�KQ6绩2�xM���8Km"f��v�S�u�Q\�(�Q� y�Q��I'���kD0p⺟@F��' ���֐"��@�+�{yE�ݢ���5���N����O��~xN6��`!ѿ�U���kOz�?.]z�����3o/�X.yJ�،��������\V֭����מUU�^�Y_��d �(�����#�oؚΤ�^0����={�9Ӝ9s^R �j�ܯs�}���~d��=[fn�ֻ�w��]|��###S�y����2��?K���wg�2�`	G�j<���e<�l#�ʜ�^��+vA˲��C��;����`�0Wp��{#��Y�n�װc�oYe���/�,��� H�f�u)`��P>�n� ���(mUMmC`�-����I    IDAT�<cOG��,e���P�(�I@@2����֍��'��B�C����
b,$�B�!F��_1=<'Ÿx'Ӏ�H����?zl����!;����������� X�9�0����:(س��k~A��ؑP��7i�z���@��B6��J�l-��ʙ:+�%�X���v��\@�k�ǳ�%{�Zݞ�gnZzء_�������e���f�����C��=~*�R��f�cM�-�&/X���]t������;�������K�oܗZu���8�>}�R6�@ƿ_�����~x�����|>��o�>ѫ������c;�667D�t*�[���r�A�+Q���-;�W%�H���T�R��Q�8>6^�F��t*3^���J�D[2J�fҙJ5�4�7WƋ�����j�6�-������r�`�%�Iɉy�Z���Ȃ֢� `r0���w����(l�ǽ>dX%Ә�eⱐ�`L<�����`da��ӀڂM�;FJ@lMh��[�,��А7a���]�淼�m###��{����Լ?�l~oim��]�z经;�5�������ի�qdd,X0%�=u�m���~��WG7�x�)�P������|����n7��gശ�E�Þ�TjcgG���|�:��G�,^�����k�N߶u��uk�Oٸa���m=��f���L-��]Q��EQs�X�%�\.אDp[j]l�n��SÜ����fA��S�y���e>�6ر��,�N��@A6�1�_��������1�Y��]���TI@���Ч�s�>�۲ys-��{*{�{�-�[�M�����­�I ����S?Q��u�7dX�B�"�?�b]
�͵|*�(7�b���Xl��}�u�DX<�e�y�)b'p����6�"C�ku�w�����
6exԋ�	����d%/��1
^ޞ6�\C���\!ra�]�w��z^�]�b:����S��'��<%�u�L@-������s���m�V���	όR �1�)�T1��r�Z[�~�AK�<��C�x)�-i����^�<��_lܸ������d���Դ��BL�v�����Q/�X�iq��B�'����w,[v��{�/\B��#�=٣�?�i��E�b�3�NwL�ڙ�b_�X,��RCKso>�JfңM��r6]HUR�J�\N�S�J&Nr�{g��t��.�J�T���-GKCC�����D�}/���oڴ��5��4Nj'�l�Kh�����(�b��� Ջ��"
z���bU5�$Ne��W����HQd
�b�`��2l�����5��S��ڂ�w=�b'm�5kVu�]����>��/s����Ư?�n�ۚ����:a�s�~��_<�j�?��/}���\:�]��ߟڼ����ם�����}�]t��6�=��/&�+^�8�/�}�Y�gώ���J�]/�%��/:���wo���;��EL�?�C��j��k�����L�G�m޺�U##��+��r�B�CJ� AjB�Y�e� R�a<���	3��ص�6�
�@�B�Z�Ж�ؘS|�pUF��e��jAxR>�����؎8�^A�
B��0#��]�:����f�奲�6��j�x��B���ߜO�����i�)\l�b�d�R�P�1��\�d�n�=�\�J\2��*j�'��\q*rpm���0/b�l�J��-t�%h�:\R����G�F.\�+Q�3j����ދ�W��YXj�W����g�rsɸR�M�Ċ)����b������	�b�Q ��֤��u�9�L�g�y܇�������vc鐋��-@6��
�If�!�ym_����:��TK�|>����n�5k��N8ᘕ/6�������y�mo9��o�ރ����Z��?c�4���fαv��ز����%���e���X�l6���(��6���O|�g��{o��3a:d�IH��ш���w{��'��j��&~r�L���$
���J�ңr}'W��k'ZhJ�
A�=���o��|&���	ʱ0"U՞*(��gYq;8D���;g� �@~���}�kO=�S���[n�e��>�K��!�t:;<<�_�<�����/�H]}�W�ؼy�T�:s��G��'��e�����u�]�,4!a��GM�:��SO>i���C�Z������r�g�,����fM{��-&�>'_J������OO}��{�_��U�7oZX.��D�Č��B��5s�#l:)RiwƽT�4cX%�RhΣ`�o�1P�^�m</8`a��|_���<<���&���x�Hs�6ln�A� �������~�e��\�2Ǫ	W`
�$ӌ�ɐ�������Rq����A�X@g��(�璛��^m�L?B���`:�u �z�.�����	'bp�^�C}��Ԧi��R`y.][�HrDl���|�L,	ó�։��6m�s��!7 �T��)��{��=#�ϕzK_�%�8�ɐ��s��i��u�n�#fKL��_�E�6��a�}�6�� *�J
����$�	p��r�i=i����6�Q2jo��)Y����t_gg׍���{��ﾻ�9}��m��6���s�w�v�W��l}���{���6�<��y�S�L�����]��	K�Pm<���ܚ�\���h�9\��.̝;�K�w�5��j��=��d\�����{W_��R�Ҏ��N���D�d�L鶼d�4�SD��u-M�P�K k��c�JS��h`&��s�d����oϙ	o����ߩ�X=��h�lzs"��T���|n��{�y��?���������;V�^����%��޽�5�y������7.;�G?��7V�\����%�d�+��׷=zlժh�]��>��/l۶�w��y7�[�P���F�~����z��iO<�ȾO>��1���+��̱���t��ؤ	,��$���=Kɭ3Yc��O�b���/$$ �ߜN����8D/s={� L�&��{3�������ܵ�K%��
���u����m�g�̦�D��Xp����!�%լJvb�-`� �g����uw�P&��C앀����T�x�9�"���eK����3��]����5+�����P��UQR�5�\�K Cc-�8tx[<ND�A��j�g(c�vlﯥ�Obt�]X�JrQ�H�ՍWŬiLu���� S�?2}.Opa��s��X�bPOCr9�`M�h2 AQ-��x���J*�� �V�G_	�i�(+�p)Y�;���������,�l�+��y�G�y.�Ɔ�Onx���G�u<�fu��O={����_,�����1P&�� ����n���`�z)�6>4#$v�>8[`����ۯ|呗�z�I��"�e�dP���~�/�J�P=��PB���b� ��|f�1h&<��Κ�4e.�aӽ���-y&vcN<P����lLF&�,1e�(]��B�.H�J0ˀ�8���|�yeG�E���v�V����)�ox*��ܻ|���Κ5m}GG���ŋ��Pn���r�Gn����X�rU���!�;�0k�#���^��W�x�߿~�v�.~E�\sM�-�ܲ��GV���o��j�:7�J5��V� �Z���y!���C�:e�EK���)�% �6ב7����!H�9˜d�]徐�&�LsT>v��o(>e@ 2HW���5�V+e�K� ѶPh��������l\xѾ�#p��w%�6S8�7��J�uY`�(�r��6�j����zp�S޴��g�Q��~��H�L�;��L�1�W�U_�
S2I���!���� ���
�4���m��%�hH���V�ʣS�Oʕvi�2�<%7��ԷRpV�EL��O��c�8��`����Wf��������vH�>	H(����Љ�A^�L�2�>.�}���X1�+��J5D�àU��@�����]@����s���yǢE�������+W�[�q���?��k�ث0R\0^�9>^��dr��u�9XA�D\;�h֬��yƌ���\`�L��T����dkj������@��9� �����y�{���/+�A����o���u>+Z���Z�;{����wFmln����J�pI��U.��ɨ`7<�5�1�	?���X��|�Y&1�)�Kv�v �
dA8�g!S	 b5D;�J'WϚ5���{��{����o�c�<���-?������7�}����Lj����q��Y�t�����/}勯�c���tͫ�����o�����<}pp�J����|�vSUlD���@��j�U(+�9��OR�[�:n=&Is�Kp� q�������V<O>u��Oh��+mYЀ��0m�n��3�����5<8���!0�ʜ<`ů=K��f|+{�o ,l[��#����Sw�{we�F/Y�\ۅo=>��M6J���k�+)3N��û��'�;ƙ��[�j�59�Z�\G��\�N�s.���D׋������<�[��<1)(8� �O��S���ೞ���c�?�m@V1�㽦���b4A���^����eq�N׶�"����{�Ma�n��y�A1\��Tu%m�1�|c�T!��, @#����k�\0�4~���
lU)�����--W��=�y������}�o�W���'ə�Jij��i��p,*%�6�/^޿��/ĊЯn�8X���<��9�;c%�T7���-h-�r�;��s��O9�?}1۴�!���d��s�W\188�|��#��8Bƀ�jJ����ZZ!�v�����/Ƃk˧
 �"�Ž��,@�0����|Q����ǟnjj��ŋ�w���޷t��-���]�X�jՌ���M?~��G��u���f�r��>�+�A���V�����n�m�c��O���k���7_q�M7��\.����k���:&��h�L\R8g��5_4�u?���IP����Y�r/��}��i�Ah�jŷΖ�-?:�k(K^N������(}Yݡ��h�R77Z���d��%�(UU�^s^�E֐���K�������@�*NB ���2Y�&���,��y�^π>�ڊ�7#����%��q�0�o��
�HQP$�K�U����oj������Pyk��-��c���.����묮��m��L�&�82�I$�%)�$Vkt�Y\Q�T��R|<��<&6#̘���8T0�'+�8�w�2#��k��.��'�+����̕��b�l-��Ҽc+
h��	� �^��K
+����������l+
l���(����������LG-M��'ʄR��I�|�s+[���_j=[>o��fWtvu��駿��˗/����'�_v ����?=��G=�P(,L����j��H�=[-&��"�q�)]����N��R)��Ҝohhj{��'jnn�U.�l��jSG�JY��L��z�+��I��W����zJ�rO�8ޞNg����ǆ���##��S�NM�R�͛773y�N�Z����6a�R��$i��[:�~����7]�q�ѯ���O��6�y�I0��իWϺ�'7���SO�w����
OQ�ӧO���:KsfϹ�k�|��/�^/��/��yw�}������ޒHDK��d�-;�e#@P���H�H ��)�!�T)�$R<�NYg��!:���q?��&�?#+_B�/K���>��-�%�f`�z�)hi�@���V^ E�G���.e�gV#��ˊK������#�Xs��r�3�,���(�����|l����c4�.����o z� ��0�H�ϑ�|h%�U��"�A��M� �o�w��F�$���P|��� ����D���V�(�� 	���b�A�\6��v�@�\II��2��А#>��Ɖ��\0\W�bqx&b#�,���yW���܁�a���K=���+^��������(�{��(�����cLQH2|<eWc(@(cV�N��P�\�ˬk�C�B)��Β{|����!����1�Z������Y���ؿ<�G'�|r����}Y��?T�]s�5O<�D+9�ccQ:�'�1]*�ք�d�Z�T�
I��t�Z���|�Zi-�˔�[�h�U�}�{W����y�m�,:�����k���~~�ҥ����֖�կ~��r��>����|�M�)K�FF�R�L*�H%��d�\����\��ᅋ��ᤓ���E���o~=��������ܰq�!�d�]������S�,�9s�l[��ޟ=�o�򕗒����/�v�����r����MMMӕ- �0F9��w�Jm{��&��N0�TuKE,���	��C�8+�pI�Ǩ�%�  �K��
3):��Jo�����h���ӴIU3yצ���fA�x�1ZS�b !�K�JD��N��GR@\m�f��6�B7e�~��"�-k]n%	l=/�Vl��0χ��1�eP��'�W�e`!��b3Ԗ�QИ<��g0�?큯:W��N���Ox)[	C��	Le�C���D~�e���؊��1�'����j�1`r��]7:<6)&��c4��	l�Z
J�H����>њ�+N	.�d�� I�<���Y��Ix�+��¼�i�G~�U��ܛ�7�y���V��\;�˕�6�cY��ݓ�OsH���>q\mpq��N�R+gϙ}�I'�p��4��s��/Y��N�5�����mmmI�{ｷx��'���!����%��p�W/�r͚5�n޼�����M�+��pju֬��{��Շy�%g����m���&)�+V�<覛~�����#��l���OT�����l¹��ݚ8���~S�c�N�z�g�$LD�"��2R����;b ��7;.�MJ ����E�,Bh��� yi�0��7�j�)/ALl�!��^e��5�=9O F0ڬ���s�3�W��=Dx�b��N�,�PًRW��0#���{���>���"�{�)I)C����x��K��P�����=��Je�T]V��%][.#Wz�V���ź��>����X^b<��ʮ�fw�Y��_ @�.ߩO���=��On�mŤ� !�������('�_�B�ɮ1��d�h�	F���b�S��[�b��] ��ȸ�����P�a�%�Z�b7��Ԝ�55O#�qu��1,���.�r���Z�����_�l���O�E�K6�d�Oh���=����o���{�M=��ѳϮ�����-�k����3��Ϗ^u��W|��-Y��e���=��3�;߹��իW�90�@Sc�m��`b�����
��L\�jk-#���Q����R@u6�}�\OԿ	�����d%�(�/+�c���,���:
(�0
]B��ǄD���!��~Af�A���3��*(�������().�+�r�Yzd�(&�����L,��K�-Q)#��!�B����hn�j�,�P�� �t���,�l�,��_ŽB�]L����LH���4�K�0�;{���[��|�(`- Z8Wc,��3�e��/��da�8�NI8{�?��d:�
��D&*ǁ�:��0Ł��Z������vR�S���!vO,����P	k��=�g�$�g�Gc���rM�� Kk�[�o�Vc�bw8�`�T��hNO��=�cc����3�̶���;w]��w^��ew���'��c�^���3�x�=����z�Y�_���l�һ?~�5�%���D��O�P@�Z,�T:������?���w�]/�.��.�˫���c�\�M�H���RE��Jt;�0�T��|�q����J���R\&x"r�Cy�*p��^��(�	�
�w�Q�`��N���و�Z�y*�#几�����JF�E�,'�E�4/Lvv8��D�3��`��\�Km�o���A�BpO�){�:�9����@��f���x��vP�
)�uޱ��� �򐵍[��؍R�v�)���&�Q}�qw(A����#*]��J�J5�{I��}�\�WVȚX")�)�P���Ř�\��B0�i�ޏ�i���ZrE��_}%�!dz�7[�O>��P_�=!���A��5���X	���������K�S`p=�6-r>:(~    IDAT��!8`����]�]���j *ᮏ���>`S5����t:�&��������}�C�^2�� ��0J�Cm�袋����G/d�oܸ���u�j��߈~tk�I;���LE}mm�����k�<��{���7���h�خ������=[�_�~�	���Md��"��O
�Dy�Y�&�1�����^6��[�̪.Ĥ<�!���V����O��h�|��G�n�*A�5�xa����k�J\OB)�P�f!Z���
d�!�p� * @�1態��G`��(C<�`�294b\��=�c�3�����ϻ�_t�2�,Wj���1WPV�����"���ewy*%u���%�!dq�xР�TMQ.|8�g��2(T�k�)�Ul�Ȩ�H��n��~�i!p�~�+*jwp�?/$�)�q��ҕ��� ddtCpU q��'E�F���y�J��.?�w�))]����X�������q�#M1g�c��D�����Y�7W��|4L�NԜ���;�=s���/��S�k���x����20*�Ħ����:::n�u����W��O��|2�� ��z���<�������n��v(�zy��u��(��e�#��#d9�၅����y�C���������e˖=�|���T���������𹮮����B�W.H%�
�g�ٶmB�Y�cq��5���l�iӬ
'BS��1����r��;�	)�*�����Q	WY�
���V�>m�,�D�8n������\���l�1������bY�Y�JUA:����U�|cM�c~������E"&G�

���#C�\�R��ഗ�(i�3
u��`�Y����{�s\C�,:(�����f}e�����#t���_����������UH�y`�c�)V��Ǜ$-�7�%�z�+���hs�ጚ�'
���1	1P��+Y�Y����K��٠���"Y�b2¹���b|�wM�z�YMڊ���h����A�#!|���k�MtҤ���g�4�t���z�i2��T*�����:�o?p��?Y�t��e˖�����ێ?���c�ˎ��o,���{�*�-,4� bbc��,YD��h֣�>�qFF\����D"����{���<��E��]�h�e���5lw�y�n_��W���O�����Ͷr+��`�
���jݺ��z�c��EaKAʢCL��U���bG�(�w��<�K�#{�G�2�5Op���B���F�ڕE'z||l��A���u/Y].���K �
�"ӵ9BIB9��x�+mV	��ŵB�\l�g;N��"�2�or�T㮉\��ܪB6O��˼�ZR^�{�-E�|ߓ�ˁGR1��ꪫ�*�ִ��.F3F�q�	�Yp���	�EE��3/�ɩ��V��i�P��s�;3o��믫{��Wu��ǰI�\�b�y3ϴ�^yR[�bS��lH�+��H�g�ﷴF��^�}Y��qq؞�s"�Q�1�N �*vE�$�3��NV��-���]�2��'\q����1ʅ�0}jw�v���\�sL��(�e�Q0{Z	��"��G�ɑq��d-f�ۑ��1� AQ!]cHܞQ��������!�������JU����2�g���TY^�I�m���W��>�aSq5��T��ot����a�.[����R#����/"	v�`���\�>�jJg���A�2�HĲ��������þ}w��6=�{��z�o���^�m�cO=�v���y`�	��WF�}��k�W	s��w�t�b��Fu�؎?�\!�� 5� c1��O���'o��)`���?�i��J��s�0����FtO�,��4@U��V7hu.���������]���v_�\{�qX�t�v���ُ�%�ǹhɞ��ag�����%�/�H�����b�`0��զK��̑c8UJq=`��j�� :��� ����ϔ����~���s�t �.��y��:�I[�� d�>Fa�.6���؁ª�zU�	� t�LIj��z=5�;��[	y,r*��D펟;�y�(�=�D� ,P���8���y$wG%��!X�1���Q����� ���{�=��6{<�P(\��Wd��Y=zl��>��~����7P�����9�Mi؉'v~�_o�:w].�?$�f@C�΃?�\�s��/?Wa���T��0��2.�����xEEE��:��ԩ��Ν���ҥ��k׮�`0�VRR�ԩ��D���:G�u��}�&�������t���H��j2�Fe�Ca/�3�P#�+L�#�ҧBC����&�v�b�-�� j�G�p:~��l'S�I�J��\�D�z��ag��(�L�N�%�PS�A�1 �]Z!'��	z�h)�J��&�R�W��5U��U��r˨�����2�B�\J�D���+U��%<���Ϡi�sƽI[�Z���%�fʡx]RZ$���h�.R;����� ���TQ�;A��D���5��p�h(��=��)���4L�8p�o����KD#�J�|�W��$=�5G� ��B��=�@�< ��dM�\�q��{���E�E�eœ�%e��L���������c���$��T��f��l.�3sa���A ?_6�����p�d�\n# ���0\���x�\6(DPw,`��^�c@��l�@���b�������aTĒ�_-��q�i{�f���p�Ì�\�v�����V���:�p-��}3:Wu���V[��M�x�N�\/H?�'r�mꀌ�f�M{��+W=��S�L�f�e�t:�/=s�\�h����`�0�?����:Aͷ�q�" 㐅�>�w*��e3���z<�6�����mE�E�E�%�%�+��KꊊB>_�)���K*+3.�;�v�s��Ş%Km1}����ZZ���zK� ȓ�J+ԑƵ�?ܘ'��|����\"Y]� _/������@)Z��d T�i!\�hI����:}�ǪMM$�p���B�'�@�N޾zsY�$��qL��	j k�#��*�*(�R�@��j�t�\������VP�$x�5�6��
�\1�������0B�� ��`5�*LK0��m�W��-`_���y��rK�P�S�\M��~�u$%�
�D<i���Iʈ)3���/R	6��E"UMii�s�8�K����`�LNW܅���?�����KtF�n���ˊ4�s��"��3�����^���x睷_Խ{��_��QБ#��VT�����nw���������N�R�L&㫭m	�r�h4N$"�D"]����d�$��UfR�Rӕ)N�M�˕����t�|��ș�`�f39������!���v�\�va�
���CQЂ�BhA�vgq٠������i�\IK=:�u����*#�v��������^wSiQ1~k�*�[���**��u�V��҆�{��=�2���Ȏ?��k��5{օ�T�#�N�V5PY�I��$�М���T"��B��U�qcU�g���g`�R�XErf�Z��L2�L{<�,d�s�\1�����É��6p&R
z�W�Z,�# �sO�4?Ng ++��_V�ՕUV����#��ґF�+��^�X�*� ���hM$4�D���0lMg��a�}���D+T��\�)I���zW�X&a~�H,��V�|3�M�+��"�S݊L2����:�A΀�V���My���!U0q���~zo�,4�m�l�
���|�����q>J�S0���y#-"m�^������mq轠������(�F �xy���ڂ)��Q��^�%/Þ
��m���qa'��țO��+ �L#�{f�(tuƗ��v��z}�<^��-:w}{�=w�r�UWm�:?�	��O>��V 	7׆�qW�����݉D��v�}��+hIO&�a�͸ݦ;�1ݡp����\2
�r���0��2�:t�e25ي�xfs�@�-�䀌�e��h���{��/'L�9���Ji�O4�A-mdYK��аz�L�e�t@$������ԏ`X��=�?��2�`}�{L��E��![�
���0�y���:X���8�-�z�C@�p��yΊ����ȏ��hl Kh�D��2�x������Gm�
�X�8ނp��C�6�j��2"kKS���ƌ6�f��4�RЦ���V���Oer�N�6s�ۂ 1�ӷi�	\(�U�������b^+�GQ�FH�-�RH3�N���W'H�ypH��V[m!�ù@��>�����`��tJ�R ќ�X�i� ��F$�&!H��Y�xY^L@�Q>V�ฐ���`'��1�/�_97�҈�~'A�4rf��2Vx|���᯻u���N��4ذa�q��l9���,����d�����;n�_xvX{[�l.�)��
�n���c`�LA��j�������N\�/lXTj����
�B+d�{���l�9W}xM��N�ز���̩�	�(@�-�hą�7ҧ �Q��[�.�Z�6"�q��W�((u�$�JD \pR�#	EP�7G��b�``[��X^%��J��"- ����-[b��4���@����0:Z��a+�[lX`�<�#�寸f�LR�2!ω��%��^|����G+$J����ƪ��Ag���bd�y����#!ꔕpg��\p�O=	�+Z%�KEE� ���N���(ȴ����.)�����I�.9SZ�+��%���uW�IH�G-EZB���:�}�q`�� Xʨ���9��41�#@%�����e��I"32iH����B�E$ʣ'�T�=��7�Ls���^����nѥ�;��ܛo�������9dl��m������咽�|ٲL��+�Bt�\8'63R���Ñ�	�81�X=�Y���u���� 0���AKG'�V�EXU�Iӵ����<�������G����^B햰U�\��9��#F��X�&Ǌ��t@�<��`���k��ح�_؀?d��Z)g
Bb�-�U�F�(l���Hy`E��!ڠNUAq!BZu'2��R� ��#�����hX2��b� CW����7��1�V��%����X�1�ư?�y#m�t# x���}t"��Iu�J#*6��C�ϫ.��H��T�	��)��ĳ��[�#�^PM�CWR�Nh��`�q�b**=4�Bm�|�ŭa�$,� yB�5T&\�_0^,�0.�o)�fe|�p8���{�u��Yee���f��_��խ�{��ѣ�:j����`~؜��58 c��r�h̘����N[�d�L��K2�=�Ar�2��6?��Ѥ���-���X���J�L����:i9;��xO���g��j��S|����X����z���\ � ���͒gt�	E�J\伷꺅TM dH����#E��y��c	'y*�E��:$-�N	�@�@D�|>��#Ays
�X����3�T�5�r�1�q�h�pxΙ���p�LIX�\(K��A���J%�
v����	��+���Z]�(9,$�2m�H���Y�~j4cV i�b�<	Fmt��t���#'z,hx��þ8&8;�~`D00VYYY��r���n��|䑇N�������9������-������v�����]�pрl&�c2�,g)���:Bj�$�~|ƒG�L��+#tܚ^A	�F�n!�٭ �^:4���7�Rط����@��[rO́� � �K��ܲ��ݡ� '�h��r� i�C�d�}@_�^������8;*]bL�$���������h�N�ﶶ�6p���`��U�B�<B&T�XU�J�8!�Z�!I�Jc6[���J��9����P�c0"E�R�N��z��
(�n�85)%t��Cz��2�G�*�	׋�����k�ؼ�I	�T9e$�~��� ?)�P����?� I�����a�DB�' ��p8�r��[^Z��Q�\;z���-���G�9ݍ��ب.��3���TL�2a��L9���yߖ�D7�\��r�nii���\����24 2 ���;�`�N���1{*���#܇@���*���ʅ l'"�6�l#s�&�F:�1�x^�Q�}�C�++C����d��N	1p޼y*V�R>����X���0|X۲Á!���;���/5!��¶*��+M��\��p�J�q)iΔ�D5��K�%6+Mp|�U�t	��
���c�q!��b~v%�t��XHT!��I%Mo(i����� ����f�*p*��s�C�M���$²?Ik����v����8,��P�ʟ��M��|Y^Q��!�3��+�n<��L7w8 cs������'[~���͜9�H$�]6��:��i*B��C�.����F���`�$<J#�
2
i��;E8}(o�._T|��6��S$�����X"�US#�}y�r�pY��(�9:�V�H�`,8<�p,Z��jO��@�%�ad�I	<���;_r�Wa*�o�<� ��́\�|?	��@��-G̴�b$�Dy �d��i�V��:��`%�v�+y]��aHKZ�����J+��AR(A�d(#��ԑ��tYk�-S.G;�"T ��~����S*u�/QA�Tk����~���n���K����9�c��jd�Us:���L�����{��N��}ΜY'466��$z%��D*H2ď1���=�R<���K	:29�����_�{��c�
�EaZ�+g����s�88l+Q�2�g:� �=�&i�귺xb<8��b�	����	��kn��[p�(�a٭���R$E���FF>�`��A(/�-+{��<�B8'T� -�T�����*�@�l���A��s�C���~���h���l'�b7*NP*�`K�C��O�)|�����F�=Am���>�S2L�ډ�7^̇m�4D��q�pP[y��	�-T`p�P(8}��}.+.�{����q�628 c#�`��t�/_~��}�o̜=k7�۽e(��ek��OW�*����!X�"N��e����ډ+q�B�I����P�#6��p?V����?:q,uVi	���5/]P��$��hkѕu<�-��%M %J+=����'���p�t��\�~8��ᡄ\%˒#���t��?V��Ƹx�^�/���Has6샨�inn�W�Ў�r0������=�u!QV�K�?SN�%t\0����8>;Sd6�]0rsi��)�UT����\G3�<ޗ���G!e�H^���#;�����`S��;��Y���5� ��4M��X1oޤ�3fo�t�҃��N%S]À�h�ae,�#(���C�v�z�����h\�H�x���>�,����h87lk����k�� �����Y�,:pp�.�3�N�V,$�)K��_��]n�8G���t���ܨz����!��(H� ��Ab�@�N[���y���xɳ%/`A	u%D*�a�#C��lsn�� ��N�Gm%z
MӨ��k �S��4z��^3�1�A#jx&0 9��v�0+g�"O�C(ΓcC᠑ˀ7�hQ���$}��t:��m��t�^{�նA~a�I9XC8 c�l�~,��g��,\��l��ť+V�w��]ѻ��a�h{[�D"U�m�4LO�i�E�X����np�J��*�B�T#JB�'	^3�/�H�3�ʔ��/O�K>��������	�J�rW�T�\S*Y�h gJ'��t�T'�=Tg d�A�%���;	�8U�T",�5����%�P�����@�$�.�l	ިH�T��j�D , xpn�mH7Apet�:P$ �g�s��+AH:�)����Yi��i(���da��2`�����v�A�7��!nC��Ϩ��F�("q������ �	���nݺ�����Q27    IDATL���vg=��#�Ϸ�9�c��gd�=[:#�c̜9�d��Eյ�WTΞ��s]݊]&M�|f[[�V�ب?�\��@�� �
?���S������N�az8
{?F2x|��I-DW�F4�&N�z�W>��.���m��%�9BO,n5�bڂ�{��p$,r��zt�.��Kp'��LjTPQS�3�&@�=�C�(^ϝ;7/���)���i2i�Z&jWeZ��Jl�ϰ��!�:��#Q!���/\�������I��J\Kr3�F!(`��>"���Έa�h|[2M���wd���PWoTUW(I�-))6rfv���g9p��e��+�α�Z��2ֺI�ק.�誋>���rE�B�UD�2Sѧ��ހ�cƊ��T8Tu�=�������p�"n%}GT��\;I�ɹ�d4��Ϊ�p(i��<N%����Ph�ș��@��(�%3M����RMF M '����A�q؈�yv��-s1R"�&�ϧl(;1:dx4�Λ�S!LM0����u��ؙ���oo�J���nH��QW�2���5��h�>-m�j��Y��IL���{1b��p� h8gF9p� z���}p ~ .�Њ��E��<"Z=z���ε��۝���<�>�Gα�-8 cmY�g�Z����2kּ����G�,X0�0���� ��@��j��>��
 � ��b8&���<H�#F�
��Y�b���:${����	�rHc+8�}$�5"��pt�������Ao�+!p��+�M�yju�*zbŌ�<,��`�ȅ�lX=g�B�q�Z ��4$�2� �{`�z1�|�.�W�4�衪£�,�d*��ؼ��K>
{�P1��Ɣ;Ғ��% �jJ	8y�ca�x�G���O�Y`,���P�#���l `������^�E�4<0�J$�-��BlU^QjF"����!�~x�z�B9w,��,����dHg�uk�4=��2v�o����W_}hsc�����[4k����dgB2 K�� ���������a��p�U)��p\��  U�z���J�#�<���j(M�����	*���,^4��Pc���D4�v�c�#�Y��!��m ���E��$�M�>�`SH�����h�-�a���W���~�H�,
���N���"=��HBe��$\���+G��ɳ���5��jj�eNHQ`*��j*E#&��y�v #�4��<y,J��T�1h+V�`|��p| ��,ZYU.s��B�U�����~��c��w�z��T2�UuuE���m�j���4��ч�oݺ�69Gs,��Y���m�����[}&N�f���g�q��%{��E�y=����5v�e��o�ͯ�:�m
�_B�p 
pp�Ŗ�%�6S#  pV� ��r��+!SW܌^��8���e�
I�   ~��IE ����ŵ`u��_T��>V��L0��Xi pI�-�+����$��ŒE�%�Fc3��_A��{P����U��QB'���+V,�s*� �)!����\�`5	�% ���4b�@�U$*I�)_��qN8�F��{/Q�!6S�֩��Р�M�EF <�&�30�猔ᾁ��/S$�d<]���T�Պ���ٮ�ŏ?��~5�z뭊��:oqqq|������+��X`�Z�����������O;;q���;j�E���mg$\���@�O�>"���5>�#@� ��Q����RMt��#a�$�'@2�	��g(��SL�أʯ(H���@'��!B��tJ:ע���X�"��N�L:H��׶���8i���-�SX���`�58a�K	����9Q�~����2R`W�$���D�T��H��d�q��F/p��l��HDcy�C`A`�r_�����0JU^^)�����e��c�Z��e��p�\�B�K+DymXu�m1_�ၹ�02E]���ƈ� �)0t�]�_�~�ݯ��޻>��{��ܱ��ddlJWs9��'�z͘1{�ys�Y��Ч���G4�,PUp�pp(��e���;"�5�� X��.����ꎐ�F��*�߳���Np���J?�`�� �%��$����4]WTm����.����֡A�;%����.iPJ:���߽����s�Z�}����d��y+�����BL��M�Ok$��j�vz(<�$��H���_���
��hv�_ǅ> Ѿbhg�Kܑ��f��9c��oeXi�2wè��߁��U�I*v	ث�IHJ�>���<MM�$qB!��v�9��	��^�����Z���A ���V~"Ll��a?ӯG_��u��`�4�w���،�����YRw(�x�8L4��G�����r?�>F�m�Ǳ�e_>�Ԧ��NAv��j�����Ji�?fg�~�M���y&Q~)�T�I.B0�D�l�"20�2a| �g��B�D��%�H}���h3f��.�G�ط$�h�F�?���o֥ vZ6/t��l,'c]F�փX<HTCvJ|ku�t �#@N��E7
�CBS��An��KG_Äl8V�^�E�" ����a��ҵ�^�t1
r��oog����-��b۝v��$����ԓa�){������;l���9q����'��1�݊�f�: J@��eiV=�P�r�-^O�������o6_E�t�?��B�$��V.ձ�to2�D)uL�:1��f�߭+�3��������ieo���sM�x��{��!��5�g�����<*�sGE�G��1�/,+l���}��-z���"P슊[Qr�,>F\,��^Gk)G�F��?	
{�gM� ����F��=�$�.�R��pp<��xC������pƏ<�4%�?��1�ɂq�λaC �!�0���إ@sB{ՇjE��a����iu�滒���N�?����Z���혬\��x�h�Ē����pbdd.5�-}{��ȅ���yn�f}�|2��������
�8 h'aQ�=ZZ� �eJKX+Nwx���(W�!��l2a�L�:�}�,s���\|�Ҧ(��퐷��jc�5�{eF�<ݟl������e1y�WI���}nrm���m��l��,z =J.��Q�7#��H-�X%�n��,�d��Vrp+c0r�veq+R�Sg��i�����IKڵ���l�A���.��H�bpb~��n)���A�F������늹9/��GC���
��$�<��,�����,T���6~m,i2��Ȝ������N7-2:�L����O�����_��Zk~+K���uD�R������ء�I�0OL�
���ξ��$��|d����`#Èp6Y�t�Kׅ�A��H?«�������*C�h7�'�u6�w��V�z�B���	��4�O���`F��-������Q
��ۻ=�}s؆�C�ODmP)�K��55N3?~�(�h؅���	����l���K�c��D�i`�Շ*Ƽ�[��ڒ�"l�R�zt�ްD��!��)�0p�o	ɚ]#���H�Й��^��h^��*{�ª�&"��&!b��ᇧ����Z4��q�(~�z�}���
pAU�05��5+�h�<&�f������e��J�֟��p� �(���Q�M��� �����[�[ヘb���0�W����-r	D���Ƶu�:^�'0p���?�*+C�,alw�9����f�Gp]>_�n�a���NA}���P�p�����0�!r�����l���6��H�3$����M���*�7
�'u���H����������UQQ�\�f��#��N+n8�7���,�>�A���G�
*:ݸ4,�u_2���3��)�������e�Y�[B�&ϬRۧ�U��lH��[��d��8���b��o7cM�zkYE�3=obd��韞&�׻
{q1�O"���C�\�@J8�`
�tp*�tb���dm�_$M��@����0ovDQy{g����?�>u_����_�L����-?�.�TJJ��~�2�$�.�Z��˂'3P^�`N�����%wSKx�>x��F?I��x�Y�,����U����܃E��D	��e"Λ���}�3���b}�]�sO�ES ѕ���/#�^Y,��z�y"�~�hC�46����䗼����}5r}x!�ֻ�B�:c+����8C*���t��n��/^�5�:wK}�ꁶ�d�����6m��-P�F�J
ЎE}�i�[r�Ɨ���NƑ���]G�B��=��bM�m̄w����pmM��1���8�
��;S�C9�8�~�hg1�½����,�G���?*ƍ�۩�:���tvz=�m���y�u���s����V�A=�}Kb�Y.�N����P���t�����g��ˇ}
��s�qD��;N55{�;���fl	>Q.�p
 �B��	u���$$J���v,,U^��Mj��`�x���,pp]�/˙Y��� 4���^���q��3B �1Fx'Gǉ6,D�+2 ;��"j��&��م`,1%*��^�͕���te;DYe,q������	�Z��b0���ղ�D�/��T�g�&�A h!�Ѻ,�o6�j2.��'�	`c�s6Z$B��q`�5G&ӷ��ZQ��)�����&�5���0�,|Pp�s����%Ҵ����\����n Fߟ�MϾ���F��������ꌱ�@v0Zl� n��/�� cF��)�nI�µ��f�>b�>	���F���=�WT�I�٤ �����58A�o��ܬ�+��T�?9E�n�8��Tݷ��=l_cv�W�z���O{������}#�C��/�?�z��(eh�4Az�s��ٔ�H p8�r�\<H
"q�}bt�"�ѥEq�#�>7�!!��Xr�U�r�r�c�k~�
����-���hR�� ��`�ña�BƧ�͐�3p��E�mº��[�����Z?F�2SR�8����K�)��9���X�� ��P7�@�|�}���R��9;���q,=v�-靓�~�e���jE��X��}�V��]�δ%:P��ض��x��<��.]N9k�u�@�Y��ٹ�H�{�t����T=�[�w_ϴ��w���~sb�-y?O���^S������;l�h*�/�Q���a_����_J�D�ѷ��� ��rH ��V�|������4$�����A�\]N�	���Cr�0��֌��I.��p�Y3� �kO�5�D?���Q��Ir�2����DR��(�W��g��I9T��	����6&O�0��\*tX>���G��S��F�[�H����&Y�W�d��HX_	�Ƶ
�8�߱��(Qk�L�J^�\��@���x�9�!z�Gٕ� �_�f5�����H��lgd���V�I{�Z0g|xg%1_}"��d�k������0�*�Y/��Ql�VS�'� �CZ��{G����H����K��<�_��r��.�>��O�7@V��i�9���@��x����y����A����Ʃ��Hg��1���6o�AU c�}A@��{�o
6Zl������5]���ka�����0s"&EͮX���OV0|�{��D�F���$���~.��F e�g(X˷W�خ�v$B�q/fUbAָ@Ke4�)��Z���]kKs��b:VS8��;��R3 !���&����{��%B�k y���}��{�i^*ϭ�ϻ�G���Aa��ҷڷ�`�.�s��L��޹���(�B `��������c�M�w?{�I�b��?Q��'L��F688(��%h�r�W:�D��m(�i�7=�3�o��	�6�����y>�
�Y/v���ո��$�uA�~7[� >z�I���+s��]�H
��L����$�55��hC��B�e\D"�̺�f��~q�/w\��}��tP��R]�����Q�z�(V��7m��*Y�zQ�1��B��Sڸ\�^ק8TZ3-1��:�S�,���+�R�-�:����?Z+�M��0A��_�!�]Ƚ�=x�m�����}�G'|T�u�y�}���#4$A��[�/��|�)��JfCmz24�4V+g��m��Cb��mz%����5�맦K�ڎ�a[�N=�$�a��uS�Ex���D}�� �Ū�O5��Cj�d�:��۽�rE��Hn�#ݯ��1���i����W���oE	#�wW�������AnQ�x�X�����l�@�1��]D D�����rh���E@�_謽��W3�$^�S��u���"�����6�) �>���3�+�L&˼���=��@�V�L�@�`�&6+ �����k�r	� �K��F��������ŖsG�b"���3X�åU�+M�F�k�|=}�8�^��9�/��<8�)DV�ǤL^���r��;y&��J�
A���q�V�LA9N�q�:�~g��s��?~��r��WWs{�.�u�ɿ�!Y�R�eN���W�o����"�R��aHwgPo��n��;�ZUU�5ɢx��t���n<_0���b��P���Y�5W�O^,I�'�qb�w���%@�"*��cda����q+���=�o<S�K��$Q�0s�G㲴�3�ODZ��\���\�#� ޱ�b���7�a؈Xb�V��pZƎ�;��x�2癐���\?�����&�H br٢�`*3|���ȴR��ؕ���ٕ&���Zi����{�<>E��6ӥAP��윣n�����]
F���������i��XAz�����GM�]�5�x�������h�Z)��Ib� �o�2"���7I�ѱh �����#�K����+u�i�?��U��ɽ	N�b#0�7��j��|Y�HF��
�7�4���c"ʀ;��1u�hS�Z��{t
ߑ�ח'���k0+T��!��Mj�_m��	�@17w.9� �ܜoc��e�@VD�,ez�}�x||�&�U����-O׶�R�l92jt��M���C�(�B��t�q9����F���,��'��T��A���T|�p�8m��(@((������DX�f{��@���y�ϋ����hɇ��
LA8�x���̑�E���\>mK�#�-�J���$�e<��
m#�ܫ�]Ɖ�#GV<N�/o�T��R��-!���S����<�fꪵ��uL�n�)����C��|��@  8c$cW�����;�%1�B�/��|��??uվ�w��3���iU谗4V\���5�j�h�ՉH��,V؟���qrp��JQ���]��9����Z���,���S{����T�^[**.��Y[��SQB��S��ӕ�]:���l�ce>��wtX+x�=��z����xT���PL{�X���^��m����E��4�a�6��0��>p�Hۦj���!3\�**<f���V��}�	u�X��*�/L	-��pKѦ���������  a��d��P��ߒ�?��Ճ�C��9����i�h��������Yuߕ��N�u�ߏ�#c2�����a;Ʀn��m�:"���8e����l/�=��\C�"	�D%(ZJ6�=�;5_pڑ�����P�Z�&�(-EB��T����鹮�-z��ބ7�;j���X����P���۲j46G7�����EI�S%�;ܡ1q|t+���Vm*,�����cz��&�����qG� �����]Qc)D:]�+���Z���쭗�Q����8;�L̉������Z�t�#�<%�0��L&5�F�����8��N��+�s���Z���US`���@V<dm�e n�'�tj7�p���C2�,��AL�Zccq(���0W`�% ��H�k�A�'�c���w,���ay�	d����Te!���
�
���>�$�]�q��y���)�R;�r���{3��k/:uԫg�f�(���޺��=�W)�#�`�0G��~���6���S���u��PG�1��������1������s�̀ �KAIuպ�AE�.��B�/!X	�F�۫��r��UN�_^�d�t���;�Zo�������"���� ���z�.����%=J�צ˟l��-�>�k��)d��V���*?�<u䯁���:x2��"���2?������%9����迪���)�F��� 7)/2��S�����x���{�椀��N�lB{H���:䲼8�[!Q����?RB���QVWkbo�	zb������Wg]约;l��{t	�M��%���G��لt�\����U�c��&����>��Ѷj�~��zE,G7e1S�0������
���;�nܴ�ʔI�1�Ê8i�40BT�\���-W�53?�����S�=�+͈��;8�_���k?�s�AOOEΔ�9">� ����U8Utq��: �� �0��Z��2aT�ѠAS�`�@�Z+h�Ƨ
QL]�PM�.�V���YR	�6-X�`N<�d	���bґ^����!*�Z�D4��?8�e���%l�J�Ά������*�����ٍd���u��ܞx���/�:ꉉ�n�B_EA) ��Բakaɾ���t��5�]���  e�N�Z�k�(��ͫO�JVZ���S�T��9o���qL�֯&Ȑ�f�*e[Z��)(�">�s��T�p�ﲸ�ʹ�0��e�㉯���+����'�f��6���@3?��ѧ�>ם��^l՞���B���AwkU}����;6��N��G��,q@�(ݼy�H�#ȉ�@IveoqD�A�[�`-wBT��MA�XFȥ�B�G�ЁۗdGذq������0l'=*^��C�=օ���u]�n�5A͑{4���\�\����[8ׂzIv��]yI��]W^wx��������_���$�\>���k�/O��U����������>�p�@�@�z�4�n�zs�邂E���Xb���ǎ��^ݕ�$��ߣ�G_�lr��������xx�x������vj}@�O�8�}B3�Ǆ�I�ӆ�����Q,4��H
s��T�lj�% y$\���tD��v�:^,$0	�O��Mo�
�v����Z�Kr3T*Dgs��LT$!�\@�X?��s3�r��ίy������:s!��j%=.��W`��X.�/t��9#�3��ד�7��~����Y�ܸ�W7[�ab�ؖ�c�����N�8̘�F���qU�ɍa�է,JjUx�o�,�v�c���������φ���w�^�(s*nI�~m�[=�L�T��(1��	����^\�.S�y-CM#�T��Á�t����B{L��f������ �����Q����QNP̅�����	z�Й���v���t'u
�`6�ӘEQ�`���f(�ˆ�d}�����I֨Xd�5G�Zۜqc4䈠k�Н�CM�D����0@�D��a
*��&PܡTu�{)���۔������`����cf���7�0�/����|��x>��q}?9��)��I�瓔N�]�X'LK���QU\r�6�`v0���.x.;������D�?�l�y�<m�P��N��(r�6`Qs�̸:�F Q���8�'-[�4��]��_�p��0�x{���S�R^o� |�WޘeLg@��(�A��CkYYFm��p,Z��㱠�d��.Z͠a�Q�OV�Lٴ��x���Y��ލ�+�'�������3$j�C���/~���xĎR�Q�4�Χ�U��a4s03����+�����EO8�z2M�����"����
	���}"��nç��Bo��=s�q�\�H���R�X�`[}<�u�C<7�8��(:�8��໱���y�Og9�{;�t��}�8�<;x��ϳ�!�x����8Hs�(|K�1�1Ē	E9�EB���i�\����uڊ��s��. �9� ���������7\(U��z�n�z����f�ev��?3�T�I�0Q���O�96�S�N�E�©�\�w}򨇤 �x������<�(;�+���ŏ�"�x���'�ę�ۇU���S]%�(*F_1�áIi����ʿ�z[�; �9k����_fz�C�7�B��\��pa+�����4�Ku�J	<������wm�S��GQ5~TV����~O� �g�w�ש,ܐ�ݘ����Y�r ��d���������[�)��O�	�扚�戫@��x+�&����Yj�!
I��]�+��*�Dk�>7y�upX3���@Ts��C�E�:8��@}������0�~r����!����RC�`�8����YB���N�i��쓓��mahlK��+m=�=���Q�X @$܁��:�W��LS��5�{'�b��FTU�qq���, ܚ{e3�� �[޵����i,ݴOѳ�"�)���(��)boNɊ+}�����^�{�'��F���G���"�"4I��@W
^�^�0���v041�'E��z����4�R,^��}L t����J,�z�}ί���E!��d�G�_YhHC?F�_�7�����}����*�׀0:7��]��&�m�Zp�& �`#�
�4I��̕)y�L�����p�T���M�_�yP\�c�����/z����E����~�Ӎr���i�dW⟳:۹Cͷ�d��Z�u���}�m4�����4�&׻�w��ޞ��]���c�sj(�8TTh*J����"uIg{f9�hl�AP9��R�go��jb�j��-*x�zN½{�������Cp'��׷i�7�(�NE@͞�����jK:��l�졖.��~�`9�i�	�f�B"x���ZY����&t[��*T�w�:�p��A|M�z��Ӻ�W�m�_T���;P� ��D�c���x��_���xW����sy4��q
�?t�1��H�qՅ����j���W��NX��Pd����V� K�&�p| "9����5�{m�����9N���񞶵����N����zv`Z���E�"���+p��5<���P��χ�U0z6褲ҞIA���E@vBt^�ZLP
�L�!�mR��X[]{wҽ3M���y��X�p۽=1y#c�$G�D㘀��";����Bۏ��G/Л^%��?����M_K���eJ�Ё2�}~f���_��r}�v*3��l|��q6����[����D��6�}՘S�[��_�����u�+q��Ң$�/��oF~[k҅��	O��l>kR�5��c#hK�V09kM?�O�"c

�"�&�Ò��#s!�큓\^�Fo����O�6de�6��9y#��)��ٛ	k88��v���t~�����,O�����b4�~���UHI�v6�1����B�)��V�44���{^]5�AJ�뽺z��
��$���=�ƒڍk�%���͟
��B��w?$ڢ��9b�.�}�Pۢb^h����l���ݭԞ͈����7eX�f��w�0zO�u�����sL�1����)��r5똕+� ���k@���s���
Y�X�,�dg��W��v`3���BH�OAΥf��׼��_/oEF��f"�j�F4韄*���E�Y9|�ڵ��8��B�M �<i�=�����F�7)ۮ�Ο�f\������rv=�H�qg$"|��
��WD����Ƅf{�$%� M��-��!�rD[5+�hi�_E_y���nR�|9�𦟋�eH�	��"`3v���X�8��h��bQl6��!ec���O���EZ��׋{1LqQ���y}E7�{����F��]|-9M9����>쵺�#��^<�
\?ã칞�O5��#�-S�ݷ��!�R�#bQ�4�Uk����cQ�e�3�`���uS�4Ѭ��Ȁ=F1�>�
ha�� ����e�Gɸc~TM��BO3��FK���f>u��/֪��9��96J����D���a���?`������z��S��Yl�:}�!��	̦���B�'��|W�W!K ��J��̕�O��p�#������uw�U{^۬�:�k�λ��e�*�z!po����!�][�������q �G/p�@��~y�&�5��$O��آ D�J�ٷd�Λ�iec63WgW��1�ٿςO>o���J����N'^
Kw"�g��a�`Y����qXЂ%�my���MX��1�X�*�U+|	uK����#�Sy�h����JyW^���w��#;�v��[�4�����u>wg�^�(/�:r�z��)���,ά��;�����>�Xo*i�v�e���� f^TV(�̄��g&�U��6��c͞�T�,�̰.�S��H���kSȭ:~�'Y����|y9OW=��;gN%G_��æ��yv/tW���k&!|��U,�d|Oϸ���@�1���qi����`��P�<���R�J)��������\b���-��q�u��ey��~c������隍�:�~TD��=�����w���o�wT���k��籾�[Ϛ�e2+hw`W��wT���V��@q����
9��/�?��ݕS�>���at���O�\P�ټ=�7{�#D�7h����W��\�M��lo�Q��M�Ty:��O�XIȁ���gH����(X-0�8������� ���2�#E����
í^"%�����Ϗ"L1�_��˪^��%e��2�%%+�/&�t�L�D*��Q{';\p�s����f�fi�
L@fc#��$G_sf�c)Ph;[�ƌsA��u�@���GֽS��.�Q`V�?�e������_��V-၎"�6t^  �?`�����Te���,�X��)��u�m��&̗$s~�������bs�J%\W��*l���� ��Ӿ��C}�e��g�꨷J�'�����ܰӧ�!-H�ֹVtZ�c?����ʶ�G� A��8N����EВ�삀�����YN�=̼Ūj.}��90��\�(�
�UUCi��x�͓N�B�3���QhЌ�ۜ��^��H<��� �^n�������[I"7,5-k+�x����]�G^���U���d�������Ό@�|�F6�����S��G�ú��ܒʖ^�@D�Կ��˵�y7��^����D��q�ndSa��^�*��@`�Ї�D���
ݥĔp ���elսd�*&�>�@b7�U�t���% �t輸��@��<�h'a}��,��W 8�VZ^`�:�Д==�֫�t�������N~V����B���HB5��`�
�r&J*`Ë��@��B�Ɲ���l����v���b�n���i���Ӿ����ݓ��W�*�a�o\v�B��?T2����C���㰙��>tq�eS�����I�I8��q���]�+q�D�ƫ�l�������#�|m��y�0��g�Og	�FF����+��:��Tn���ӈ��Ϗ�F��4�nx���H��UWQ����{�d�U2Hx }�P��0^��oHa!U�bD5���,^T�A����/��ꌩ9�!��J����A���R�LZ�pʙ�s��p��j��Y�+E���^}�ՠ�x���U���Ն��)L��˭�����߂��қ����Fb�8>;:#V�&�
k�������0
���֞Η(����oh��J��~  	??��	�U���i��'�31����&�������W���JC�?�*������F�私��]���U���ve�%\�CP@&)m�!#�VO�~�z���XF�i&�S�m�h�O��J\'$��V��SYd�иˎd�0$�$y�#�^� �9�h~TC�-3��JY�}$%y�xL�F1���Ԭ�+���z�0է*��A�|�u�]��{{+�2���Xi�Xi��Ӽ��l-.��I1�"dȿ�f_�~b���@���E���N`leeeٌ�Au,x�3</�)�:�u�?5�=~��r[�[(YX^6ʥ+X����t�ktiF� ��$�ea�G^	P�_�1�\M`�럘u��7�PH4��Q]��1����!܆d,I��bٔ�樝8��e=�tD~��_��K�S�'�i����h�z�����*�����6�
��Q��?���ZE|��_zA`(�R{�L�ˍ�`Ħ����d�J���k��>'B�g	�����T��f�\���J&]�qT~'}�Fc�b.�Zqe�qF��o,�I��A:��c�r>[�y0WM��f >��L_C���m�z0͗lG���.�3�Õ����>����{i��7��Y�sEfmv ��R�qw,��ܱ��"��1A�>&V�3��Q��o��JF��}��;-~�J�EL<�-�Y�>�lhM.U�G�3j�<M�b/����x����a��R� ��U��H���V*!�y�'n_'/�9J�|��s	��h���)]���gN�Q�x�?~=Lh6v@�$��k8�ý}Y.�	FZ��u�;朧2��q�$��MG����a|� |0��������i�����QW�l��ѥ��/�uK.]0Ckeo0v)\}#��tV�X!ln�׭�4E�ii 	�_��c�=;Q�l��nG?O.96G��CT��r��)��&%ꚑ<��d��$���s�Q0ɋ��D���I�n]�=H�����|��E}��|١L���>~�p�$V�s'$E�d�?.)j��P�O�^.)< ���� G���S�_QD\ϡ�399a��<|@�<�-�U�"�|.=�7i��r8����KO���N���˩;T���?��\���4h�+[������T*�Gv���8��Z.����c*}�^��V��Չ�Y���J@�:=pz�ҌυAWm��d�y��v0v�׌��U�ʣ n���V(���^N��ѥm���7�2����_u���%>{�n��Mn��v'����S�����o���t8�4I�Y#�i�b�E��Ƴ��%��a�'�N&�V����h#��l�y��E������D~?Vlr}5��@�$�6?ٿM���ie�&H2�R���H�tv~Nl5x����Br����$>תCA��(��=+���p����t�A�^s<�*�ޛ�U]�?Y���`�RI'#���d�l��� ��şY��.~t�w׫�Z{��9��LɸG�Z|�h	��̒���:0>d�PR����[f���k�kY�]�g�M?OG����pR�������:��(�v�,'J1>-1U=澹�x�[4���D��j�e Bk�=� ?U�6uɰh������@Lx��IC��	F��{��A<<������\�Yyz��:��ߔ�����x}�#U|A�_B�ra�
"6~T��.3��V��#�'皧f���A�������]JN�A�}����C��TY�n�g`6VZ�}�]��7#-9:gα��.,���e���9�,�a>Sd�S";� y���b7��wC_�8a4?=��ѯ��嗻e�<�?��}*[Nm�zv�z��dbҲo��&���C�Qx�I�w#H�����4c�v�w�s�)�R>pV�G�c�%rf��8j�P��p����31UJ^�ąF?�⿑8����e���P�!j,��C�e^|�`���IF�8��ޮخ�_��	����g 7�y��a�4�^��:��]%�>��)p�G4*�&]�����}3�����隷V��i�;�1�d'ǩ��=T=���7	P�/6��Ƞ�9�p3G���2v^%��Z��T(I�S~ǳ��x=�8qpR��w��:��D�����I���'��ù�g�[�y�~��F�}3��Vg�#��T� r��� �ƎW�d���]s著K����<+I~�W+b�)���[�"0��޶�������I՞㞾yο�����4L�w����ῢ�+�!�x��5�����V������Sé�\ixv��`��)��{��a����VCT�A�~���E]5�N8ha�z/r�,�J��h��T#�_�Rb��8/iF��_�#�WO���Xt�k�Q� x Q�O-�u6����"U��g���G�Y6[�w���C��u�����]������6�u��n��qwlQ9��WԊ�'�>1"qE8�G ����.@��4r$&,�@hK���1�6u��~8J���`on��~|I;��E��O��[s?M]{ˑ5�I]=����4@��y������\߫q���/�<����f���솆.x*?/���"ofM�K�`��lK9�Uu�֤�����B^v蒓 ���}�����A�QۧI�x"�_���7*e�i�Nd��������q�3�%�a!��y�s+�um"YSUx��Y�D)��ʉN�c����а=q�f�閭�������$����U����ʙ����`"��V���!�a���mS��G�ElB�%�k��%y���+��2RK1��p����e旯r�]�=p�ߠM~��w�U����)��Uџ{O�\��%�V����n��� ��{�������@����FJ �a���Dv|_3�ƙB�R�(4`T�E�n�DR@���`l��\V��&O�dk|Ǣ���Cei�e�T�)�	l��	��j��v�{�_|�����%2Cױ�(S;qD�Q��R�@�G�O��wA�g���:
Q�O�����.��?����G�<yZu�{q>^���P�1�"�U� A���z	<��w�w"��LĺU��_Ơ�`rj��Z *!�eDd4�!��g-���S�nu�����!`U�sg��qp�x�o����z�rh��?�>�(�>��*�G?�����K(�S���0�eBN�X�!#����8��c�߱_���5v ���w�~�+�>��I+�"��j!�Ћf�'��,CCA���>��b�t��jq�Yr��S�C��+͚C���o����0`��9y�ձ��Kϧ_�Wc���cr]>���	of�G6'��w'/�QC�Gn_N�Y����8�QrQu�%��2*|F��e�'g���̸�
$��h턀/�Q�h�=�1wՖi��(�둕��˦ך�y�᧛t�U��l����4�wt6.S����Y�qW�2��ȟh�,j[`�!�7T��*����^О�yj�d�̲ �J�W��5�k�ś�����Œ=B��;6���<Ϟ`ء��
���A�v.*!�$_rڄ����Y�Ɵ���u]���/����f5%�\��-HU�]:ǥ};~Ĺ/^�m��Sވ9�}F�����ӷM$��%�x����J�Up?�?�w�8�g�+p�ȯ%��9m���);P{Z�	�JG��AL��E)4�!��K���Ο%��ث��C�c�9�| hNe�x`�h�Yu���7ܟ&>��be$��΃��i�;����¤��l�J++|gji��i<�����M�i5��q�k��S�7�XRm �`��l��';���"��65��]��p���N��=���	D.���'hrc����K(���`,hp�-�5��I��'�ضQ�
U:\��O�e^h��Nɟu����aV�%b�&�����ӕ�}d?v!u2mk�hoo/h촐�����Q��xp��P�Ԭ���VҖ��k�e5̝�(X³ǡ��ѥ��~R?Q�"���L�O�"��⤿���\��<�GW�l������5Uw�UiG��R���8���՝�](�37��u3���$ǿw���w���]��+IWTr�;������jj�v�|�)X��7����1�֤�\
������ӊ����d�&9E�]�{>�\��I m#M�?C�<gz�;Er!�X�����:��i&Z@]܆�A舞�����?&�����D�d�:"�`5���3�AQ ҵo`�f����s{��	�R��v�����k�tOb%Ӎ0��3�el�h�¨��l6��>��*�(�PS�����&�QP&U>DVA�nd��Q9��@��e�q��P�j�v�U[3��?cէ�D�Zm���ǗG&p�"C��[R�2p	�t��\@v$@���$�O��m���� ���xx����%z1"�ٷ��d1S�z>-f������	�Q�(�$q���cc��`m��{��� ѻL׃ܯ�9��uUN�7��oȚ�L�Yf4��]d �F�dm�������(]g�(vb����<D�I
Ll��h�����,��A=��U�b�Ra�He��?����L�<�QT�.GY���W@�{9�]�Y=��e�oF�~{���i�鿲m��*�����h0}Fh��2�-P6�-��|y��%I=f�ă��QR�ui�%&߾�c@������/����1���2����=�AO�����qWI�Ȧm�%6^9�O��r~&&���}�]z��0���j��}S<$�/�h�(�� & >�ƅ�����bW�7+PMb@]^�WΖ��>�۔�d�V�;8�X*�ӡȘ+v��:�5�#<�o�x�����6��H�j'r���U�Et���;������APr)�nX)Ab)	A�ei$�qD�%�Ni���}}������fΜ�9�9gf�y\Ek�9�(�j	j��:�������Qf�}��|W�6�"6nΗ<�.�E���9�W54��ƭ����U	FK)KN���Bo���`�8h����d�Vl^)�8w���o���'p%�ؚY �M"���i�׭߷LjM�;������+�Ob����nc��H;�/.�$���GC?7츞�L,�m��}��S�W fK�5�&�Vw&�'��bK��`��"�� �'���2��XoJ5��h��q#q(�����Z�C��﷾X�k�Ct�o����\㼘_=_���0Ȝ�N�l�z6B^�l��{x�O�ठt���W��"rq�ĎϷ�*�!]UU;-gx�݆�`)�@��(�D(�U��$^|�*��͙����}K��B�վ���K w��βg��6HL��3��j��fn��r�|8���K��/G�HD�Q��x�VM���Іh�=���(o����p�>��H$#`,�r�H�Z2��8��2���hD*�q��Mbzln�Y
z���C��f���A���g�ò+�rin��,��)�`�n���_�T-r�<���V�Ŭ�;����+�͜�4��xll�D炂�S3�F
4��5�l��BB�ܛ��#|<C��������\7�P��y��#������� �l�y!\���`�����:�d^qs�y?��|�����R��a>FJ�pϫ�_���L�W��RG��bM0 �e�6��άĥ01>�`3�PرP{~ �]2�^W&Vp������8�r-G#����tO:��ؗ˛[9$)��].K��ż�v�P���PkZ�0�,�6(�Vy���6b0�=Ъ�Q��3clj]�p9U{�
����e/3��|���#u�����A7����:5�_���*�ڛ>S�3[~Z��?i�-}�P4mN�+�ͭ��%�V�ZT���������� �^�T�,c���7F���*��z��ej����M�����o�����f���	�G�/b�k���p
B�fK���DNX�V��2�����mf������d��(�I�H���2:�`�)�S���g��.7`�_v��;e��!�߲��>V	���\�v�ש*�I|�znR�B��g�;�4�,�1o��&�T���pU���������Dd~���r=��$�z�}d!��|Fw��R�W��k?8��os�� *��3�{���-O�A���u<M�r,-?���)����Y���-����;�`B���^Y�l�R��M�B�9���l��l�&h�k��x'������Ň�Z)�:h�{7?��_}]Q��R�����G$�]>�XǸ�ňˀ
� 17�1�|���P"�"��cji$��0ꂬ�cd��%	��zqa6�l�}�@���ZM�����؁P[xa0����-���Y��* �ƣ��h��6����Հ�܈�����ɶ����2]�zn�����JQ�TJ
	y$J��N[�OEa��֤��U��*H��;S*5W�����QT�Q��w��vj.tqڣϊ
�$��# t�;��$�(t�����e^�	S?_g��)u��6ܶ3h�.�j�~�ձ(@�G�W���M��~��r��`	1��X����AZOb��7r�>��)�w��]�N�,�iT��`�E+�fT�V��1�p�������|c���חǨR��;k�-�4w	:��� �[e���F=�����f�y�]�a*�Y��u�T]���FgN�笚E��h�&dҟ�.�;���h���~d<s�|!�� T�S�5�u�Ib�	�Ó�l�^� ���g�3��i1=%�;]�w�B2y��0�m��h�y1����_��*|��@F�o�rɭ~R�K&E�n�LZ�=�m�6����v@l��}��ZS���4���~wP��wN.泷w=�=��f o�����`��H����k4*	Fb>& O�o6
y���O��w5�
42��K5����͉���� Q/:llETE�PK�ţ� ��Ӹ���అ�iSu9Cu�q8p��wwֲ%;�S�t��杍�+�Ώ��ҙ�:`z�X����N�ԇQ�j�֪�� �]Nn�QxP��}���ܰqR�}N��/�>��k���b���i���������Yk�	�g�����w��ᕕy८��f�!���ϟ}t9)Zg�v���5���O��
�%;$ؽug���9����x�	f�𮱰�k+�pH���w�J ��ܞ��zհz�b��֦������o�t�=�mU���*���fs7j�Zm�0?��!��)Sʹ�f�V�57�E��-u���375U�B19�>��!56iM�x��8�*D���T<2x�A���O�	���Ȋtn��T� �#���S獍J�H��ܫH�;��4���c�a5x���$©�[_	�+	��0Z [��d��St�~_�59@�ȫ_r�Uv��'M�8>f�ȿ�H�J6ڟE�".0iY��&�"V�J���nR���	I?:H	<�B��v�hnNU��ii*ɡ�e<��?1;���pQ� *����fi:}��9���GWW������و��}��K��w�g�&?�_˸�w��5&�</U}�6�C'��Ic#������\��ε����l�
�|��!����b���F�W�e MƼ�/!((�0Q�ϱ��o�]:�k����:�3KϯJ|����dl���3��n��N ����9�_�T)P_c�p�IN5�ˣmZ$�o��M�l`��N�;��.���B���62��w��nt����b����Rhq>&  �C@e�c:��utt6�3WD��k10�\�'���
C������??j`�)"�ޛ����r)隃W!���|<>�љߣ��u#�_{Za�q@,��V�#�'�&�~�[��ϓ!1�q�9��$�P��Ҩ3@��3S��^���45�aI䡠�&MZ�Y������[&CB���:<�^ݯK��U�Nvu-�+̝��a���qQ?��􇖚�\v�x�m�i�"�w�8�Ƿ�ʾkeڏ��j��W�{�*��idK�P
�T�)8��[07R�t�=b�Lޛ��n?ƕ�N����WYTd��/�|sT�NӁ�	p���y�z��"�Wt�cPֱ�<=�����*
+�$��_r��e��;a$bz��)��P�f^+I�]��[��
�����խ��ߡ!�[�iesS9H�a'�*��m�c'dK��P!�S�3�4��O;ǌ����.b`$�����!lV�X����[C
�	�iC�Ʋ`�6s�1��S|����G(!!�!�9�¬$O0�B�-�������5�M�z�;e�����6���IH���Wv^�Y�w\�[Ӫ�*-<c�F|&Er\`u�:\��=|�VW\lwH��������nJ^�Ӆ��\���w�S2P����+k�l�@�Xvc��H�I��{�d����'ϰ�oHt�G�S��~�l���U;�Mq��uq�3#�3�?�lmzJ�Q$v�ִ���X�l��?�H `�����h~�s�+C3�uȟ�kS���?x�?Im��Ō|߮�����;����!��Ti>Is_92>�ό�E��1��4%���k1�rB��%��ԙT&c�D��uǖDKk����~��pm�[�k�\f`N'@�o(�#8���8|�x�BlHq�^�Zn�eT��dڸ�G7�XS=b�{r�?��T��ӈur4��}2�
��[���?��uB�!��)���|�r�-Q���:]���͈��0m!ܖbx!a����� �?���	j}i���p�E�wR����~!NqKj
��'�M)3��*ϫ����AวJʐw�R�p/q��c�A?]́�����.�0�w��]4Ќ���dE�En�J��O���]8%y]]�'-8�4u_ma��~t�����5p��~f� m��s��!@jS�h-�o��z�����߫���ǴL]w�ԴOp�z�܂h_�/����G�����tz�;��٪�_3���d��Ɉ�i
-��N��P�3F \���9���t.▖�0}pZxv�.-Q��j^նw�������R���t *����s�C�]xD"�qI�[(����l��"�aM���F�,h�>U��4�BG��q�Zt��T�Ӵ7�����>���UGi�;DV�j�,Y�#�:�ҝ����FFFA��_k"x� tw��n���;�������x�9$��\Û�������ƨ� ������#��ŽNv�����׵��^��W������*�h�hrFD�E�ǅS�ק{kAF���At��rH��,:������F�N@�2�{�[ȳ��ၚ���Zw�&7���b���϶��Ob: �{D�� ��4~���L�O�5:�;L<����,�h<����?�Zh�b=9`�?�9�X>�m����  {���?�C@h���l��O���$�K���=�kR�?]P��m��PK   ���W|�߮�  ��  /   images/61b75eda-77d0-43e1-8746-2b678f56ccab.png���[�A�=�J�R��PJK[�8w(w��.Žh)��V��w^,��<���x??��5��Z���׬�{�?*I��R�b``���H�b`<����=�]`���EUZ�l�z�!+)��i�����T��ҭ�v�q��8�@}r���h��a
k������?�'�KG�
' ����"��N��[�m�<?:Һ̼)�r+�oß����Y:Z�3�\y�����
�A   �I�Z���� ���A�@ �z��VK�w������y҃A�xu�l��� R��'���o2",�� Ab!�����ygų�oA �)�!ZУu,=��5x��/��Q�'�������_����p�-���Z��?�ѣ� n&����������s��9��������i����؃����~����=�9M	��� '	n.[�E��չ
�c�g�j�-X�[<,M.�����ɓ4��O��^n��WR%���BB�9�o1R�-y0*T?��U���$Ae��sT[	ޑm:봥lI�o��d�ll��=�]��T^)�T�[7�	sn
��B��uH�8�G���>A��9r�N��>�G�]� Xwа(�
@mo���sW���tvϮ�&�#�����������IƩUF����b�6��GR��Yd�=�#zc�^�ş�����A`�\չ�����ڜ#b�?�l��{�1{�w�2�џ����z��2�X�uk0�x��Q�9��Ər,����%U$7����τY��I{O^s���eK �"[��%�YQzѭ�eȮ����Eo� �WQ̭����>�2�"�����?5�8��os�M�C����I�FICt��U<[��)7z��O��[��
�<��	�2T��;���I�*�:�Rs6~if�'\4���l��JԾ�nS�@�W"΍��CJ�)��֠��1���������竞!6�6�Տ�G�<C##���F��������N��(P�ss:>�Q�:G�����T@���q>���+�#���*�+KIr�߉>�xòx��������233�}d�e Ir���a�I�*$�3{Sŗ/hi���9��q�Sp���Ip����l	��扇d��G�|%q4辍Z��/�;�$�8mW���%}̙�����哑����6����е�/���"c�=���FLE��@cDR���In�,.�\-Y��$C���1]���:?�����l�?}Fr���6�m:���W~=�����a��T�p���Oj\��*@@���XM�_u�o�Z�r���%$�H��)K�t�D�gԥ���N_�ffR}\����q���L1�n�cr�N%}~qa��k�+@��ӝ��>�����s}�����9��ri��*��*���"p��4!���Xw�&����#��<1���2�x�ގ�wo;jw�~4�C�����M=Պ��
�������pt�����/u�g���5�6��.�,�����<|ó�]��FH������3�k����Su4��:'���!�<���PjY{��t�����Lzn����C�֞S�t����R�g�Z^w��Ь��f+٣V	�J�_��;���m�~�ݩ�Y�]����q�rss�v0��@AC�dlii�.�0����=��((6�.�"'��6���#�D�c���iq�3���̶m��c���̎�]�+�R7\�q�Y�f{�`�>;o�}Ȟ��7�e�:�A����Z�ˀ��𮱱1�M�kf�0�\�Y7���Xs*�jG;o�����Ų��yc
��ΐ!��~�+
ZuQ����:����M?�n�E׬���y+4ica�1`Z���t>��.�*����lnn_Y��АcF��.%��6js0��,�\K���@%�P
��5��� �At�6İ�V;M���򡫼j��zz>���_������45�L(�\{D�\�L��������|Q[ۧ"�$����0���V���k>��:��d=6�%8��e�[�M�H��������������i͂F��͓4ԛ�Y�r�t��Š��)ԭ��^���Ԩ��v��f�|h����~�"o@���󴗷�?^�XQ���d�����q�0���]�6bv~���D��n5�r�r�`y���Va�H��^���m^#�a����ݿk�d��`A9���ō\��`0�vw��_KkFB���0�qrr��Y�}����a�Xh�X�n�R���]8�s6`�֦����$�38b>�ŸSf��p.<�+L�s�\廬�<a玕@�`�3E�")�����/���N��\"���B&N/��.5�	q�T!o�E]�3��X�l�Ӳ=��
��Q�Ue�Jbe5��\���ăo��>۔s�w���o�(�7�'��Q)x�h׭Fj�쏶��"��n�O>�gh``�ѿ��.3h^�g����7q��m�E��v�ۧ�Z����U@�N�b�\����N��j4�4f`%旊hϏ�f�qm�p����MUC�\7,
qc��9G�^�t��K�l�K��n_�D�`~,6�&;<<�4�[�]�D��J�)�ݽ��t�9�G����dxˡ��8e�Ы�s�Ѯ��⫞�y�SR �|I	�iK�������C�ݵ�����N��v��?����G���k�=|~S�-��PU�<���7�x���c�*�1��]�R��CƖ�y:$�������.F>�
���=^�&����WY@>eT�>#d8�J�~>�a�����`d%������S�X���W&߬w�$��'zh������U���P`��x����0���@)Azղp赏r�/ �WA�P�Dc��(�VU��N��s��Tԯ5��G��H1�vˣ�h���FCA''��O�j�g��D�L��2��=l;r������E��>�Q��`�QwA���n�N�sc�2�X�I�XE Ɯc���u�3j����Z��}~A+�3L��f�� _���Q��f�d�Ip�~�wS(�yZ`
���dk�!	;"��;��e�s �B0NW�H;qiÄ�i��_;q�-OM�:�����bEo��,0�G/?U�����$�qX3q)��Y\jZ��s��UlqAH�Z,�dg����U�W���G�[��y�@n��s� �z�4�ߋ�yA��	Qn�Kmߦ�\��E�dOPڑ���9Ց->5���*���H���Lw�o�ͩ�G���	-�u�����[R�׶��?��~}����v�oo��Z��HR+���OdT�b6hZ+�gbn�����1��y�����?��x0":XPM�R���.��X��gd��8q�Hh۱��6Z�Do�|~޽E���n�ۏi.�5ݼ���L=��cߥ�vt2�=��3C7��x��؃j��Co��=�gԀ@��^�E�5y�f��t7����ׅC�M��F�HW_���]
����}8!�s�E��A�T�ʩ��^.�L�޺Ί`�Oa�w"��6>xR�4u�BSS�����`��SӨ�%���6y7=��������a/�ҏ��}�S��k6xů�eЇpX~Z��mÒ/rܟZ9�d|OP��[+O�r8�]��%�1��x?��6.{����L��>�`�djTB�-Ź��VS��;���e�kwPIh��ӭ���0|~�$ܟO�(A�ɫ�����ʧj�ie��rH�����<�E���m�g=/��F�>w2��s�\��J�0�j:ٮ�}n�}ۦ\���Ű����㲔u�v��\�:���q�W� ���P�P���-B��Mk�̯!������^����ƻ���e�h�"α'���&G�A.ॐ�������|�Ժ����XF��J�����A4>�����ĳߵE�,�I������t,K$�5_J��]��q�'���]hA���?5W�sO{�ǥT6�с����L�Mr�����H'��_R/T7T���˼�}C��m<�rU�u������[�(�*BJ����Ί����{:m4�ڮS��4�n��*AJ�W��jǵ�ǯٖiʏ�m<�}I��32���e����d]d!m��� ��	�
IYD�9�kyH�}J�&�	�� �Q��X�\`�}G�ū]��Z�m����H&əU�f��B���ڻ�A���H���Lt_�y�4��YK�_O���J@�FH5.jIf�8A���,�ԝ��pg� ǩ���r��pkW���A�EN��gFGF��N�a>�ǃ_�F$en��|#���$L���w�Hܜ������Q�X����A<���M����4L%>7�{:�S���; �(:�2XY�6ڋ�	�"�%t3���U�@Rx�}z#NN��v��&��v�Q��#��|��i�|ꠊм?��ط���b���"�E� �?��	�{���D����u��Ǣ,|>Y������ο��+N��n���R�by��N�:�fd���QqZ]�'D��:���|�j�j��r�v��n1�栚�o�s?1@`��}���_g��h��x�E��O���|y���[�3��%���#�d �{Ԡ����7˭�fw��k6�ALb��'������qptӗ�yC�R�tP����[�9j@h�"x�Ǎ���-q�ȸ�g����!�I��M�Z�����F�O�I�X�D]���*��o�Q���%��~�!=�����.z��;�ނW2�*�/ݬ|Q�����d�X��cGb�$,��V���Z�xX����4H���k��΍a��r��n��S�H�P���mg�>j`�yʝBPQ�����c�J�iUO������P>�zM�K(�}�W�&s7;;;�J�����|9W�?b���t�)�s?)��&���������ÃF�ې�ɛ4P@�� a���0/��&�
��j d��߿� ��߿�l���Wp�5���ɗׁF��ņeP�����B��,5泷3OW��o>8�;��
|E����G���|�9bva�[#'v�����*$����?E��[��)F�>�^	_X������I�����sՙ���r��C�e� p=ҥzW�ѡ���K�we7;_�-DM���e�\̊�%55�UD��*ق�a%���'-5Փ� S�[\��`i>1[��~�����=��=ɮ���3�ݓ��r��!�kƜ�I._J;z�CK��΢F�3a(�!��[M�C[y���5�����}����x�[��F-Rp_=+˅53�J}K��Q/.���J�Z���G�K�G1N� ������w��f������M�07b���Ց�$��0X�l�8o�b����z�O�t>����U�o��I�
��D��In'��4eZ�C(g��l#���Mvc���i�����_���s���i�t�7�,N�s��=	����ܗ;"���z�J_�Iʩ�EKG��n6���n��J�&Z��kyr�c	��:��K�����Jj$7���|�]�HY��w�:�S.6�]H��'���WF�}�i:S�Ԑ}3�IW���
�z��GT�t����-�W}���5xU��RrgfL.�W��E�,�i5a��XZ��TVV�~uK��!��t� E�٠�^���p��@�����=������8Yѫ���������ӳ���\�ዤf��v�z��!�f������������
I�j���&[.WհҤ�}�=
g���Ltċuyh��P-��u�x�QS���S�ɦY�T���hg��s�qQ�z�-��Vn6�]�:Z�]�t�$�#�J�N�M�٪:{=^�y��ŋ	t�����W!Q��dV�8oKKK�#� <<���U4���7ӠT�,bg*ֆ
�����q��8��N��~݋Jk�ܗ�{;�J����Y�۟��n��xmWv;�w�!E��v��K>qB؀�e�9�-���n<ZtF��&  ��q��Ï?scM�p��k��-���:�=W;���BO
"H��w\�X�I�g�]un)sY�?'(gʘ>E�� RsF����ޯH�k��ё蛈�Z�Օ�IhH��**���R�2�%\��3}oKςn���GY��Xm�<���ʊ��
Ү���3q��fB�nZ����@S�}�ǳo2L#%e�m��g�k��8A���������#����J����@�h������Q�j��,^|��+{�舯`�@��|o�2\dp:�Amex��u���8-�H1?Y�l�m:�W�u�J�������5�SD�;-ib��~��)Kb�kT���a�Ȏ�1�Kjkk��`�����K���@� zs�Q��|���� �dU7٬��2?�8�=x�C ��Oz����4-���S�V9�W?>��A=M�uF�u;&s��&�7�˱kB�����Ŧ{��W�8S��]��`§!#>\�����
5��ճ����ȧ���ۑI'�T=.�E���&�����븜GGR�$Ƶ�ޑ8�c_⥡����������`���I�o��)x����KyI�1oooyò-�$SPD2<�Z�I�v�Ot繳5�ޙ�t�~���6M���ͨ6����J�y�^ ;V=�?�2�
��a��P}ͨG��R��GV��^:�_��ָf.f����ɚe�𡝝�2�*�)����y�����Ac�0��Q��`r�OAF���Z�;�x�dr���z���Ҥ�&OH��#��/���t��Tw,����:��?�l\�Zxl����A�����m1<��d��Q����j. ቪ���[� ��!nC���}������$o��r�T=a�ÍR� �Xvr��mX����������t�"�3�V������ƞ��lD�v�۷�Z�K(/i���L?(.�d����'P��(�4.��s)?Z�
U�,�b9��+���2�7���C'�����;�Cd�?�P���9&�@c�=5 �6��a6��:p��fs�X��u�|
+��o��,^��m��8]b���6n�����	[�Sp�p�Ga�A��y��6�5"�U+3,x��a�t>�hmm��Q'b5��[�Ez;����{���W�.����p��XG|Th7�Ǫ��M�a�}:����h3kX�N�Z��c0o�?��D$C��X<RJ�5\�� �c��$���.�8�9o������5�).>��̤�VA�F�vRRR�����媲�/�PL��r:�62r����Nw@꾙�#-�</�7˫Y|�#�����v���]�:�՛+C�J-ЧU�G�qb�#>��s��S|�P���
�C�Xc;�4���RP�o��F����C;?�씄��`[Nc��p�'�oCK�)oe];�
4~E�_������r�/(n�ݵ~N��� 4;���xx�"�4����-�G����~,:��R�N�������P�ЩJ�&���f�tR}���Jc쯢��������v���Q�����'8�j����wʓ�(��7�1Ŷ��@~ �N�#k�����?6�������E���!�c򹝽^����A�D冭7�6�%�+?�u`Y}�"�sP�D��AQ�)��ďU���/��\1�ܐ�D&>1b5N��$� ��V_~�N��$�L�d7��=�����g^3�uŔ9�4hL	6�����$5J��:���4I*"���T
C��H_g�����<F��#Ge������aUEu'�aK[���ӽ�)�W�ĩ��w��|hx�«<�P�N��m�W�88�L��kfE+��}E���G�*$�a��A����{Ռ������Μ8L��{NE_\8k�)L+�|�O�q�G���U��0s�y����W]�V a^N��-�7��g��t7�.y����T�a��8*
	Ǹ���ĆQ�BF�]L�
��c��Ǝ��Z�LeX�%%M�����!s4�F���>��]y�ߜ�.��;G��ȱJ�CC��d�?
�3D��p�%4��ː!>����R6�(Ay��"`�ˋ���`�@	�Ib�������o�0�4VY�L�fy�B��T�}Y͹�d�h�}Z������e���������zZ�e�Tf�ȝ�f���R�J��q�f�-�[L�2�~l�W���ؼ�O��c�|�ͩ`'H�WQ���|����}�)"{Ĺ��@GN14J�@��%��+?_��y�'
7]�Ͳ1���zV-�<�θg�!`�8 � 3<�>�1~	�������v�H�H1Gl���z��M�8vӲJ�5�[aXx�-���_�'����N>=����/�q`�n�����&�}a�g� 9ϏnYW!��>h
 �R uލ��먵��X��Ax5���k�"�&��h��Oir�/]QD�T���s��3�&���'J�O��I�H;���-ʏ����,�;�#���q��đ��V%.�S�	'�ӣ�zP!��E˧�11V
�	��:V�8Z������%����c��hk����c��'>�U�~5 ����·a;xX3KcA(^�+����B��_�4��)��d�Ɔ�
R����B\��/걹���0!��ve_�W�Z�-����\��K��"@�c��������e��"E3��Y��'��w����Zd��	4��{���,�λ	����맾-Y�λ�_"�nN"oN�}D���+u���3M��T�A)�VlDɿC�Gi�KŲ��O�l����G�ׯ�d�'h��C�U����y����Q��~Jߏp���ʋb��i8%ɈplL�Ɋ���+�dd��?���5��	���R�݇?��}
e�[u �-&ˑ�T �qV��B�퉽 �W�=����/�����2����xDfĢ�8\��E5�����뇝����2~}U���;0q)�&}�n�xJ!�ٿ�<����RD��ΰ��R��,1h��Pm7UR�/��J0�|U80:d�f/��6g�EJ����.�#�^� r����,+����.N)�Fʾ�B[�ч�5oaX��/c�X��`�է�(~�-&�f�bbO�NVI�M���L��2��Y�8}@��Y�����Ã���FLd�|J�V�:�F���ޔ�Zg�+���kJ�2�by�k�[��\Նb�Y�|T������A��3z����"hỄ �v��p��@Ny�����y�@�h��ϟ�|�Ւ�1a](Fk���XjB�v�D���g��f�����:�]������/V�_)���_��I/S����\��_;�r��9ν���iO�
���+�:.*Y���Q�|AnJq�����8�O�a�)6�����4>^ê(ቆ)B�pFLdqb�E/��y��"��������L�\npΝ+�0p�ޙ�8��U�������������w�a��B+�J|�^��)�J)��Qƺ�<�w�=���$��/!m�Gaz��]F�;�ӗxU�I#>qS1 �h@����:��|/�p��1>�MԘ�� [��?�u{)��(�Q���{�-3,?>\F��#ɔ���E���-5RU�O�D/]����>~v��r�䰤������3�}�e̦�Ԉ��}s��h#�ǀ4�I��~?S^"��z[~��5�C�gK��+B��*#">���[jP 7.�Uص�s�_ ~c�q-?\�G�� ����� n�~m:��$�h<�V�e����'�b��^zz���j=��B�V��$=3����M\���P�%�ӯ��vM�=�y9��� ��n�e�Q��m;7΍-�e8A`l�{���~�7̈#і��n�^���C�p���C����'&��in�V����æ�lԮ��q���4M�W��'߆{�l�8�6�{b�x�^��Mܨ�,����O������v���)�}9�c�h��|�Rq|����͏|�m�*F�`��`0��g��P5^��fTuP'���8{��3�7�=��j�`8���7�cG���F�Ԥsv�.ڨ��%MeEf<)���U$U977�ɪ!Z���)~ǁ����L5�֍���r B��%n	m�+M^r����a��\�|�xb�f9?�iD�����AG��o�F����}Id�x3�#�~k��c�F�O)ۤ�������K����nn���^�[��E5QSc;�@�y������}F�|bL��J�gQ��e�QI�ڴ�|Z/��rY�MҎ1u�7'��·Ē�+����`^9���4�uMY����&�e��Ԗ���ѡ��3��<Aj��_�<qF�IG46�w���m��X"6U[�5�O�IK2E�|S��_��������I����B��6H�k�/�f��J�T���Y�Co1w�!Z����<�g����J���١(Pa�Y"��S~���ݛX"V?��>r��<5ΡDi����f��"}g�� <�jSmY�wC�E}>�W�w�3����R���Lˇ���'ߎ���F	���0>?��'�Y�4���S�������=fEg���'6�@tc��G�9#֬���X�9��
�1���`W�?���-O���Hp�JH�:�M��ksN��j�Q�_e��Ꝫ��e�f�`�o9tퟕ�[-/��x���u��8��*fZy(dd��mA(C--?�9.-���}�F�S}�\�"� +Խ�g�/w0����۳aq����|�8�����w{���΅�1�]�J;>3N�5�&�5��r��ZWt�J���\*��+L#Ag��H�@�c���Y�nC��B��]���N�W �}nqr�Ѯ�5:7�:����9��bĒ�_��eׂ��{�2j����)"��ȆX�������z��cp,��C�df�2�}���I.��l�󇰰����7���|��o��I���]��U{�"����v������;�w�oAo�>��)���Z�g�e�Ȕ�2^�ԋ�|�����[�B�ִja�T1�{���+B��Y�����D���e2�M�����������u�:pw�^1��y��ҠL# WV��F�xӣ}���p�e��ܱ+!��}�	k.��Ƕ�Ve�O
ĵ<f[��z��ۣ���gEj��W��ζ���<�cq�Sٸ�eϚ~��{��؛��y�IBz��g������rf�E�F]���ڲ�R̀�第"<�-�r���z�)�wfNQo�i��Bs���D*�|eN�)��Qx��5}A��\y�T{�-�y�$7���ef�l���߄��9T8���I���A� ��q����H�_^>$H�\�E�	��C���Q�&�f��n`áwi�V<���YHj��������և�+��WWg�2O�e��/4��Xp�K|'��5f�5��D�b���^���k؈�JTM��0t��z�$fG�^��Tm}���i�m�z�+�Z��i�l��)�.9{���t#z?!*��Z����V�X$?�&�� ^g8.�8�}�&�&U�Y��e��}�+X���:��ހޭ�yc?ق�?�k��	�������l����G��Sr�Y��-W��0{
b�A� ��=��x7d�uDy[�Yq"���кA,�M�Wؖ���jH�9�����H�'�?���� ����\N�H=�x��܇��&D�{0C8���qǑ- ���ˬǊoO[�U�v����"�xHX6�k������|�� ��H2��s����b��>U�َ*�ep��Jc�2
9~[�pnQc�M�]��V� ���{(u���8x/,���Ծ��ę�HBذ�AAP�_�tN9���N���	@Q��ܺ�2X&[;~����E��Ģ����X����khE��*�(�]̽�큇�[�9����
E�X��?`/��CE��d��Q�MEWS�=�˘�:R7��)�Y��E����)�8�`�%��Y�^M{{{^c����*���n�����:���(׺2²I��"����f�Ab���5m�ӓ}ӣ��[�˴�׳@9� � �nY�/�Ϧ���U�}�#�R�8nc��y.�Y��2<_���󏴦�&ρB< ���_u����v⪓8"އ)�u�Ql'<Zۉ1H���De(KL6�G�Y	���T��YY���$�K;;8��AJ?4�q
K��}�<��+�[�C��˵oa����y�8E��NO��c�G�~���䙸b�\���/����O��#����΂`1���G��~~�Yd��x'���f=�>�6�6s,9�N2�]t}�P<�P�'�$5<� 2����pB<~�$!���A��Lw�Z3�iIM���'���)�P��&�I~G.F�j
�,���W-'Q�� �l�pG@ܫ�	�EWTAQ�T�"4�O�Q��B�~�d@�S�*�"��� 1����ӄ 8e�{�;��g��d,��t������}��X���;�t�������U񎤬`�jI��/�������x��ۜ��<KpeI�>I	�EuT}g�F�����`^1��~�"�y���-�?:Gj
t��gt7ߘ�Tɕ�Čl!����OR��ßau�K�����љz�w���V�x��I��	����e=>x!���n���,Rnė�W��.>���l��c�SlA�:&�F�J17�m}�G�j���!,
f�}�~=</�I�b�pJ��ԾY�B@#q����t{{7	�J}�ӥz�wf���Ј����Xc�'%`2-�)5�?��˽�T�cЙ����d�����v���긑��qu��~��~,���&CbXe_rQ�d�%t�� .�l��J�A�͵=��5Ϧ��z?�,d ����V���$��]�����֜���ϒ��k�m
H�FP{��#� 6�M���p�d��3�鸨J��r�;c�Ɏ��`�7��g����W	<��k�^�";��p�aOz́�^�?�)"�KK�a�\H�X���|��'�	$R&�Љ_�*b	4�7P�����g������~��I��ր�K�2�=D ����N-����n�'Ϧy�mI�]H��vo��«�|��5v����-'捉盼��L��ߞ�2�)8$�=yȍ^��g�j@ⲤnT2<�6�Č���i��z�si@L��1w���7�-7k�y�4R�ﳜ�����r'(��^~���Qb�����ܣ���I�8�"�
܆�~��}���_9<<l���E����A�/Y���c�σr��U�7*	����~Y���#I&v�>Q�хq�a�pR,p@��9}F�I���8kp�RN5�G��H��R�I��"���x9��¸]ߛ��r�d���_D�;j��.UC��x$}\�2�4���'����p�3�^ھu��� ��D ˞���(�"�B'��E�{N������!އ����\�i��xc�8K�z.��7�`C>�0Tc^���-Id~���5e��u,V��xS��ڨ�����-Y�叉��yy�Ž>���D��<@�f�V¨e@̇��p��?̵��MjA�������rȊMy���1b,z�䎪4��Z-+��ORaL���d=�$θ�qJ���f,sFj�ir�¹��"�`i����N-czWf�W�6��0�7��=ƈ@.�$[T5L�c�|�G�s�T�~	� �Z���!�p?�ژ�H�0������:&#v���7����/�m�5A�>���բ���*�t���~&0
�гJ�����m9n�y�Ĉ���e��H>�Vl��3�k�U�s�o,��..�����Ի��_��tMװ���.$�a��z8�w�}����=�����Ӧ]���N7��.o8��n�v��d��a4�(=��C@�A�>�h%���Y�8��A�JAI�s��<�A�0��_�+!��<�|3]��J�F�](�+:�d|�������ǉbm�IW�F�;We�э6//¶����Go�/���O�}� ����E:�W�C��i�G���?�p���6���;�:0����F��2��|")aA�)^A�����bǁ-��Y�媇�L����Xl�NjW}/���,����7&}v������N*={}��<�_��d��%��I�QYI��\�蜾HPu�r�s�I�Cpt���%�r�t^�{���|�Wz�nDxۧ�z����b�0Ŕ{��_��V�.�ZWp r9"��{m/H$�����|F�HV�^�� ��f�6>�i��{/����5��ia�ū<�y[��q&B��,#��J�Ī�\+�-~v��!Z%��ḡ���~T`W���y{r/,k��ɽ�F���g�n�7"������'8Q�A��B"�pV��[C(�9fj
�6�Wbl�J �$���S�q;��a!��պ��>�P�硾���@�{�W'���޴=��̈́X!{���cW��U�+T�$0;�}���=����O�b��&j�zTP+�4�Qyj�ܤ�4�����i&
����Gd��*CWe��L�3JD�@Aa�?�i���xQ,^%u�F{��a�/_^͡;Ī(��S�~�)�����H"w�i��5������N��w)>���3w� 99��\��N���U�t8'n�r�='�����4��V=����W�~��G�ສh:6 ��cz��v���wAo��t�$���.y��������.	�XBp�I/�pz5Y�&�e�J��E
�n����b��z���|7S ��B��. ��^��͈d��|��-Xt��h������P�I�����X���}�� ��o��&���Z��7\TT6z.b��K�îrX0S �=26���1�$��&����Բ�]�����\/�i�u2�3$
HjP'����s���$׾��J_f�	���C8L.J�x|ب�r_E��n�x�Y�nߨ$V����Xd#B��L�A������T�>֠�2k��\Hm X+4���*�糝�����j��%���������f�A�'?/�A�<�y^E<$3uB����a\��4�a�������o�X��RHH�"f�O��`������5Z�,�k�#�]��'�A:@\Pm�{]�>_�#M�qH�����ڊS�(�}�ܛ���30U���"�  �A�Z�ש��[>�N�p��";rN�.���t�(�Oլ�;<#@�iN,�#}>��v��`���f��r�Z��a�ڳo�}�$�_5L*���"��zj�y�DJ

�o^� s�b�~=�k��w�������	���t��� D�20�}lqY������QV�J"�\��ǫ�]���;l�<M2D�sRV,5��v�l�.��쇧p���i֣xH��2�N0`�9Pֵ�#R\�O:��;%�����zB�EbMW���X�N�
貔� L	e�]Hӹ�D���0�ɢgB����þ�K�45��F�¡��D2o�qd��Ҿc`������d ���틾������jE����x�r�E^���`�c��'���H�M D���������v����|a��.Z)-zWB�L���-��\	�$�n�t�4��ٲvt~I�Q����/��&7��\�\��;F`��B��k$�0B����Y�~�J@bK�;!�t^a���Ġ���ʧ��� (8�B���;̵�`!�,���d��
fz]h���� �*ǋm��*�K�B��/����m^�An�B�n䴓��}�74�GB[���9��+�����(����$i	P˗mZ!s��+1KD^�����:x��)��SOLyŃ��)Bj�b1OG���f7�UX��a�W=)I��������|�-� ���S�;VDÙ(!��z��s ��c\��h���N0)7�?:(KD�Z4!�'�H��7�g�e�(z��G����ӥ�SV�����Q%��}a�~�O[��T͸�)���s��(�z/_xj�'ɑ��[(��B�M�xWP��Ͼ%�_7�q�Z�}�Բ��1�6%����ԉ������/w�R��Č��8��~Ѯ�N�\����~%둜��[ňSC}���*�]�	;�7����% Q.�':���͌>�%�د��`T�i�pWM?Qig@(�v�v *�KY���:oQg<��|���q���-��ÉL��d������ym|���{ק&����N}��	$��q9E�~8����^��O�����<>>>H��$-e ?��{�H�0"$w ���g�e�����o>�e�����j��ze������֑� ��9��.n��i~��f$�ӱ�`9	WVǑ��i�?���RQ�(,�L�6��'��b��'�!M���W4<Y�SDk�$�c.�s5�v���8ݯ{��wB�ٔ=,R�M�3�,9R@Uv�V���^�E����!@,r��)-��aT�-��}ľT�܉��LP��H~��s��SI����Z�v��f�2����+�j��Y��TT���߈A�i�U��m��4�yp7����il�5���]��1kS�B:3����,���5!@�o��b-n��ݥP
ť�)�^ܭ8�ݭP��Z��]O�o��7�=��=׽�g��_��hf�!]f�[|�����dXͷ�?�`Z�,>է?.�S�i��uSW2��hҒJ�ֶ��-�� �p�\��'�5��r	'h�"E*0��~pCp����	�?+�wv����EUx;�+�'"�yw8W�P��,�SL�s����W��w�d$�@&sW;�-�PyJ���r�����x��@��N�_��?��ĀC�2Xi���c��7���阘_�:�L�D"��[��Auλ��]lY�ǀ)O������r�6w�;1P����zAu�jG�3�C�q�1n����ă�
�9�)<6�[� 2���՛
q8w-�+�*{hl@� �tI�S�{	�#9��xW�C8�H8�Xˌ�!�SM�K?c�cS�C�O����pe}}}�/*�F�J��D�?������j����'�� 򮷫=�2�q۱����%9~�a�����)�緖��Z3�墩\��M������瓗���E[������1)<̕���苏g��,��yd9�60���76и7ᴂS��T��W�I�L��.�~���Q�P|�&��ᇛ�S>�����t0/H(�w,I�+��CT˕m��~~�A�oD1�S�Gn�+R����r�l:� Ã济��/e�Z��%�k2'KM
]��}��][cL�̥"4I��K�0Su�̋��5{p���1�@Y6&�o;j�K���FZ_�T�T�-k (#u����d�<�IT�(���gs�\�VL��'/i2����)������b'Dd�]6����0,�~�~��b8���n*@3�8�����dj�s�}u�-�,��S�M��M�E��@3a�fuT_%T�lv��"��)w�FBę��9R`�xr �K5P:O�7P�%Ӓ�g�X����K$���}�-T�GL�r�-�s	[�>@��F���bsFE�W�H��[���/�|&ley䄺�<�Y�6]:B��b�0�[��H� fi���~՘����E	���F���k�#B���O����~���#sI^cY���
��E�ȇ�E�]Q�P�QI�k�:�������N���u'ްX����)��]������21��&[ܙ����\b0�Q�;�H\~��cD#_5�0
���J+�)1�^�ǜ��H��BJ���t��C�o�G<l����>�ĩ89V�3���S���j"iCA3Ύ�PK�B��PN� k�~�{O��)|f��+���e����v����-�E�ϝ��:���Th��2�Z	�a�m4�݄�V�v��z�@��&ܔD�I�K�A(x C�EU���\�#-k���K�ٗs��4��r�`���q��,B'��*;�fn�RI<��KC|^�[�?���y���ʊ��P"�:���cqqI�cD[kk�����[�{�
C��y@z� ����-�ը�r����?�3GGu�e�E�1��n�ƬO��1#�s����B2FZ2�GӼ��R��>�2q(N�ݦ;�pAN��*^&"����leA̽m��\H?���sk�����B�Cy��c��Rk:Zs�Jд��!|?��1���O�U�g��|;g��
�7�+��%0�8��wm��đ�����$|0�r,�sa������9�]d��m������g<!o�e�
���6MMF:�2/������3Ӻ�J�i�3�����{Pnz�Ư�|��Ϭg#�-F�ĉ�8*̐5~"�Xm�V"�����8����b$�"'Ǭ�s΄����]R�]$�Ytgસی'����%/�BѬ����(���u}iu��S'��E�d�����'s���}_q&s�Z�+ڝ��5zs&��G&D�_��3l~�۹?*�L˿=�y~��g\2%�(޻�RG��g:��G//�IV��"��fcfJbՍ�҃��o���L���RFal�~pO�@������cs�r��x�ɟ�	mL�ϼ�	��/ OE�<�cF��5r7�^�m��N��ι��G��/>�FAG�'ծ���O�R��D�l���t�������A0�W��fo��o��@��#�&��)z�8pV�؊�����m�<���+\3d�G�y2�Z9��X� �8Ւ勸�߽s񭅐�}����L�6,Rg�����J����<�)�6 3s���ia�*BGtA�F��F�®��@��%��g���
�2��6#����YA����Ԯ�5�Td�rA	u�%V��g<����e�z.��Z�")����Ӗ����G�v�3Mo���R3��/TMQ��|�U�]�8�*\�cu����}����
&iG�7_�r��t܌ޡ�&�u��(@��_΂n9��.}���0-��/����AIN����l9��R8>l��A�B�u�7N	��:?�Wm��\�k/�<��С�3d{�����u��t���*�8�"f���]���5�h�d����*π��+@IɅ@�� ������Ë����'�Q�/+���TL�v�0��ɿ.�+�_��]̑�v�7y�jcs؁�ka�d�U-�����=�R�J+�4p��
���t��1C6"�}S��Ƽ���|�M@��������<SI���Vo$[����l��Pʩ�|�ѽC
H>8j,w=ui��isq|d��1f�/��!ߔ2������-D�����0
�S@Œ�u�Ш$��Ӷ�W9�?lhQ)�"�t st{�	�h���7vNw���Q.�;�@����|�>�ԟ�JBO�a�۷}�e��S-k4(ңK��	����(((,�7�c&��}��#�UI4	|�:��c)(��͵I"p��b$����x;e���*���θ���BQ���a;��y^[k��s1���J�cQ(\���ϧO-��4©-G�u���H-'�P+�#�Z�]̳�c�x�E�`X��'R���F���0�\H��QC�^��<W!?�ccɬ<��	4�t�A%	k��g� 6���<��������y���x<�}�n�Q/I�	+��������Ι���Pe�qp�5�`0�~���}8���(gzT|\�Q�\�m��<=�1��,��B���� `�F������_f_ө��Nߧa�X�녇��֟<����-��-�l�]B�����Fhs��,���/��p�"�$�<!eGԸ��}���s�b�%��?�ʠV_J��%��p����"7F6����:uS�.���ְ}�)�'��فUX�B���s�����Ё�8%`��_z�y��ȲdJ7�c"%�����mx�9�$tQ���f�.k���?����J����{s��rW*M�,�{O ���<l�!� ��Ag�'�Q�N��Q�9�����c7d���o��Ql��]M����D��J
P��Z�ϧtE��#yٿ�qV��RS»Ӂ7�ؒ�K���Lvm����Q��I���_���<.�S�/�B3�|:��٩ (]E��!����愰�� ��)|�����u��(�IU*��>F$����K��p�nDQ��d��Mc������Q����g�T��'Y��1�:��T� -�^zܛ
�$e��q�R%
�!���D��
�!I��5��T��O�hDBq�*مc�>BR��/���#���LIL��u��#���O�'E�ݥ��9�l��&&��N��hsonHw_a��c�C���mmTa5c>�&�|���ɻ��f�f$'ߔ{��s�2�
q$	����Y8=����k]�L�+�]i3v�3���m0�����	�����]��Jƒ,�yw��g��|��o�Cps���=��m2D:)�������<e*. >��4����9�S�[jtײ`���n_�g��ᯠ���p��+����* �B���x �h�������Y������Ԇ��0�kY/�zK� g�H\�_���S�+�ȝW�F���� �\� *[C����ZS��Y���4b�d�M��A@,i}��Oh2�-��W.�T<���I�2�����l��^q�o6���?@D��i7���CE��V����Q�� ��������ގH�+�us#�f͉0u����i=O��NB���Եy4S�
�im6��s�0C^�q��O�=�GBh]�S����ЀT����*{B��{'}��|�۪%�r��9���ɳ�qm��Ԉ���E#07����9`y8|� �;=���i�<�U�7�D�Ȍ�C���MH
���I��~^�nO��pe
�I�q�=�Eə�prW�o��%�`�!�*v��(���WR�k���N=2���]_haf^Üe����E�����s�� �}q&��A��ϐ�IT�H�c��Z���]�:/��gF�r�hѝ,�G��G�ӕ�)���Exu�������T� ������h��O���WlD/�33.���6s�C������)���5�����Z;�� 2rꐶ4�'T ��^�-�1H �`K����"�L��+��N�	=��!����[�u�WG�o4��fM�����s�Bt�!�F�� �r�V�*M�,�/:��Uh�m��h�i���[�O��U�}�9Q��j��~W��ġǾ�D �O�;���WUe�QU�$����[�� �pf�6�+D�?+}�*����KHU����`�+����%�~�U��m�_=�e���QQ��C����Ӆ��!0=�C���PM =Om(�$�md���N��8���@9N*�@M� ��NboL�(����:@J��/F�߿��$��� �Y?l��?dTK���pŉ�6��	}� � ��+�c����N���ֿ�U�N�:O��}�ޫLَ(��
��Ib�<��v����O|��ʇQ��X�`ПǴ�Ii�5�FN���J��Z����,�T��.4.���#��L�m�M*��Xs�ÇY'u���p� �G�C�� ~�|Ǽ^�W�U7�ɵ����}���ƬM�.�������C��kFaA�>�z�eb�m�4��B�fM��~��]M��e#�[B.�A��7Jc��W���%g�D@��Ӱ��0B����g�huX�Zv�L/%q��gVH�P���q&���=�cr��)�g�h�w����,��ͅs��#���DSG�9�Xd�>�x�7>Ј0��3x��Z�c�b;p���@������!5Z��fԑ>]�KՉ��l�T�WLC�ޮs(�@q�����X!����-6N3J�c�P_����l�V���_��޿��+jl�{϶N���R"�c+��y��ݲ�?j��ؠ��kّh�^/��3��7���7�{�V�lG��F?��f퇘7P��Q�%��677���c���<~�GjV����'KvG�H�n��!"��
E��C���}ʮ�4�1R�fПӖ��Zd��mvo��}�N]ɔ��41��=�Z'�Y�!u:�ա� [%*Y���(�����d9`E��c���9Ş�(�N庍V!�"����m��M-�%�0]���$�YOƊ_�:Kqm�#�A
������:̫����ԞTZ��<g���o�褰�;��s����$�t�X�� ��wc&�¼��lL�鵙h�RP!��8�(<�Y���{q��8��/�ϕMK�9�����˭�j59�X�S��e�N#ʻ%�����#����9��jÖ󚑑��Cq��	<�X�j�)�v 7Y���>{���:|&k���̜#QUߊ��OZ�J�.��K!{*����{���q�h���J�1CI�?��>l�i#S�O�J��,�����xJʏ���� Y�e�`�c��$�3� �eY`�Ikmj�^�#��p���d"Ũ]�Е��BRb`��s��D��лO/`У� !���a���#�o�(p��{��q�q���^VH2YKn�M��Ob |�!l�2�:d��/�D~¾y������=��5�$��曷��)�1�J!���wK��
����c``Pq�B�*����K�g\6������=�Vf2�?�c'����9x�f�#_��{����#8l�
⺩&׾NC�Mᔆ��u �K�$
e�Lxa�I����O�1�b�-V�#���m��������
m`k�jDSJغ�b�
^�t�6��@5�fT�u$�GitU
3t�[t	����E��e1�sǔʮ�۸�� ��.�G�s��e���Ƅm���Z��d��1X4���kz<�]�L5"6��R��2�JI�9	Ѷ�"���.��ѷ��c�;R�(#�8U�\�̎Y����̮��L�.e��ց�����>�$1OR��W���D
��R�!����uBz�!��0�W��P��u�e�������L�0e�_��Rt��7�pO�O��t+�``�,�cB��f)6���"���P,��t��8��{"y������~C!KP�QLp��y���H�5ʤ�1Z��%vV�֝��ƕ�u�߅/p����I�^���o�T*ͨv�����胲��ŉE؀;CD�T �/Щ2��F�f�!\����k�TD �H�Ɂ��B����b���R<iϨR���1�I�c��߃]/Jo:�����6�hƂ�	��&�4G$
�]uM��I֡ͫ�<����AF��\٥�S4����̽t�g%�%�h7�����~ֵˠ�r�1N�aJ4�uU��i][	�E��B^:ݞ�1��6`�ǚE��U|܅���D�a�<��i�S��8嗔vU�^�e
�77�!Nt]v��I�m|B��-�z�e�k��] �v��s���?�T��u?a�O{�ɔ����a�e������Y�^w�6]���_���Y_f��`������Ck[�������G���E�.뚄�.	L�-��{8o�U��ck���k6��_V$�?o~�[մ��=)~�9o�[�vP�U��' ��&Dݖ\|RIg]b*Hό� O��|=�ΐ_ԥ�<��6�@�d���	i�t�k%ԕ��"-z������� R��Ņ�4+8lGU�Ct���F��l-t�Ȓhs��Wt
 <�}61�1�����a'������Q�6���8q�߆�W���V?�*(��$�HP���Ϟ=XƹY.�f)�E�AJ�g�H���7���c��}K�nlkSPTT�Hf	�)�M�NF����'�}p����]�B�����P�������fo����H�6>{��2nyk��(�B����ƯEEyx_��S.wϻ���H���vK1��� ͹ `�I�3��f0ћ��t�*��u��w"t��(�s�K޺?�NR�{�d��w3�o�0��q��\Z���S��ygN�65$��Ӕ�B��Qa;�,c�]1%�q��0GVlO(c����>|÷3����!f{����4��SKС����[<�2�

ܞ�q=�9-aUf����T�y������q(�^III�|��N� �'�f�bcz{?eKt��oi�WeU�,yX�P��+�o	�'����V�����ѱ�9}�R��� ����(�r������!v�l~�,q�^uO_��Y�o��)�i]�#V�zλQ�f�:=�3T-5��Y��a9�ҝk�!�(�{��ŉIW#�R>�
]�����qŒM3��:���g��p%�����)����Ź���I�*��ML��$$)e��+|d� U��PC2L3Z/�wd�����K��rӧ&�Z���z��o޵�j�z
8Ew]@@��!Q�o��&��NܼF*�my}�]T� rz�qN*�	� ��{�s*�W�ِaD�����|�[����X�w�s,�Q��ɭ�)r��Tߗ�VK��ؼ����2tÄ�(mC�������@�S�z�� '<u���z��G�^�;:���Gtf�.Izl6�3Jص�W����rt��a���p�-S ������,c���)#��R+y����b ��6?C�'O�����A#?�2aq$9(���8�i	(�p�M̮����������z�����'I��sl��Q�8����(^��e����a{!8��5Y��3���01�9 �D ⺎����W+�gF��iCd��a0��1��&o�M�9�y+���H����{g���7��r��F�3�b��q��(Px�
��x�����9Z��-���'�a�*k�:5�L��*[w�I!L �b ����=�V�  ���#�x�'0
-D�#i��7����F(��v���g���>z{�~��)ߨ�����7�h�{9�s�<s�r��W�`����.��O0l�p�=I�w+P��$"���a+O���d7��="6�����l�c�E�;D���y��P �DE��uo�3^ش�bxм�̝�eK�w~d�(��DR�N��y}IQƘv:'�A���P	
�ő�7��	+U�Ui�2��^�� ��A3�e}��|B�M/�aP+����T�s���NK[��Uh� 6�#��S� �4��_w��(Y�c������"@qi�h�i�fǏ���r6/��	^�4��&���N�y�Wy�.N��EN��Q������L(:37�fT�a��S<"��o��x�h�ԫdD_��X2�%HMJ��\7�3�׃�j�m��*d�����iwN4	C߭d�0�6��w*�{۴Bm䭏v_�����@Mn�=�� vn�<r���Ɯ\�i�n����ya�4$ETC~Jd�V����<��>�F 6���\e�^���r/5�{�(�#/!�$o2�{�c�h�q�/�Z�!H�M%��D����nr�����&���	���`�c~��U��sT		m��4�-�5��j>���}V�����N�`�޴x�)�1�)��s�����ca4�D�IlO����6��HR��G�����.RV�'�Z�Z^u�a�Eh{�1���}��eW�B�{�H�Z�L��&��Ͼ^���>����&�KQ������\�J���c7�`�,%5�31�I1�.�D_<�S�]<K�gje?�o�,?^E�+��ݻR����"����3�X���.T����<9�$�Di�f���_��w-�2}>���UJӾYX��>Z���LV�F��(E�]���]@z�X��v�|2 V�{A��I�]'��	@���H�HHᷛ�U�-^Q޸ *� I���/_�5H;P =�t��ԏ�	��-c_W]���R1W�а���Ϫ-�i����c���B��V��1�oL�ῘY��6kˁ��mE�I@�HP4L�`�GX+_�r���ç�<�y?
S�/��D�<E�An�ә�����f�AO�TcK������UZf3���[긋IQC��s�.H���Q��p�:����/�qą��>EA�$�	:�x��D!��YqӮa����`%L5�F��??n;a�P"~e�=_��Kp��o]i��aF���P�U����/	u�%�4Z˺��,A2\Z���~?����mq����ns� ��,w�QV#���a���|۸ �hȭtWNƏ��1�Ԥ����qi�d�xc�I �������c/ul��]o�#Gf*}MKNҍ�LT/Z�h�����@��L�eݮ���b|.'���d��1 =z�i����=�ˎ�ᕆ��L�Kj�X��&T��~D������c���l�y4h���C�kJ���X�ơ��@;a}�J,�)4�^����֛	��Z�	�3����$
�.U���W�Q�^�vŜ��q�xad��h� �ܝD�����O�tN�^�u#D�4�Zp���# l�����sun.�<�g�y��j�,��G�+��pӺOb���&7�%Ϛ�W�|���*��?�pC����� �γh�%�>�jVX~��;tiIh)%��;X�.h�5	��/l��a���E<q�tyھ��$Oh{�44��c_j��GZ��\P*�Aď�Q������gZ*i�}P���f�C�̢����|�UUU�����4x]~�S)S�{KZ_t٫l
{7�'aO|>� u��^I^�׊��[�`$PT��n�����l���"�;J�Wږ82 �9V��F�#1���;Fe��HR־�d����'4�}�n�i=)q>^����b9k��U�O+�3ı�{C�ȝ��w��
��S��[��z(u�,OOH����
�$�{9pךl����L0��b�`X̕kQ���������X�H�Va���b�m��@�A;�3*�Vfo�d�C�:��A?j},q��|��&d�UU�U�`��l?`|S���{6:ƞE����-VW�\&��c�P6��A�<nhX}���ab��U 9�cD��J�8���D���̬��$�J���v���ʹH���p����Eʞ�n��ϼ��;Ih��n0Ğ�8bk�Yw������X��W{�N��Sv�q��'�So{�3r��h�i lM��-��Ų=QI֗o���v�8)�	jf2	k�2ʪF>�6aj[n,�����F>�!�4|\��[!�V�A���z���pzB1�>R��q��=	�H�엍H�R�ݓ1	��	���k)``�E�rQͮ�ױ �9����a�7E֯L���_]8p�*AC�7��Z;H�D��Z*844T� �'Wi�5��5�|��k�ٹd̕Dx�~�l��e�i+_��AB�h�A1&@�Dڡ4V�������S����/�6�~qΖV~�^M|Pp�,o▴<ZF�w�E^�����M��u}$��,��P��Ϲ�&E[�󭡑bp�a�J�,�橪�^A�(d[i��TTR���<q3�n�&���f�ÿ��`����IND=��u9�T��o�L�	��ш�@ٞ�-˵�]����^���t��}�}�\-|
B-�m���%K)�&?��I� wbO0�8w.y9mW�B���b���bo����(�3�]s��GR����?�q��	��������yP0C(��*���Z����Odh�4P����h6�!Ԅ;�����"t@Ϯ���3�N����7���Y�82:I��f`Ɇ"T�J�����9�~b�bN����Q8��
��� 8���v<�Z@u�I��>BN�=��;��Me�\q����[��K�?;���F%[���W����r��SgB��丯���:l�U�t9��<.��6��m�r���w�-�d[	������G�#�n|=cf��FjG(i���CS�LDU� �)���`�o������J�s3�s��qv�i��h���1��IǞ�I�r��i{��jkͷ,�0A�ˌ&�*�f�0,6�M����U�LP*0�A7�:Q���.��_I�2��~)�t�s,�ߐ�x��&�#��9�_�����R7�>H��`�W8�P�cd6kVtA�5Л#�*�:�M��d7�mk�����f�(r@霧5=�#���j��#�@2	��ƨ�r!j��A)!a�y�&�Nō�9 p�������!�N����$����d�+>��=a����>�k:9E�"�dw  >^��~���fa��n��͸;���O`TR�7�?����z�y�r�!k2��,{l=�u݅|��P�(Cu���F⶷���Xw>ǲw
e�a��S2m����Q+@.D�.���a��g}jg�X���B_��N��(���B�$����|�\���G���p(��1�.��L�/��������� j��E���_Ә�z�3{�R���P���
���;�m�!@���F�J����h��dQ�j}��-�������I��s���O��?�X����{��$y��c�#[F�YO�XQ��2�0CD	�`�����;�q������~�Cg�{V�V�˳������JWA �`��j�MxA��8>H9>+�0������?x���op�u���]J��d'�����@���~��}�.���l��z�>���F�Μ��e�P%@��B�C����꘮��BP<���$4���W}
̢G&}����/J"|��_�x�E�	z�_Wh~� �y=0��^��lSeR��wA�<�p��L0���S�y���^����g�6����\�3�[序�M]&w�f����(�	�i����=H�*]DE_�n�fBϷ��\�?y��9�9��f{��۵�A����k�-T��0[:��{UIqhq��0M���`(�I� A�
����w����&
�o�DÝxއq:䪴#���|�\��z����l`��KJPϥ�
���u]$����!�u�~n��!6��I4z� 8>#񇳒�12��%P�KO,w��υ

9�7�M}ӈ)p"��Bw�Yu������[?)�����m�L����N��Oh0*** �N��^�������J�֛�	�9��w�r��Ϗ��{���zEujK�(�ݝ+�k�������p�r���~-Z�?-5i��!�?!���]D_�;���C��>[���8XY |���jW�,3n�gj����7sZ4E������7݉�*�2��-`�8�]j��}Y��x�zGHV�6&$q�6�ؙ��#Q
[��9L��O�|N��/dM����·�֩�I����F�vWZ4��C�	��ŮN�]�(ե�O���RUG؇/�D��]�[e�6���$�x7�Lf(;H�X=���*I�-`��*�aVR��G�=iZ�;�|w�?1��6L���)gg��@�?��b-�b��>�޳��ݗ܏%�0��^5wv��Nr(��:$2��{հ��\�vg��z΅����?��i)w>�����ڰ�|@i��ɀ�0��B�U��	�5{������e�<��c���1!������X�j��b,��~A@�ʂN�p��f�M�k����`d$	�r��}�\1 �����ή�*�!�T���ff=��:䦆t���&+e�Jx��tN(�u�����#��cgf�y��:�K<��|�~Y~���v����ȉ�Q�WU1>pH�J܁_���1���X8�US�� �X���C��PH��8�α�i6��Tb�_����|.ZZ�D:�q�O��z��b�%V+ٝ�.�V�'��W6�k�.���*9��O����_Զ �1@@[�F���:x7����NF�A� �UCu6�� 8�(�k2�]�aD�1!��K���T��lKB�ƍt3�!��\q:���l���;�����v1m�G�	ᥞ�v��ȑ�u^N^�V�����o��"����HSi�^�n��~	Q���/e���j����ꞢL`����X<p�8�R��)s?6�v�2D6B*}��L��،%�$:�d��p�띙U^� 
ҍ�<��*�v����I���>�rQ����p���N:����d�
dɃ�P�8{|-4@?�g�j��#-�@ @ÿ܁|/����a��T�?M�+����EZ�����9�b��-�+��5�?<�S�?��1��?I�����첛���G#�?0�)x�`�y��ظc���D��"�{���/�Ҍ�1�kW �2R4��d�������(5R��ؾ�����([Cc<Hbf���.��z���894�(�ξ&Cz4]���K����y�X�;.��BC��t��Io��}%�-��Ȳk���E��2q��/�����ۨ�0{�-k5n��0]qq��3و�q��j/V���,�V�f��b�N��T����J��
3 �eɹ ��[^������P�H8fOj�H�m����L����a5��[O��~閻��<ĀJ���]��8M�^?��Q.���_��e�5` <�����i[&x��O�b��ֆ�i�F�P�4ʻCf�݆/%1�c5��
��8�)�i�A�	�45�g����Ė�I6C�?H���z�߾��{���~�ds5��v��t�1�E�ؘ�4����5p9�����m=���7t��rU��_�,�Ǘ�����f�[>16s�H��,�y����H�?C�[A�7' �T��b
��"�u }5�D��Bz��v&���#���P���U�ݹ��P%�"���^�(n������G:Yڹ�����v�~�S�"�"5��m���v�~�5H�@k"�9�m�+��8�㻡 m�S�z(5���D;Vm9n=J* �KШ�-+T��}���Bs鍃wgA�����-��<;fO�a�]�͸�+*[�ޢ�GR��i����1�@k89n�в#ا(�I��Z���*i��Af��������B�ȹ���:k]�PV23C�w��e��� ��Q��#*���y��& ����X
:��MЃ��"���"D����p>�y���p`l�=��E0~F��a��z�����������D6����&���?��1�3�V0b����,�~�,ʶ漰�U�a���(�?�J��nƈ�/e�lȸ���
ƃH� �Ig�p>���z7s��ɼv���|�\��������4+Ε)�.����������p79����.W� 7�G�,��k�;�ް��{�
 �lU�#��-�>�.93l�a�hP��^.H��^���?�#��$]�%Wl��0GL�x�I)Wf��A6��/*��9�L>����Ї��QX��Y�/��>n�WC�WSM�W��޺������:H�ӌvh�	��شh������~A
 d��OY\���&N�������{����(E��IXj��zx�SKIӚW����p"�6'�eϬ�^0x��6S�ө��|� �Q�z��b|�9�6!O\�m�1��Luc��,���h�@1#�H�T��6lЌ굲�ˤ�ډ��F��9��/@#P,� ���� G�Ǎ�1�wO:?+"�I�@��@���������ݾ�e�$OZ
��DgR����v8�!ϯ�+���y�s�G��:��ɍ����j}�,�$��8et��&儫�q���[�NȖč���0���luү��4U;|o�9H�4��	,��'�B�"��ű��M��S|ltX�t�l���~�(m���m���C'	<�bٷ�[Z�f`!�8A�y���m����A��]/I��p+d��Ԭ��rwK���G�K'䂚�T���!ʕ�| 
��N�+Bn��G�'�B_���S��sD�%��rH2c����ݐؐ�Q d,y�:��;��3��,�@,��L��8�v&���	��`���~���W����S�'o
�~/'�����4�9��ֽ�$J!�{��]b�m�K\����i�B�.s#����R��߿��&�3ҭ?�ʨ���������[�ѷ���Q7��a��v�G�Z��89�e`}���۳w�07	����Q�%�볹p*�����:9�R?N�D���nY�QO(5�ȤjG7�=��8�R�c~	�'Ӧ��m���l"��k��|%2l������R�߀ލg\�ٻ�5��8ٯ`|����Ex����q��ߎ��U\���Ϫ8L��D��R4����L쒦�Y1���������.F��2�O �z}Ϳ���5ے�\��離�g�ܥX�������x�D��|�ND [��`'�wR��Wf��[�$��?dqt�
���g�lReZ �&�,��>/a�*	K�r���o�<��sWA���o'�Bk��"��Ti%m)�y����,Կ]	9z��^��0�uiY�g����s_b���*�FD���/&��o��v�۫(i���"jo5Sן��^ŮWS�2I��mT~��cV��!�V��G.��p�S�Ϥ޷*[z6\g���T������Ij{$k�v����N��JK���T�Y���B���/_1q}K��%3c`�^����T-�� U�K�������U�6��0�ˌ����~=��/=b���oRk�M��V�DT,U���`O���p�/���_jrȀ�C��k@��B��a��@x��+v���K��"�΄�� ���҂���d*,���w�HOq��v�O�d�2�� ����
5�����n��{��P��bԼ4+ˎ�%��Ta=�k�I�7�z�>�T�@�*�0Ҍ���%Pd�j �&�G�%��H�8[�q�u+��'ԙ:φ�lH�W��&0HmA�` ]��Wk��M&���`V�tz�?�n��R��Wo�a�Gl{\,%�^���}��k>]�Z�6���b����Q�(��}
���?�%��k�@l^��y��F�D�>e�*�r��c�ʺ�~��8����K5y��Z;�f����O 
Wm\�?��މݝߙ[V٢��*#$����}b�pՀEP707����)�b� ��n�9�=��j�2Y�|�[<�Ð�n�N8d|I�e�L�^k`��wJZ;_S�^=*���.�đ�^x��Ħ%�4o���׾W?E�}�ò�.!KHǒ�
H#�tw�R"),)���"� ���!KKJw� -� _^������ܙ;sf�3�{�s�̽�B:��Ԡ�\��mC;�	�x�˂��3Í�@�&�HA{y�6��?7:�
 vp���ٜTZ���O6{�m�j�۝����8�:84쒒�W��>>^ys+IMk�����bk[v��}lU#zB;+ń�m�6��)�C�cl�c�&EJ�Hz��#�B��.�bą2ӱ)��Ķ��S�m���J���.}�"�Zp���
n2b1rU�<;O6T��d����t��;m���`o�o�D��(����]P)&e)��C�1�����9X�i:�k]���c	��-y\o�'_�ۮ����i@��7���fB���)ŵ����Fԥ��-�,�"%Mԥ����&�5_y���&$ro�m�e}v�PL{a!D�N\s\uӥj6���J��1����BO7�a*ժ���]%~�mQ
f(O�����Ƞf����p�Q�?�!�
��[n�X�䝀ʺ_ ����hg�I�K�~k'��z���r�狒� �d�J4�_<�X"�JȮ����7��"O��Ne��+�k���C��=� +Z����A��s�]��Z\$R�A�{6�	ɟz��)jGV���������ۓ92�!D�T�*�a�~4��odl���G�
vʹ3C\b(�qY�~%��3��!�Qgb����X.�Ck�)�@��"��b�w�]�Ȧ��}����d.�?2���:��S~lu38������[�aV.���1Ip�y�w~茅�~����$�AN,��Oy�Ȕ8!-g�2z+����.�u�.��h�l��K���0�%�����{;ND��?j�'�,��k�F+�u=WA\6\��8
Ca��ix�w�cn���l��V����P���9�)Hnq�_�j:mҖ$�40S9v,�a��>�>�3�/��O�T����$9#bB�K$+y�[UHϘ�=���ZMբ����i .�5>.3�Y�J�������(� �0%W�{G�N7���bɊ��>CJ�3r�LQ[X*vh�}X�s�[�d3�t��X'��в���ذG�Fl�T�Ϙ�xd�s�^{e����){n�\��&F�����^\J�Z�]�X6�y��(�}��6s�xT�7��Q���b8��J����|6V��sV��k~b d�]�Ȅ���/��\�x�3
H#(�5�)�_�ô26����ſK%����C����v��߱?� u!�	b����.[��&�[���DV֭���6l{/XC{��M奣���dߖ�ۡ�ٕ��.�6�`9��/$��a/����mj^z`�Iq�-�K;%��v�ʖzې?%qN�O=�t�!G�m�
�._�Hۼ-�D&)�F����s����G���M�SL�t͚>�|,��(fV�!(=��z�\��u�ٳ:�Z�e�ٿ� �H�~J�=U#U|w�^�3�����)�b}>�����EKH�O/H��h�Y@]���)3E��%��zIԅ��3Fd�F`N)�3�XӺL	+�az��i͏����ӾR�5�j0��x�����Ҕ,�j�8��������~]�uh�F��Kjd�s�"+����̨�������㣯~�*����B�a{e[��0�=6I_B"��gf8�ʲ��i�Gl�z�����f��������O�9b��[���	%u&驸I���ْO��.ĴU����'�~"Z������<�?��!q;#��?sJ����G��D�'��ͺ�1�q��<�HP8_�y
�kPl�Ǩץn����l��"S����G{L��@kH\#���g+�{��65��8�n��>�Vs*��m�� jy��d�~�{8�q9��*�φ����ƪ׮7)ǆ�v����]O�qbT�q�����p��Վ�k��'h eՓ��>>���N�@��3n�;�b��� ����ܵ��ע�e��/T�E{]��Q�#���oYij�*/���p{���߉
8S��s�N�!��i]z�.�7L�Z.�u��}�|�%��v�BL�ϏM� '0�$�J�V�S����+��.��w���W�iC�f&��8d{V���X!�%Q�� ��~��(� ؎�� �L�g/���|l}��BZ��c�b��Zr�ϑ_NEZv:x&�p�ޙ�;&�51ЪcE�}v��i�1G�|TL�o5%뽄���.$?�4�<P�ׅ�l�>d�9ك��Eh���Z�z�X�C�"��^�(��Oys��)�:Z��>��Z�/nvn��;�:g�~���Sc�89��R4����hI�-3��_}��G���0�<��}/�������f�i^�;�5���[999K�ľ㴽��.�(�\��p�N�K���Nۇ�+��i2��+����V��Hz ���։y!�]��T[�d�I�z�CZ���-��Ʒ(-���̃�����U��߉_���q9r�!$�4u��}����n~Oć�z9C�I:f�g�X��E-��g�ۆ2m�|Ay/�u�ln��C����� !/:�-��Y���UV.+5�K��d�u�I�w�x]����!ma��=��[^���� 0))�L�17ZF0� �/ӚN�f�����OH����Ȕ礲�tV���v���yZ�s�%Z�ǹPޚ��V	"޼o�٣�]]]���x������`}�z���b��ğU;#� ����7�Є�B��i��7��{���6�-�[9�g�}�jC:������\y��dWڒ�5��-�/@p��?���&ۮ�q��1oDC�d�?|b���f]����ϩ�lg�Z�#kNy8�[c�{t�>��!��񋭵������Mݫ�S�#�d�17֍����坬���ؒp kj�K���1N���J淢�c��g��{z�b"h[a��<������	Gই>� �O�$|����oޯε�~?a�:�{"4~�A&t��Ί��.��;>-ƞz-X=�����4}�� ��_P�o�g�+�E�m�^X��P�����w��ǒw����DƑ��#S�O|�
v���L-=?���F���M����t*��̔�Qz/�����Ɲ�}��h@�<��z���f� �E�I���|�]\��~�����]>�L9���R+
5�jLA���������*c�׵oHl�������ϵ���K�Q�JX8n݉8,)
��iܹ櫌Yr⛌�r��Q���7���3�`�o��
bGD�RK�����4��4�E���.�S�>_B���4��P���2�+*غ5�5آ�� ����B,W��|F+HS2ь)p��5hJ�K(�΅!.�?^=�΍b�t��}��Ol2�����]B䅊���"[���]�q�΋�Bﬂ��|���� dsu��B��������s�[����W�',��u�L���Ɗ���ȋ�<�0�J1{�~Ӧ�T�+cD���	���9�Ig|��tOꖨg�=7���^�����߿;���k� �t��V�d9bF+�:&�*�?z��9���Z]�]�Ҥ�Uk�A"�D1�y�:M�=$;��̋I����ؚ�$-쇋�A1bbb��JP%+��X\��Ӹ���@4)*��Ӥ���Ļ)sfY -?�7��,������;��oi	�yę#�ǹ0�D�Y��9/A�|�0R�d5����~P�������Ь#��Y��I@�_�~x@ve� �k=�E+�%�v�^t�%���_��1y���)�ʑ$˶�\����=Q�N�����=-� Z@͈V� '�M��9��Ț��������\(�B�Np5sޮ�|�;�B������[����T���ݓ��e�?gR��lݖ�=~�������k<F�b�lr�T'�9�=��R*ӆ�V�6:oRH�<��ǒ�s�3��O[�k�jg�w�������Y7��=e4o�gw��+��m4,I�z��
�g��c'��㻙z�6wL<���uq�k����KcTYW!��V Z��VQcn�L�"s��=:Y���Z�{�v�A�HIJ{K�~�(�{��^=�kf� �=�$�'q��,�E� =f���@G�EN�(�����T��%���s(���f��
�-�$0��ԤT��jrNH��V���Te?y�_^y�_$2|#�;�}f��K۫R�޹�=p��t��^�^����%�h}�"���Q�x�k뀕�HΓ_�H
&��w<+ׄ��323��HD�{��|۝���l~.
�Sy2��
}�-?�l(�ȡ�=���]�`�?�r�&�[EB3�\�`���'��߇����H!�0�����<���2b��)�u��氾q��ʪӞ�O��j�JP��ai�D�M�e�cc$����F���^��Qa�R����)��d-;�I[|r|*ͧ��?������DOM�a�������|��Ԁ��P+���HX=����N�%�:�����W�*��_m# +�)H�^Ő�κ�o��Ƒ���̎�ew��M'�K!Ui���/��}�'h�O�<p�$�'r�����"if����ʌ�S�ˀ��֠RzZ�`Ɖ�������� ��e�\�K��w���g��j8�t::�xS�)�.1")���ʵ��(NTt�{�T_�k�?ϛ���-��P����&y�џw�����V8���E��A(W�T�D��F�+��P`n�*���Z
xH~����"�]��=v����9�>�G.Is��;[��Y�f�xO���9��ܝ5�
��u�������>>2���A	�5g�H4�������E2%sI��ѿ�`��Ǌ�.:�{������_ZZ
F��͇�Sa�`��f
�}?~9��󕋜I�N��#��3����>e1�Fj�I-P}>���T�l��)h{k���1���l [h��Ù�k�0 � $���Q��JpjӉ�m��P���1�
1���oD;-�t���
������!� 7i��B���� ��r9�$��;�0�Op��2�ÍD�^O��K���E*�\��7U�������G���TQ��a�B:A���t�謵p���ƙ�~��q�w����=�v�E?n���l ~�̵�K��^c\��^�:x��wc]��������t1����<K��������{������z�)u�@�s��6��o�\y�c'�Ճ�� ����κ�����ُ���yr��~��Ҩ��W�cA�r�����'�6�U�E��C��,K��mM2+6��J��m��墦v�4ʕ�;f��Q- �8D�sJ��O�㽂�_|���>e_d=̈́S�3.��&p?��'�E�٫��z=�B���Bh ���r�M����=C���]K����5�3��Z��_*��4!ͪ��������C�6z��%���e/Pnj���d �{�O3��
(�ӳ���gm��˓�8;h/�P��{yl	�H�y[�r0���L��r�YwR�N.�;�V=E�{a@N�[��{�&9%���	*p���� ���+��˪9&��٧|ߝ�����������ɀb��֍���A�k������a�H��0��q|
yN�D�Y豐j�����B=�y~����>M�!G��K ,�*��4zF��l�Q~2�]G��tųW�g�+��oXP����՛���a�L��.e}�Ƿi�^����l���/a��n�M·X/{(6�`;���Izޓ���^��XK^�r�	;�����Y����"BV����K0�c��yM��sKII2�T��nz?!4(,��2I���*�R�.��K�����N$�`fJ"��c;s1��o;��Be�3u��F�z�y�"N5��	���e�	��,ēLeM���ZkY�J����[[?R$z�x�q'��mi�J"���
�4X�r��߿Ǘ�"��@�߳H0��3NV�90��U�8��O-+�aL���uX�l��~�NA�{���}�O����OZ��W���u��>�$|�d�ĆB+O̘u��AZH&(�93� ^ ��u���0����Ҫ457_']���R�ǐ/p�3�a��P{:^�nXʸd���}[�0����<L��evx]M��(�����_pje?�/on���_��ٱ;�x��@9�SU�e3aU����OC��Ab��D����.�_��=w�$A{ku<	k�2��/`0�g�`.}�cwe����e�y���x�~Y�f��wj���`&��\{l�a�:ݗ��}e-(e�<9�a��FiA�Ee�Mj]{ނrK�����g�X!�����ҕE���)���i�& F[���V��$����#��	ﲜ����v�s�W,p�z�G�������5��� _�#G�"5,�韩�z�BYU�ϵ�����Ԕ��ͧ���1go�׶ġ��i������*V��=K8�C�+j&��(&���\��N�q�KZ���9��V��SM�n�v鋙�bE����f��Xk��ȅJ��j9��'nA�T�.�G��h��]0��`���H<�,�\1!�����{�1W�J�� �U	�|�]�ݟoݾI!��%�N":���ğ�����vԻ���Q�ʨIo-O���ㅝ�=2PMx��;/���5���7T{�͕�ZY����$�jɬn:ۗبJ���8A���u��Ď;�<L�eQ�.s��K�o�W���mr �,�֐���#�-w�6ī+���H�ı{!� f���"�;\X7���9 ��_ݢ���-Nߌ������d��Z29�_��_���5�(���v�ֿ��$3jl/��n`�< �8��"�e*�Sj/v,�
�}g�5��;��\�o=`$_�����:���%$�_ΩG[��vvvRg��A+'''��Ք�y��iBN�&k�>V�H����ۡ�<.$o���L�mNS�4��|T��rMT����ghQ��\F^�&��S�Q��=g���[�T(�m9d{����L���f�������5�Շ�������w�g�iy�h��,W��١�W7��Wr&z�K��Ηt4 �V���'��������`4؎��<��	:�@M,U����=���}�E��4�(��_HS��r�`��W�6z�1�1U!�!krl.a9 �~c���t�J�]�$����V���ls- S$D��+��q�=<�j���l�p8t!B[}��;�س+�r��a\�Sk������ʡ�fj��TD]"}ǒ������Ynԍix��\ʟj�F�Sp:���w������}#˸}Fw����PP�0���k��g�|�䇦���o`rO����>+��>5-m}�ƮNU�G	�/<���t!���ޥ���58V,{E��C��Dd�&�H�WHgTG�\r�5Z�xxbNg2�\"��ٮz��6r��M�T1�-�1<ƙ<7�k��ip=\�-��4K�h���c�Q�����u�$�Z�3\�5Q4�`��2̓noę�M�ґ�B�9+�І:�糢I�z��͗&6d�m{��Qp�)F���H�3��_� �Js%y��,�ٰ���(�)�j���6nE����vu\>�E��&�(�?���쳴{�mo�������<�A$ �}-��@7������e�f���b[KC�p�u�-D�y(N�Y�<�(���n	!�щ�i�|�X=�rc�s���撬mbJz�lwp��G�o�e�,ޠ��<<�b��Jpއ��X�E�3��#9�k	C�aGG���"�w�~�:�G�Z_R�Ǔ.3*E�'vG]�'wg���{
,+Q(\&hR� �3[�3#.'��9_},����C* ������L��X�\�V
��������T >��2+ �;R�k�{kd8�
��	��K>��r�vWjp�xo��4�q!v���?������MpD?����������P.g�� PK   ��6X\�
�@ 6 /   images/846d17e9-ef90-4979-be28-74fde6feb977.pngL{eT�]�61t ���HK7!]�0tJ	CIH� �twH" !�H7�����~�]�Ǭ5?�Ϲ���u��H�7
xؔ�HHHx`E9M$$
$$�_����KG��5d�ʇ�o#!�"�夵�M���R�{�η=l�̓�����Y�?�R�� b#y4��8�x�y��L�|��?$4�F��Fɣ��D#[�&e��d7�vpoHwn��1��<R�u6�}�~U}~c����X%�,��,�7������,�ak��n���X]u�[�l�Ծ�e�}����1չ}�^o���Ɓ��10\.Hw��v�bZA�ee��/��Q2��A@x)�$曼�����ꔧ.|�v�̦+�i��Z��cf��6d6<�|4T}�z�e�%��⡼m��Ԥ�)U_�p��&�!!T�?��ʆG�e��G��n{\�EEE��_�/t�d��S��2�ݭ0�2���g{���W�8���<��;t9��nc$����W!ua��D9z���%%�vNN:�!���}���=��x���ݫߏ�b��c�(��Țh>�|�kB���.�Ѥ�)^@�D�*:���7�2Oo��
�W\�������N8��8Fj��k�ު����֢>-ה����=O,+?8?^�Nz��k#.J��hAm6�ʼ�Y����BРg�K�§M���������7��yZjDN�%"����y-bE辪UF;�/.p^h�I5�i�#z���o7��0�9����hb�ZB6�?���Y�)X-G�&�^k(�"=o�v���Fը����ŉ|�y�Q1���t6F�;���u,����Xу���k����o;���m'�S���o�qm�E�EHE��uzGt��B�.˅⬆���8�nS�ˡ�k��5>'�u�ʖ+.������О�����J8t�!�����B�ds�lU����Y%�2;u���֤�Ñ����*U2���n>w y9�B)�-���T̛��d #�"��>��aHRr�V����X53������"���w��S�N�<-A@5-���8�6�2�9��]�'��%E�*㧑\����grc�i�L�ûLljDB7C��[1?�s�T��q0���_}�, 1#6W��Z"���J9���?kYZ��ZS�x����?��"�ߘ[��۝���'K
�B��F`�Q�=�}���%ҊRIZ�(T�6P�$��QѾSr���ȋ�7ʓ� P>C��dg��*М��2de]���QQ�u���-�7���m�.x5�b.Öc�q?F�g]��EJ����W�@LZ4��2m�KÎBKAu+~�o��F7����N��9}�_����wԳ�.Ol���u��3��Ч���;�#�:��`)�����|�-}�V]�[#&֘���U�NX��2<�R�UJ,��+�p)����-͆�j���d�~����^��m�5�8���l�s�JX|E�ɬ�����J<V�{�)q�����j͖7 D��4��w��B��{5+��|�4��h�E�t��igR���|Y��pw���
�e����B� ��oe�|�[A�c3\J 24$��MBzoL����wn0mx7Q䆳9�6����U�Z/��Fy�E�[ڣ� �n�_Ǵ۵��+�q�yo^��x]�x#�0�м��K�,��Y9k��Ȋ�K���������@��c��6@ļ9�~?�ӏ���?no�S�.��D���1(�����ҟ��t-��Z�xp�!xln(][�3��1������n��p]�	��ݤ�ut��C�>�F���҃��2At�w�'��|���F�N�:\���ѥ7����|�B�YUEN�������s�G��7w����k����pN"ĝvZ����n^B.�C)N�>Ke-��%z�Xo�e�D���1���5k���n��U'�S�ɑ5|\_�m��uD�¨�cI��T�[� 9N�u<��sW�e�K+�E�d��ˇ	�ͧrԐMI7�4�%�[�n�X�5uY��ߗ�Sb����J����P���\ܲ����T���j��?,G2gm�/���߅���!M�p��ji%h"��m�&��O��2tK�N�'�,)�Ka�bz�6d�˼v�J��ϳÙ���0Y�+��m��������N}�qy��q��ɋc�E���;j��c_�E??�m���=$�'�@�ȏh��I��k�@x�E�f�uX� u�:~HvM
Y_��GC�v2"{��k��"K.�b��Ԡv���.�{��w�X>Uͬ��᠅f�tk�`����zMT�#J��k�I�yӡ�m�N��qQ�_�1=V�g��Z,����?���k*����l�c������ׯݧ���$ͦ���|���~��4�Wh}�w��i-b�Q��{�w�b��k��X���˗��~v�*3]�hKsϸ$	c��r�ɂ�.�#$����g9[�Oo>֕Ko�J|�L�4nv�3���鋹�l�j��he܃=q�ƧļL<ov��P�{V�u0�j�[��F������T�
QTS�RرQK������e�ވ�-�?v����"�!��ὸq:������|����䥎����Vo�$��YQ��k�:;�g(]���g@�����o�T-Śu�lKj����l��s�8���c���X���٩�M[f�ߗ��hi��،�Q�_o��^�Fs�]��>g���Jx����Nߟ�y����B�&�0���`�kB'i�4�o� �	8���!-�k$��Mr�Z ��p���i��xc����ZB�p3�n�$�|N��$��M���w���w֜d�RD<�i��vV|���]GR�c&A�Fq��nR^?�%�K��<OK�����9�d�+Gt�ɱFo
��_�w�j�J�t���9�I�d���I@[fV��_���~�3�3xl����}�X�P5hܺ;%���(���?G�G�GA&�w�����U ��������%/��1(F�Ág߳[�`�m"��ӒO�R󼜏�+P+�$������t<���1�O�1��'����L���>h�=�[�uY�̫�F�0ᐟE��G:�Z=��"Z�&����S$����RƉ=~�(�����(�~Gok�Q���� 	��ـT�;����������8"ŨM�+\�|�UE���Yn������d>�//�?��z�����b��q�=�"���;.�/l��^g���D���gJ-|{��n�<*_�C�hq@2>\�KW�6�������~�aSѷI��H#K���i�*��1���u\Y�ˋ��ϖa�0ld��L��o�y>"j:��|�ܠu�
�c}��!��'��F�(�M�����?[_�R�y�� �N)��'��8�FB��w��M��r��V����*�(}!�8�2ڬ4!K�X������W��^�A�ԥ��F��X�y�Ƽw�)�m(���r�.�周�>�&���g��p�����0SB���Kl i��k���v����iiS8N������ƱB6����[�7��*h&.r�Fr:5�$����N	>!����6W�um���^i�װ�r�����ZH^�f��m��|l�O5�ښ��/Bg����-��|
�xR�G��׊av��SWY `�^�R�%�ի�	���Y���ZE������s�t�����~�H����)o��<@�yQ�$Ĕ�������"wѦ���C���q��s������	�M�~�!�������~�vm�[�0?��[Q'O;��_
B�տ��9?+����%��bϯ�>�k���pXɾZ�"��*��X��~�4G�D6b�X�Ș#۲�|SRr�w�k#w� ���/̜`���$oBX��)=h�#�)��X-�B��:(��A���-Yٔ��qsU�a�[I[@�V���t�X/�.����{�d.��Z���x�!����%I��9�7ʋ��$��b1d��v�;$���핆��T������������X���ZRj��a��s(��C?F��|Ξ�_���=��c�������E�XsX�4���f�<�F��V�e��[��J�#�� ���:���B�&�����?�`?"�7d�V�pV����^���_ZD��֯;��TE�ޛ���v7ul����`�������I���ǂzS��ѿ�Pp�_QQV�e܈�g�D.����i�9�^>��YCH��z"���L>UO����Ǫ_�:=��Zڈ_�W��!& ��i0P�v��;FKJW�I\0 U�hfr��9T�G����P0�H0D\���X� �5��)78�����Q\={G?�����e*o�2~�ζ�c���o]���Fx/�bgW�X��)��_�`��D����3�ۃ��/���-��Ί���p��h#:d��Jk8����P�L*��Ԙb�~B�h�7)y8:��u={z��<s����7ʼr�A�+�)���?b˯��w}~�P
���e.���6�;�;`���	�����;i�K���G�$%����M����B��o{�{��z��$��nRd0'fQkl��b���FU���u�v�W�y"CgL�:dx^�Oπp
�A_����[�A�i��W�&�j��i��ň������K��__�L��*��� d'!��?�����~���-O;���a_���I�3���9}�H4�6�m��<��A����.)D�5�������F_��G�,6��9�R�Qr��e%>��%l�G��*4�'�6L*)������_���§r���;�I,�j��m����ڍ_���� 6���:�H��"�i��F�W�C�l]��ʹ���L>��Ī@u­P��#��K�9���t�遐�b.�5�쥊�{�c!կ��&˽��$��l�)�t��G�B�lBK����橃��D4l�c;�����e��p����?����&7梫&��U��AQE��ۂ-�?d�C��*�)�yd�	�)G�Ak~��2X�>ʎ�ю!�P,= �pr��!�8ҽG8�}ǁ"���2�T[[_0�C=���o��H=�9,�xj�<�hfg��E����*,>z��I���;N΂͌{ooX��4RF)�$�e+ L�Q�Gk{�W9�7�9#P��I��+g?��f�$�z��X7����G����gҵE��_�h`�N�����q��k����n�?���I`V�/���Y�G�c�(��{����f�*M����a��$>���M��D���*�+����nZ,��/Ӻ���2�\�?��"��	~��������Y�F+��@��C��^��|��Џ�w�@�V�dnC���n��3�S�m��ܕت/�q�y�0ٕ����"w��#���OrŜ���铓�?�z��~��L��ü8	��	);p��c<D�� z⧰0�Bz��D\4:c2��,�K(D�FL��I���($rL�<l����O�0TI�<�����3��K$����	[TVդ��(���QnP���p���l.v���N~O�|0j0��F�ug�������c�����7���'o���#�G��[F~
�]-��SR��`��ت��7c��ʬ�~3"J�\6)ܲ�������(��f��#���}r��9@[��*Q��L (��N�qVċ�5Ɩ�S�Sx�"VM��(�}i*�X,D��m����3u�HI��!�"G���t1����,���m��7iqju��lN���0�@p�ϝ�3�Mc�������Ϸ(�T*
�wܖ(*��:�u��7Ю����6��X���e�D%n�������ۏ�?���p8��(�Ni1w�;��g�A�Rs��g�&�_��r��&m$�O`#�4~c;�j�U��
�BA����bvwh�T�|����w9K��*�9�Ns��@G�S��Y),=pC@���ov���H�.gt8�lQ":��3�YB�~:\��@�z@ڰ��$6P���m��D.m���Hs����:ǳ+���'�I��?��~|}�쳑O4�����`9���Ÿ�o�ks���6=.$[�Ą��#���N�|Xn�``�g{���!A��[��ULY��1��1Ê��
��-���x�te��9�&O+��{�U�x�.Z�o�*,y�o>�Ni|�޸�5�{R�O����z<W�_�ɻ�XC�oo���}ގeIs���Wb2ueb��vN�{�*��K�c$ 2�v D@�nm�8��MD%9�da�&�[5�դ|k�Z�ť�r����Oz�Y8f]����4���Ҋe��y���3�?��\us����4��֬L�+o�\��~�^<�sR�p��^yTs�5�G�#Vъd��ג��Un��^��S�Ѭ���_2V".pX��l���'�.Lx�mgK`1*�����ID���3��}7������%S�t������񻉢{u_��7��{<���π�ʗ&y����'u�^�4��㸏J��rw��v��㣌a�b�����N�F�[E�9JC\ ߇�����Z�������B��)ɐ�+�$��&oȴ�i�%T��4!g'Z����H5�;���X�dt����3��}�L����\��T�Y�x�S�쒘I�{�g����:���Ϛs��o\�͵'�wv�T�/	XrI�<Rl��W�^������H�q���� `�hDψ=TN4�Z@��P�f�g걮��N�h�l��ڵ���<�r�Jm��)�L�N�Q�<�l�J"�-C�>�\�z4<+V�~��M*��+�gBc���b��٬����vSg����w��а�Zu�����k8՗��*�O�Ă�..�NE��)�H�d@<Xb݁�N��x�Nv�ʺH��<=�03.I�)�
�dO4֌�Ѱ�� n%ê"O~�Į3�Z]���+�x����w�вF�u���[л���{}�l��,���r˃�,�[�'!���E���ƹ�c���ǥ<o*���s�mc���^'�X��(�W��n$��5{`��Y�%��x�\(J5����D,]�L��y��]%$�@ϵʶ�A�n���7w2�z���v��VY4�^YNc��U	�����S�5Z�aJ��>5���LjY�ӗ�k�{���E���̟�b/��՛2Æ���xoB��*����B؃#>����C�A�2<�����(��>�Q�#����=,��ҧ-瞤����"�1�G��"2$� �U��_�������[��Tg� F�8�l��j4������vb�O7]qпy¾�s�O�C����s����qAW������S�t���J ����uB���&��İ������`�RSv"�2?�zfd	r�	tq�-Dŗ�2�8��L^1$�[�=�#�&��
���)�r���,�e�xyD�o�~Q˖X�ٜ�3;-`�_{E�F�n~��D�و���jo��%ߥl��dEe3=&�*7�]����9�n���:�(i���*R�¡Q�I�'������d�j�Fۧ�����&.��7i$nx��ԧ)�L���w/@`W�͐�O����U׽�)r�T�A 
�)�a<x�pl^��AJZt�i���N���bw�"��w�=N�\���|���������g�ټY*���7ti��!�I�t�+.�O�r�H&���5*V
�*}��n޺Nu}�f��L
������F$'w2�D�a�� آ��z�j�{\�\K}ٶ���t(�6 �2Ȁ�|!;�Wm�HCK&��)���0�	��GuHs	��7{l�y�����{m7�[H���x��=���t�ٴ>��綳sC*��7��!�Og!s�uu:���b5���7R�&�:U@)+v;�S����>�_�vw��f��VKK��O�,�S�Q�A�5_�j	S
˶��A�;�{
��o����;�z@`�I��C �#}��I�z�e�}�PBA�ˏk�fϞ����9�++�/N̏tn��me����Y ҝs��ê���%&��p�d��-�x4��"F"�� ���{�Z�d���2�9�j�~�O�|
PO�>NK�h9��G_�7��gI�`��='A��dT�O��u[�Q���q���,6����O�nK�2]0��ء��n�R?���.�B��}�����̈�|�E�7�MS���Y�&~��t8�8O9�����s�����p��[s��w=�ޙZ�R;Bl��߿�7����P�l��#�g���
�`���n��L��w<ȉ����#8(r��>�4��k-��s ���c}y�J�e��N?}F֍#�H�w�:ܾ9P��m����ޑ�&4�Ƥ�ὃ����t����^����y
�ʇ2c������⅋��/�.�����b-����s/��L�w�����e�␉����{�����=�Ú�!��]�X<G������
o2�P��D;���m���N��"�ޫ{R0��,^���%��`�:_�0�E�0�V�<{'0����'�X�����S��5���L�����%u*�֦�����c�kl��-�D�V_M�����:?o/}Ƽ}�d�G������m����^������]���j5�.�_%a���\R�˶��G7t b��ѝ�1c
1�� �_����\ʔ�c}���*p�N���9L�T���d�ǝR%L�l�]�p
3gv�ܰj�F�e�����&n����_e�>���|�Ȥ��r��Q���9xc�vXvy��d��ޝ�Q/�޺�L{5�PѶ�Ь�,$v�bmOm��P�F�l���~
�ąZ6�&�g:	����FԳ��83dE ��[�i���f�.̷����F���|vS �{z���'}e�XM��!�w�2���pd�$��0xך�E,X.���"z
�9���`I�EM�O��<0����pc���7W˩ qК�d�e��s(��в]��]����K�����H-��{4mY��-����z���7�w��s�cA�t��I6>��cr�uR���U�X>�e(<�G'�a�_ˉ�������nRю��r��5��p�f�t��]W�#/��(��)>.��#�28�S�o<��X~�E��>�+�;2� �������A/��Z�����EfS}N7�R~��}_;f��;ی����
�`�	n�L z��i��W���@��8!<�Ni�Ų{�׿vv�_�o�v�����/Ihc�JȠ�f°N@��s-	����y|�r��
D��Q��k?ОZN 	�Aā�x(�%>�k��ޱ$A`)u�_��V�?��{�;8$�1gp��FsV��p
 ����8���!��{zp����g#�&c�T�f�JIER�}$�ԝ��c����� �]�U#�FU�A; ւiN'�H�zMp!���/P,	G1�q������5I;M�иp +��0v��X2��@d��/��(JU���7�B�Kg�}$Mʶ�p _e* ���3m��BIiiF�q�Hx�Fegǭa��pS�ӿ��`�%Tv=g�����<���V?&�s,��wzE=�T��֐?a����&��ٸK&�@q���.)�B�k���7�،<�B�?��^A
�8�b����Mq����U����a��a\������UQ�MA9е#��!�:'Þ�l�ڸ�Y�Vo��jധu����-�vpS?5�K,8����Rp���1B��uՌV�$*g'�g���/�d�fl�u A�hɽ�W� "������de	�z�c�e�g�.�a�v�C�s��j�Ù�X��cFi��Z&���̄��Cw�#b���K��^��P۔e#�Ow��N�Q��T)J {�K��S�?
����#� ����ol-�xA(6il2(�2ύ�O��x>�u��S	� !�at�p�i�:clȬz���_�8��s��q?u�u7�m@r>����I�Ά�9.�]vA�S�Aޗ
��I-	�;�r���̭N��������/F	��*f����V�}R	v�ԫ^��݆�ϥ�W� " y4,ǰ���W�B��2�&���@�l���+O�`��xQ��n���pf�����KA��x|�S���k�Ӝ��_)��ߍ�,�":�����1л���ɥ�\����(���X�\1��t��n��I\?M�d�}У�q�w�YE� w�}&��A')٤���n�.,�5=�-�T�,��J��U����e��z)lZ�5!Bz*o���95��U���(%\dy8
�i�`4О�~,��[25a8&!���fjz����	ol�$���M8�}�5��,�6}1�!� �l����볤Qgf��A�4"�kVvu9�*����]�ل�55l>]�?���0T�8N�^H�^fC��@v��_4)���9Lz�Q���̗$=Pt�]l��1h�(F�a�S����K��&���`��U�J��	�%�m�����*qL��:�U�0f�F��QJ}�ѩ',�e?��a��zmQ��B�1"oo_ƄX�?8·�ָ�L����]I?ˀʗ�7�}���f)�o�d��Zv��w�+7RpdF�M��ӉWS�Ge�,���'�U��8����U�_�W�q8#y�9`玠̸�]�x�
ؙj��mmŻ��B��06�z���l��J_NH
'k�M<��˹�0M�y�$H1����ڒM�;:k0�0frPBN�N���l���I���$W�uq��G�4��"��I�YL_��-�������27�~��;�Mo^�����V�:2��i���H��;�jT8�zP���
��<�̺�����|�o��Ґ���̳�hY��Y8l��R�0i�pL`z�Q�
�����g����D}��t��x�x�]��d��`�9�5�̇�Zx��_x}c ���}/=�Te��b��3t6m�]�.��U~�3-�;f����PZ3��KP��)�6/����+	�$��co5FOY�P��'��U�)o��F��&��{�l~  $�������Bb�(J�b�Yu�cz3��F�m&5�x%0W���G��|>m\�v����Ths�����N�JUL��N(3��uMv�w�� �2)��o*]�
H�&�yR���eC7�Klb&Q�/���%�C�1��g�yA�e�����\V=˝�:��E���zOӱ�rx�RQ�M? �}~����OƝc�Nϱx�q����1��
��.������8^q���{�o�����|���(ok;,��n����܉#O!x��t<M��C�<0�>��A�6(J�*�1A���&t�	��}�<?�I]��+�uPzm�{Wh����\?'	�|��#�c�,|���7'�Sl(u�C��D��g��릑:�d ]����6�}7P���z�tm�N*�}[��<���9�[^�ty�����C"e����u�����0�}��Sk�6��[6���}M�G��U�g~<��#{E���~��h��m� �?c����c�������2=�ԄSz�{�܎��IC�]�dE������b.ubl���oKp���4����ت��q�R��l���{t���Dr'�1��9n�΂�J��V�ò#��؃����T�srڨ��h)9xF�F�a!�ޠ�F-����<P���F�d�U�;Pр`c����]տПq%7JJ=�7εn��#�(ûn��$�+b���QA��e�-!S�ζ����>n@רLEg�(Z�.���Ђ�D;���oF��k��C��Uޮ�4q�I�L�B$���z,[M��R5���X����Qk��H��|J�h�heQ:��K^^������a�Y��%F�[\z��/�ݱ�˜�ٯ�F�ʕ�7?'��T`|
܌��V�/���7��P�MZQ&�X�����_��h���ޛgr���
�$1OP^t�q�v���*ʐԦ�
�������RQ��lڛA���FK���޼7,������G��at�i?���Zl_�<��`�}{\�v��Cz�Տ�΀PWE�����b(��ʡFMc�}�;B�	�R�Rp\�`�#M,�[�Cy6r�H��̤��{U�Y�|opY�������u���P��S��jAO���Y8�"7��V���gt�D��-#G���$g�9���	��$�e(��ng?:܅w�^ƋՃ-8�}���_�Ú�?$�������/�F�+�Ǫ�x���S�n�_�ձ�YI�s���?[˾�S�~�y͈*�E���H/��*<�EҚ>I[II�]RG�.�'
D��CG`�o����&9��;(���6�h����b�H]Ձɥ� �f�F^��)�.w���mI��\����o�P ^����ݑ��&8u"v��t
���.�+Ӣ�kn)�Ϛ%�U�8.��{��:E�*~L����O-�۟�������W͍��Kc9,�كO4�o]�����KC	�Ξ�&��"x�4~4�#q߯��n����Nױ-��0~fVBT�L�}�]�D����#ք>Ev��L�΅�~w���`����z�#�Z�5+����~tZ�ē�y+5O`t����4�+�ި��:�mF�n^"�f���@�bU����4��p\6r7N��ySQd;�0�j�F����$Ʈ߂.�Kj_F���ј\�!�_C�DS����+�kt�g��ڵ齵��帴&���:�<3?���ŉ���#����J��1WA�L�J0ZL���%�`^S��h��	%��z���
@��\�:��>L-�� ����6�i��+g�����E��a��@mM�X��[dWa�e����M~�ْ0PH��� �=i�=9"@�'�Ȉe�eﾓ�b��!fK}?��ޢ�:s1��-E޸�W����K�'Xf�M����7��,T�6셇�|�#|�������[5����R��|;V¹Y'X1K������_��2��O�&�(�����0�#>8
A?zn�[��rKd&c*�R���"��횝dK:��Yj�ȓ�1��i�z{�+1�ϗxg�P>D�j?kd�G�U��m��,e��b%3yfƘi�a,��7ĉ���>į���2���#K��3�U�/�A����Ez��m�׽P�B�3Q��KL��w�)��{�3��JSU�q�g�#�I|�g04��-�d}*T��ϐR=7#kGWb���F�f�H�آ��)R(G#�1�RkDho�@��!Lޱ$�n�@���k]��J��{��	t�_E@��H5g�ߒ����t���!F
�x�A�Re��Q����xV�,�C+��#���"t6��TN��f��y�R[�{Q�y��sy�d��`C�F�gǫ0�v���B�y��M�)�7�(�C�����B�F�q9��Zc�MK]q䥨3�@!�{��1{��C ��� O�N	-�h��b�w8~;�/�Li4X0�Xo�l��  QB)����x�[Sp�k!�Ď�m�f	K�"�@ǜs���[�����}:��NB���A��a@svD���=2k��k�G�f� ��*��Obm��d�	���͜��nU��T5횯�C��N�JKt�a3��L����}ʹ��<�̓G���[���fꜸCP��,��� �2��z�7:9��-�L�X6���uw���Sc��3*g<"�~Lt(sI�&�B�"|�_�^��`x��MF�����x��'}G�7�$�8X1$��i�q�*9��:��
�ܙ�M��qV��[)A}�t�P��` ��lW��1�c��h���]�H7��hZyg�B���GkF�ǌ���?�|�/1��'y}�J4�T��<��@��sz�&g�\�^{F�|F�q� ��}�11��wG�$��E���v=em�<T1hw����;���
gj�M��p�tHFo4��d.=Z9Z�h8��i���K|�?oJAD�d�A���R����Gŏ)��u���c�͎'��C,��ʣd	O^~���u��G��4��ΊK�H�����tz��	9�����$��J6�S���+ANaV(�#ᵭ%%��Yo~��u��lZ��vY�oID�`q��إ�>��co���N���)�7	,�Lv8����秼[�]S����؝�Z��y���4�!�]���ἭT�B������x�knz�������U�q�L�B�/&:Re��Ma������6�-�5���ϝ���;}���z��	h��o��s"`.X���#FWl��5���L����1r��iZ�}�)��1c��{���z8����%����R�lCٰ�޿$j�G~\��o)4B�̖]������0\0LJ�$p�ש����@�V���z�����9�WǓ��o�G�Q:3G���͚-
$ME��$ڮ��_T����HG�-�e��4,4|}�����nY��(�4��m�����~���綮X���t���¦�FZɑA"��b�]��R�71�ci�f#�~}��:F>�k�6� "��I��H��x��Ɠ�W����C)?c�/h	a�1I�mw��%���|���]�O$�u����qA.���I�NإAk��4���c�BD�y���a�A ��&a�iC8�0١4����3�e�'i�$�q� �<Ǆ�r�6G������H^���5�Z����)G^���y�aP�NU��V\��6�����m��VSg�@ �*=}�!�0�i�<���yA$�60����"`Ǆ���(�`^���`�|���^�RY8H��huqc)KTn�Sˢ���wtM�K�[�T�z�����-��0���s�&�"�t�=�8 کu�P�=�|ť�0��2y�;�����Y=�?�1�u����V�k�_�8O�Fs���XXKG�7��LB����&��#���6?D�]��S���8&�㝲h ��Nb��@��������f�b�C!-E�?�LP����Yỿ㙯J��<CvШ38��w��Q!=,+}aG�(G�>����?�;8 �����ɇ
R|����^(�)!��d���t�Z	z�6���T�$D�4V,r�v#u��{W^�VR@s��uᖛ.�M��ҥ��+��p���H��1^*Z[	j��w�\`¼L�"[iR1sx_�mgfk��S��ݏyG��P�Ğ���:o��_Ҭ��3H�Af��~߾1dw���nQ5��������Ϻ�T!h?�N���'N��]��oW.wx T����A����oD^��b��NH�ԍl�Hȁ�Y�Td��N86f0������[�0FF"�Ѹ��°܍qY�B�ŊU���;�,i�
�0��|H�'�_�t5�*H��a�b�<�TM
�0W�Ia8��R�2%�}4D��݌���<݂�N��y�AO���r&.%��.�;t��6d��<��Td�L^��(���ײ��<n�T��)�Y�m��:��s��
�d��Y`P�p܌C�W^k;9ź�2��M���kLR�d�ݕ��Hb�Ҽo�ϴm�m��z�y��xF�UNg��lP	�{$]�ыUd���^-Z�T��	R��U��O>�;D�q�w	؁�n�U�����ߵ�� N#Sk.��u�4g�r���1�I��\ǁ�e��P��9:wV��c���5�˅��wZ]�Z/ׯ
>�o~��Dˎf�=���'�z�BpG�TI,�O�_d{�߬�i[j���vq�l��M���{^B��{�#!�����S4��:|̙|�-��3�N�sM�PC�w���s+�@��[e�jQݟ�z:ߵ3\��؜��
?1.�ǲ�6}���C��<���'���u�{K KQ&ۂ��eǗ���X���1q�H��<���Zw��$�:r�gp���;	/6�?1�#��U=��d��̡L�˿�
��YBz^���}J�����LiT��Z#��4����u֐$��a��E׽\`d�J(Ǖ�B#�Ū��a,��2MvAB�c�Xڜ;]s~G��l!»�Dd�q����X]�x�Mܒ��q�$�5ƿ/�:˟���k�LDwW�icE�E�3�չ�L�î$T~w������, �f<��h��<r�\q M��ڱZ-RkAz�!hr���ck8�pl��~�z��?(�P�H�?��.������$�@��\�+�t}$~��j���i6>����lE��dwW����~d�aS�u �~��������ʼnT��L�� �/$/(�����݆��iޯ���r�rz�tD_U��[��{L���H���Y��=Mjl?	,C6��t��ɖ�TG&~�:��W�����q)G$i�`����|$�P��t�mZ~$e�u�o�BR�9
�F�������]�����;�@�%�_ ��Bo�ֲ ��	a�1��i�G� �14*�T�NNǞ��� ��*�J*��B;NA�G�W�� �SE71('�x�8��Sn)����6��O�P�Z�k�{θ�hW�#��7�:�a�?\|Qs4��O��0��I�϶5W3�ӈoʟ��S�W��3���fz�����LFA�qH���z붨��{x`�������A@��CZ��A�[J��NA���������~s]���Yk����y�$}��h�F��2�	O䗺>��fH�����hv`�E�"��1�'��6鱙���"{��7����>�H�W��qr��I9gqON��Y`$^Kmbq.4���P�ØO�����5��@;d�A�1���(:
&�Lr��C���ٖ0�r ��J������x�s�yi��s`�nGH��"F�e/���V�w?�|<Y2��(��Ɯc�?e����co�K�i�qɬ��%�ު(�u����b͏T��'�U�����ݽ�w>bS����� ~�r�u�H|$u�t��V��'�I�q��L�+^�A��`��,�c�]�i��n���93Z�p\�е����	���7�
�m� �{���	�?�������~��%	�#V�$�{H
�|ԭ�R�(��<�[>y�w�ZX�ib��O�E����m����n����� H��G�M͒{{�x\������$|�`���lq��Ub;m,�-1�~S���D`e}����X��!���|^��6�;|sծ��-�('C��%"�����׍|�_��&��,�)�Yyc�K��q@���w�C�J�_j?'K楀����S��q�	͘��_�����}��!KC�O�-b�H$(CE�����E'-5ۅo�К�'9�W%h�`u<����s^�����L��ȿ�|M�v�F0�lo���c5�M�y���O2��-,,r�
>��d�^�5rfP�$ u� $�h�[6��S~չ	U�,��<�΀CQp\�p�st({zZ�(�C��u��B5��w`ߊP͵�-�0�>�7���S��i�D��#�c�d�f�7O��c�͸�<jQP!@�2Z*'gG�^�i;�<WQԷM%|p�5M"�;e�U"���`)�*I"jbB�1.�M^k���'���y���h�U��A
Ofh�������t�w����e�{�*hx��_ϣ�
�YoQ?;���/VRP�!Zz�C�k�|�Ǆ7#4#3���DV�$�q�T�\�iDBYQ�Ѡ�d�Y�:��O� L�( �S�p�K���p�}�1>4=Hgw�W�H��B��V.7��9Z%y����,����Ӊ���<�ٞe(*9�9B�Ƣ-�S����K�|�P�qd�	c��糺�:�9��9:�6�R�j>V�H�/�L���eIOA�b�x4s���ϰm��ݑ�䴾��Z�Cn+^g9?�	��1=6�����t�c�h����lk���l$������k o�\��I������Ya��K�I0Ӄ�K�/0a�Ly����u˖�g3`����T;��r�bF�m�a�,�J�\SFo����%O���K�`��${L�ܽ��E*>��ًW'��^�7�(w���څ�T�}���[ sy,!�h���<c{Z�
��PtzT?X�;QBQm��V������r��?�Ko>�&ƀ����t�VS% -�������Ѓ��h�ر\�r~�{{'vՅ�����hڎ���Jy�\�vJO����n:��d���3��G�߲¨������8��JBK�,��}VDjn�)|�/���h/n�_��__"yX�IR�O���[��Ҡߝ���P���� �m�I<k�z�ѹ'�/D9���e�3K6�n�[�������O�����A��Ŝ�I���pp�����ܽ��0$�Y|`�NX��d�0�Z@��ƤC�������&���\��*NW���.�V��M�s���uz����>1�lB
�a���`��c��v +�~���Ѡc�8oC��ذD�K�k���«%uS�%�.��'����YbE���Z���(�
�@iΕЇ���"=H���5_m���'π`�-�8�B�qr���$3�!8� �$�((
!�ljGD��go�؄���B�O��#A�:�QO3%F�L�� 	����㢷���vԜ[o;Eks�܊�q�ȏ=.-�ӨA�P�L��j2C����R�e�l�����smC�U ��G^@y
�|,
>ƾ�.N�~��bT�r��"��.�>)-��ǽ8�\������xeJ#��1ᜤR%]+j��Ȥ%��QY��Q"f����.֭��M�DYMM�&�����o�h�*�tָ���5.��X֓N�|���W��c)]TB�g!���,E[ri���K�����XZmB�
0�L���B�E����Ƥ�o7�Ѱs�K%��V
�+$��w&��Obw�����_ZfP������pJ�� �+��\3���"�ay�8�H�JQ�(�`�ێ�c�H�7�
U���!�G
ͻ�[_j%"�����$���P<43� �x'G�8%�A-_Z�u��B�N��E!5H�B)��˜Q��1JU�59����^���6�	����Ah��nY���ls����=OL�%Oժ+*4��+�i�AV^h���|��I�kE��V�҈9znfɹ���w#E ���L>߉�Ƙ��(�F��j�$ѵA�'?6q��!��0�}�`��+Ή	`��C1w��Nv�7��y�P&0t�w~���t8�*�bt�!Lj%�)7��(�9`��S.o"=�]����S̅ޣ!B�=���:p�XzO�8F2w<����L	~:��q@Z�:�"Cp�4Sn�����h5��t�IR��^ӗ������u�V��zA��ژ���Je�ϩ9���7�f�ᢿX�қ1�Ci�=��A��J��~����z��4%�`׮��B�6d��T�;Q�?��t�+Q��!� Cl��n����}�#���l���.��=�mt�eQE��e~Tn�y�D���F$�(�~��!Ђ`)��y������� ��M�!
���V`y�ٸX�t����6�J�a�m�g�����S���6-���4�OR0dọ���!9�B1�D���R"��N�|K4[\�+��K�$��rjݑ�����)q��e�������F���̾�����Rg5z,5�� $�/�w=�o;ik�%�ޣ���#�G�s?u����g��A\�3\�^],��a�:�z!m��B��򅑣������a����sA�s�2�MѪq[sg�L��L0&DQ��[w�J�6�����n֛� ���s�O�׼���t'6���3R�E�F9�M�)�1r����>[,�C<�f$B�k���8H.��O�+�V��+k76p�����& 2� � Bˠ�7ğ�E��N�c��//�`�qY�[q�za˫���oB�ӗV��=]���J藝����I}3_����<IrPc7�K�|v�w�:��*i��(�o'87�{�x��{���z�a<@�Y��	V� %R�JÝV@ȃ�1��f�g5NXy?p� �R�cM�ՙ� /W�qΟ��18���ɳL�Zꏧ�m%Z\c].��Cbؠ Nu�̓�8��� �Fƛ_솒&�+d�(�H�#ΘYe!	�p�z[�W"Ʊr��j���cj��F�?<����a��6�-ŉ�.몊^=��״��_�d�����}M3�՝#9�����p�,9�:=�\�|����~��ֈ~���𳲠a�n�R���RYZu+Q8 V�1b���|�
�B�B�l&`��'D5}����h(c�C@NH �d$�h|�"�7=J%���}�/��7����[�[�o^TRk�!p_g��8�`�'��������H��`Y�f���P�7�q����W{h@�ߐd�%�0o��	�h|�hP�b��.�r�|ǁ�Dށ���("�V
u�'=Y�v�)��v��շ����eH��ӊ	DDs���}t=Y�=�pjw`S��ϝ����|��-{�ߵ`�Dٰ�j�0�"�L>VնU��_k�X?�B�f
p��`��ЛҰ"2���e�>�ÜV��O��1b �q̱�ĀT�o_�Qo��l����i�JPl��@ڷfhj���G��Q�,?J\� ��]$8*L����GK&��Ʒ~�e�S���z%ԎɅ��W��ia�ޤj�6N��-T�G+->�m�;d��1�[����:��.c��riҋ�����rE2u�h�b��}"L�D3_� �k����/���?(����S��j�RD�c^}� Q9kY���m^i"f��ϹQ��=!z}�_��Z�K狆��=l��L�:�̒�i��2Y>�c�ͻ1�U���ۭ5kqAF8z�{�9,?�3���(�[M�u��0�1R
[�g����#�bC�F�fQL��Fie�`l�("a�&P�)~�<��#%K���eE���_��t9�.ɊU��O�)\:����V(#���%!^�9�R!�/�����$ju���\�@�vq"�"��\D"�1�� �pI�;�[n��|F_B��C7&���Z�r�zB��_���vG�I�42�͉ ��o'���`2�u�!̖ᕨX�4���W@5D5W���xJ�<��D�j�{vB%.�/�/.�$b �6q�f��$0��m�B4��k-����r+.�θ�)�R-\��^�o�Ѧ;)� ,�a]����w9Ǔ8�L�� �{cl�.��U��7�T)����`�m����]���.��ASc�`�4������H�Q��z,��Z?=�u��W`#�=gU�f��D���Z?�i{px����+n�.C��o9-7kZ������ku���p�~������?[�
&G�SZDI
��!f;�T9!�c&�,�U�������%
���aP.ݦ���@$�6u=���!�ś^�*O6e-�I$�i@
�3� �t/�9p5���r���gW�t�ݐ�]hd&*���6
椎����ݠL#x��!�Ť�H�MR6���|@R�ow��7�X8�Ey�gʩ+cF?��_�)N��?�_D�J	�1O�\�+)��A�	�q�`�Kp���S�����?�.�^2U8d��w䵈����%�w����*G?�w��Do;�=O	�MV�oe�`Z.׷ԋ�ɐC �|�_�q�}8#@��q��d���N��k隶���:2C��>D�hF�x��im��@��U�ϟO��`Y�w��"�u@g���ux��Ð�tP������%�{Ggi�u� }�L{!��쳽�p��S����@���[������t˸��N����F���ܢ3L��0Œ^x��U�F��@�[n|��X��?���[��e3�(:�o�A�ATn0�Ӣ�_�n��犱�ͦ����4>W�C��k_}dh� $H��BN:����⁝Xee���Dg�\Hp5.0̿e�NQ����z	��\$�2�f�Ơ;ۂ��<R��Mx#���5�p�)]��)[ 똻!���P�nT!o�]�z�e�'K�����f.�O���Pj��-�e�G�4�W���|�q=3��#Qn�4��$���'�û�����3�n�~�֌8�c1L�ؙ�z6a�F�Mw�h��� ��Y�����A��5�|�%���<Ά��"�ލ>T8����g�M~���ޔ
����E��:�Չ�4��H�۩����`+yٜ�Ue�edmE�D���
�ze`���"!$�Vۥ�qF�KOr�-���Z��Ħ[�XG��c�c����̓�I!���?p�%��6�'�#���:�j�w�J5����(�T��Fӱ��S�R=�B��9�w�wFݿ��S�	i0��o�R�U)|���� ��y6��d8A���(�^�%.����GK���5~�����>}!�9��5�G]����D�X���m�0	�����e�2�@�b?	��C^V�m�Iw�Y9��d�7��ʢƴ��7�[�^�g�9ڟ½j3��{�\E3�Zj��_��V��3���"`�v��5Jk��\�J	rM��"Ŝ	9=��h2jQ��<.U���Uq���b��U+�E�A:
>Y� �7�#�yѻ��7q6�/DƏ����K�ZԄ-Π��{y�3�<ň���B-3\㭂�Z&��r�ȣH�?�����e�r��P�x]�,�/p��|�c?�d�i�1�4�3�ݺ������$7��)̸�>�y�N�� <��}�<*���,0�~]��F0 �KG}��@��I��[�6���Ӻ?� Σ�
�܅N���!�}��o���r��m�ux��4�ޥ����M(�~�Ρ�w`zu�HB�oB�>��6`?g�'� ���"ܽ>�cDLʉ�w����C�1hM�s |ZBr�/ԝ���4N�f����s���!�x��_IPS�����/�,���s��#������x�u��۰�v���Q:�/�b�:ڐ�i�T���俘?��qyH��=���q�nV#k0�U��s)��7�zq�<�}@�-g�Ʃ�QkhA�O���	�o��>��/sVg�M+ᆵ��2YZ�[�ܒ3�� ��Ȑ[��|�H!����X�3&����e���w�9#�tu>�)�e)�ޘ�IⰠ�n�$ϵC�X�ǫ����:��	?������7�hUו�j�c.����47�j��*3��#�n�1k&q�<(Ύ!���*/e���$QJ��NJ�=����7v���I�x�en<��(W�oyzO)��";>\�HZ�8�F�����@�` @�meFi)�/�D������?Uh��q����� �Z,�
΍����i"i��\W��og4E�>*�Y�3"�&b6g�����͊��& �V���$Zf�HLP�Q/:z��?��Jd���e���<`���kd��+8&�'	�K��I��i���DD'#>C>��T2��>���j�叶�	�c�_#Iiz�[��2��j���xԾ�/�@���=Ĥ��Y~���i��}�f+�O�R�v��"�y��o�٬wɼշ�=���Lf��^�S��_�U�bB�	 3*
T��'�ϴF��~V����؏����U0���(d��e�ьs�^����&��=a���מkώb�g&����T��V+z+6��LiW���:j�~�	�|![�?pbb�0m�*-f�`��?��җ�+5[E�����8N������KI�o�*� � <J��ja�j�Ӳm�@���"m� A���s�mU�"�pX�C	F�@�<ii�t���[/���Su��v�_Q��X}�/b�����`��>Z���e���!w� g3c�~�������B;��+<(��*�B�Ď�M2���*h�Nkc�l�+E�ٌ_A�Er�P{���Tfxa�t&u�IО~s��_���&>n��Ո��dg�B�_�A�Ҧ�����'`�S���g�E:y��R�l':!��L�@ـ&~�UH�p��'�G0g�D���i"��"��f`A
Q�F�
��b�
�mr������5/_ϓ������)/���D�kT���H�R���H`L:�M����l�0����5��<�s������9��s��v�Ls�Yj�UIQ��T�������q̊�#�}/�[��d\&f�t�bF�|{+���������Y��Ht����Q:�g�M�y<��́�T�����c���*؄�D�iS�ሉl��gFlC �o݉��g)w�9A�d���m����1C|�$'��b�-#r���6�q>YT{� �:5p浪�tC�&m�\� ��-�<��k���yT���h�GP@��)S�2/��ܿ�t9?�M�e�����!ԑ���1 <g��;_�R�;�D�z�4�}��d���_����s_��E����^䆒��e�V_�C��+�D�8S��E���@в���TL�b�z�c"�C��5�Z����q$���Y}��4���B��A���`�͞2-\Rg
��i�!N�H���t��$�&���M�]���F�[W�.ܤ���t��kò�HW}v^��Rk�%b t�_��Lu_���LLG���rz,}�}5�M�}�h�.��u簹Q�O���<��و=��MumͪØG-V������L�oaר�o˙��R?�8w��~u]��4x��'�k��Dn��2��t���Rnu�=��_�5W��A���T����'��K��WX�Y��d���_�C	Fe��Q�OJ��>ʎ���N$ �M,�y] 7hg�-��
~���I?%��'<S�Ko��װ��k�8�׆��Oz<�qC���=j�p-�1�簘yI>ʡ���o��*�.8���)�oY/b����Y �bR�WYְ������X}�A����~e�]����T67�-Sl9YE�$�ry���Z��)�lB;��r	=���>��yjK�c���#�������s}��o<&�sXՒ��9�-���Q
���1"2�"��@���E<r7y�^�&���2����Ю~c��B1����^^�/�4�)�5�i��v;7�����+�������o����Fdv&%qt̚�g�w6��U�,����
��Vj3'��d��Ҍ$��rU������.Ӎx��BȂ���4�f�fD4���n�>s�"���3���Ӫ�E�*� hV��o������!�thZ�8 �#�Ӥ?a��x"q�+)�mª�]����G�ƙ���@�̄��ѐ
[��s��dl��J��"��#:Sng�����Ջ-?�(�~���ؔG;� D���Qs�Q&e|d��������C��}o*�T�R-r\f\�ԇm�o�D �@,�8[=݃����]-�84�d����*Mx���N�M����~��=b����;��|��n�ݏ�X�]�n�-���{������Y�'����O=v��.wk���4�?	����`����,�t�(�DX&$캹��ei�)�aKf��ű>�Y ��'-��қ��U��'�+vʙ�$�u�r�]��7��	�!�P�I�@� �+�ǵ	m�������'Hc#�ӨM����AR΁B����[�Ŵ��AM�q�qw�ݺ�6�x�16���U:w~1���(��1ə�Cѹ�.��̢�K�FI����c�5�x/g���h~6���yYЇ���Z#3��� �K�'��c�������8Z��vG����xE��i�q��x���4����σ�۟�(q��u߻�*������(���'�f|NV�3��{�G�7���z+�X��!Vȧ��0�U� �x���< ���A4:U�����s����g�JK�,=#�Wi�`��C
9,�ib�L�N��1SB٠�"��2�����4�8��ױ�8�����Ku�
)��~}��e�S���,�����pW�J����(�x�t��л��U��&)�`1�{�D��0�Xe>���1Cgk樚�
9%�v � �)���M{�y�T:�223���b�[�pW�q�z���hۥ;�oɌh$������-�5�F͇���)u�!��S:�\�mS�%�w�~����Z◿4�������>�H�/a�����8��1�-�/rj�)���:��܂�ш�M-T��t�x��K�g���+�ޙ��?eʬ�e ��if�v��T@N����q��A:���Ε>�c�t�g����-�B��f�K^�ß�L@'��K2�iaTК�z��SԶ���1&�Q<��y��_�b(΃��}9s��7F��C{���j��p�:\Wd�,�J�p�uƲ�"9J���e��CrƔC~��%�3� r��'A��d	h��aV�X1dor8-�](��{�;h��zq�B� VuT
�}�s���*�G�'�4w�K���x����g��'�z�N?�%�~!�mij�>_�����K�:��� D:(8��٘�(E��,Z�糧���W�V�4�dD1�\;z:��5a���4 ��z�����i,jŮ`qM�ȴ�=�_�m�13,�2�TZ��������}Q3Bk6l��-��c�	R�;���Dft��TC'�+�z�V���p!������)3����H� ���w�F}�?�[3i�z]�>f3�$��4��U���R�B� �@b(��
���u�t�`3�n�g��P�4��SA-��R�j��a�xH���4�B�t��_0����5�/ٞo�QpL�M�������սư�}:�������h6�i����oY�S37M�V��uP)to2Db�2�ò�=K�j#?ނ�{k���
ܼ1��		��A�]���+>Q���f���-HV�~o�� g���p�}�2bF����؃����]
@=�\a"�둄	���D�1=7�ZF�{�ڃ8��j(9��h;�q.�"O��sE�IɉS��E�aaa�30��� ��F�o��ũ�p��\��.\�l\��\���js��u��e�C�k�*h�J[c1�x^��P�lr�1X�,G�2fkw�_Ј��*]s�%A��TU����i-"�Pa�c6Qm��&tX˙6;77�|^S�v���Q��f��]8�Zֵٻ��u-�#-���;���!��6�L>'Z<�=͠Ypƒk�o��E�O�ި���Qa:�raq#�V���X�\����1 �I���h|��,j�d�о^=|�`JLYχ}��t��=@�BD�����	]C�D1$ꀐt4�!Om�ִ<hh�r*U��������s2lei���(�%����`�`\����0�s���x�\�@�u���H���T�A�AFM!>���rW�a��P�$���r:�SIfDnQ�gq��o�l�LwcU�[��\��*�K�B-�Uz��	}q���l8Jze,��Xr}f+��}9�c�͚򣶗�������N��+�)���[xj@!��ñ���69���F�=\�_��.rA6��Q�M?�v�V�ۣ�Z/�8�# �5cs��Y�	�� ���p�1u�j�Z��L�]o��N�ES��\�{8����kq�0���Π�s��*���R��:�zT�9���G��r�Ĵt�}���_n�u̵��:�+9��͆h���а3\���kZ���w�,@���=~�9�L;�;�^j"�,�(���E^�����W�25AZ��)oa|P �4�S�@�
��J4?*�T��"3���P l �yN�����F>x?�p~�'�k{
���m74x���,R��jZ����|�ohv�c��r�A�rw�2�j�OȰ�ɓ�����>ٗ���ȡ�,6æ�{M�z~�l����}q�Eu^��7��y���>��Q5�����g�S�/К-�*�����<�AȘY�0 ?R.�,X�r�{�肉���$�"!����'ɷv���b��<�"
NH��*�'݆���v�J�d��B�ϟ&�uZY ۀG,�M� N�� d�)��V]��e��2�f��h�uC�W��*@q�}!?#ڨ���m��i�9�c�����xZ��}$�<j��ESd�&�A�hg�/��*����Fo�!;�RDIAl#�ַ��MM�כ���B$h~(�����{h��x3��m���N��M!���L:�x/�mӵ�����$������ݼ|U":���3yT>����u5C�Բ�z��DXާ�D��[�7��	Ͳ"�X[�)��o�hz�6�����*��"������2�������]��!�3N�\�z��R�sYPv�W~���������>��DW+��_5r���esm����d��4픩�P9��&�*�fE���S��;�y���Z��$��se���ˁ^U�X�������'e|g8��������&�H���ȿmu&�)��pD�S`��!���u�NQ��y�l[���-=���|�!���ß�ꖍ���+����%�����:f�uX@����gu>�ܗ�<����]��z����[��nvSt�x�����;����h������}�	e�X�?��ȽtB1��4oi
�󇦨b�!��՜N��$��_=��*|^�#�H��p�-��C��+pGz�W!d���h�(	H4oÐ#�g�ɳ�t	����@������Ud���8I'ğ+8E7&���W?L>�l�T�1�VY��ܦ��ŋ���n�q,L�-�L�!�U����{k��U��x�[��F�ѱ���'qJ`��@�[�~��52��{V�G�f
�jq�!Q)37��g���7iqOE�'�>g�������ٙ���pt��K���m���*�|^&<ЩIo���2lrX�f'���wX�{��o*�v`<���r\������o3�f$w���9g*v�ҁ�83s���o�%�ң�|4�w
M�J�ohk�0� ���k���SމP��1R����%���#�ғ&؇��Z��߭'=��~{kS-���'���5�>hAp��gb\r�r�r��BG�3'�W� n�/w����`���Q��K`(�+�p�V*��qz�ힸ��Z�a����,��7�F67g���H0ě�����l�9�f��z��|6[���Nz�!�R�s��gb��e&�30�H)���-�F�Ӥ#��m
[�-����+�{�;����7��u�8b���b�coYt�O���K���%/�s����m��n� �m�A���	���N�~u@L�A��U/����(�/^k��MUX��Y~W��ή����p�i�8���ɹ��0���a)K��p���ŭr�w��3�����p�P��Q�U�a���Ҩ�F�=[�&1�G]�^�-0W���7���;�(�7QK��s9=-(S0�IjA>�!$10�����k>{[��y���E�Vƣ\�����-�˄���+k��w��̛B�k��b,r�3���ُ-���_�Y�� ���?�?.Ċ���Տ��we&��:���tX�*]�V���ϡRҬ1�p�P˄r=�XC��n�(�(�8�$)�#TSO`0F`2?��bDG/��[Kk�� (f$-���e��������M��rb.��F?�|��3޹S-<b�u�87x�u����@�4�O�����P�����؂�+޵�6z�R~a%V�^;�����ʡh�N�p^��ߔ��z�S8��L-�-MEeLT�e��2^�gg��55�gP�]g�^w��\��:��R5��s�D/F1nx���X-���"��k	��ؾ�`^�V�jSn�?h�s0ǟ��S����b�"`������,"-��Z����4�h��U�X)l�z�3yG ��J��}�\�knyc�\dޱ?Z�\�7�=!��O�����1��?�ny��I�	���PQ>�E�x5~�c\��$�w����F��&g����v���fz����@0)��)boƪ��"�d&�ׯ��M�)�����G�g EO�I����:�5��6��V�#z���q߲En��B��-�����"��_ �Ҳ�*.~���E)��)�n�f��Y��P�or�r$�h��d��������][��H�F�?z�F&nH�K�]4�H�U�0�ﺕ��-eIH�	�O��@�^�Z�94,�U��IPR�s;V�7�@�;7j�1�X���ч Sy�~x�M�m�՟��VT�v���+�"J%$b���4��S[�d�5!T��Qz��]G>C�O�]D(�e��dB���8�᲌#	����U<��i�S�˙�5� C��8�������Ħl�
�
����Z��H�gjW&)�<��{z�偳Z��:&�#��QX_�N!���y<����]蘾�탍���Y�gy���� a����*sӅu]���zpabK�jrX�jL��'�$#I��-����a��۶ֺ�U#O(�Q�)�w����0Keh��U��X��q�{q@�Rs��s�����sc�x-2=] ������#K���MM�ݬ����\���Y�����/�a0�h���O3�^v�#S�_�L��[�6�����T9��6���ج�H���}^�d=�6�p���ףQ�!?�QC�C}�G=~���Aw�`uj��X5�{ؕ�!a6&0K}g�;q#��3KV��'�*(<2GbE�XEJ���Ob���@
��"w�v\��搭�D�q�aÑH�ӟrrT$ԓ����N롬�.3�8%�L�پ�|��5jQ�d���2̠q��Ե�������"Z�����5ct���m��4;=B���a�`���Y� �	���pY^����>�f(���i��,p�~��ل�n��h�qA�����tݐ8Gȃ��|�4��d�cαy��;�ɧ	�e�5��i�;h�Rg�_�d��:]�K�@\�RhcCH�0��}�Yr�#
�`һHU��L�������;kZ}^y-�S|���a����XO�s��8�V""��d��98$�Ѿ"�<,̇����#c+�e_l��.H垿;��G����q�VX��
�(��?��D3~��D�Ud��Ft��l�vJ�Kfu.A�L�I�:͙�� B�o�ds����:(�#n���G�� uj����}KI@ ���WmZ�Mi��kŃ�,�w����D�5��'�`	/c�����)F�9�H0 Zq=`^k�/�ʌ�)g	��D����2~֫�x����
����d p�g�=��+g�o`�=��8n���1�<�nW:��La��Wq8�An}O_�PA�������4�����ʛ�*�/$Y��Oe�����.C��W�ſ�j_�A
�&�k5~��u��Z�T}=�jLDCN�ǚ��S�.�^>ީ华� ����y�J�m��R��aq����i��(�=��l�|/'T�e�Lt����gp��fg4ѯ$˰�A��9�H5�~����ʭiF.�Y����W���>����[s�z�vf�Ҏ�3��y�!���ff?z�'���֞�hP��Ȍ2��R��Gօ]�>%lQ0J�F�K��M����|�w�pv�Z�p"J뒽�L�O%��s���+�CH�T̬�~����fc�Kv�p%�'C�+�[!����f3��ǜ��bl,���n�?[$џ�m�"N�]GFFR��B���##}��W���Z����"P��^D�B0���
a͍,Jy�T�8��O��M�s"�@j���FI��EfHK˺�(qV�>=^�ˉٽ|T�[w����f	�3@i.�u�7��1�[���/�mOBA i>Rm,�S\/�v���#Т������pi�+1ek7���*�_����%ʙ��G'D�r�S<P!J�`^̏;q6]�[<���S�_��9|������^B*�p ��H��'�=j��H"=���/rJ�4�My0b,�T�_f�������h� ��x
��5���Y�`,��!������=�d$�i��,\d�yr�5�N�Ψ0������㎩.���~,��",����O����R`Q�]�S_��)��R�/J$tu�^$��x���o�?�8t8��k0�3dd�wP����d"��48����r�kF2�w�[L�P�7,G$RC�d�p�*l��8.R	4Nf������A�$j�v��UU;Ev�w�������Y��D7�����͢p�Y�e������.?l�����_U�sO�$����=���;��Y�~u�D��7���3�u�|,]���|:��%�]���Z�v���ř����/ō�g��w"�nWIS������1a���q*�����e�`v��D�73[��V�V��6Jq��.��zΜ��)mIF�'�L)���w����ç6++��a���&��e���o��v��{��Şڻ,��t_v��{�Ղ�|���n��O�%�AMi�T7ș=<ɖ����_0��C�ik�iY�w˾�1a\�i��ð����Q����٨�|��>A�uV߃�
c�0������ϯ4��������YQ����h��j뗇Y��iEv����h�����ˑ��[����F�2i`D�� ��*L��j�k�0l$]�{���$]p�Uװ	T��b�5솧�� �nСs��S�c����u���0*&J�3�d�M��{�D�$�����I�WӿCm�˓l���]��}fӿ��y����ՠS��D%�9��:�ptE����@�^�R�]���ϒg�Z��mRɵ��a�s��x:g�Y*�R�^�U���xhh�������$��h��'Jl�P5��X�L!5�&���'��D
�2�,������Y�.�n��ҧBs� �!"��X�O��Igi����g��o�r����Һ�����y�ƻ[	>�^
�8�z�&p!�煮/����K�w�������@��>�Յ�*~��'@#H�Jq�T���؀I8����|<kmy�;���@G�a�DX���|9�PqZͱL~�}Z���_��ȱ��	��.7�Y3���؆��2+++׳���Mc���\*u�{XO��`�Xq��{U��!��A\X�i6'ػ�ޱ��(�Y_��Xr߃`�U������fo�����0u�m�d�N6'��S�5�dL�9a�m۶&s2�����w]���^룵W�A��[̨��#�!��8m��,z>�{S�t:�-��#�qߩ#H4+ђ K��k��J���T�N�E���j�S�'�˙�&��ƒѣ��V�����.��8b0H�(�)�d,ݝP�$LZҙ\l�3�!!���
`>�@Sj_$��h`x�
s�e����dqBE�r���< �іQ]!!�G�r)�z�P~�cg�?8>B+^/�]:���A��x��Um�
��a~�ၐ���:q��`e>!�9Ů�n3K
�&���JnP���{*�ҩz9��8��MUF���*��wC�0I�P�꠺E�MW���&����r[�Mel��:2FlP���Z���H�|c�W���Ĩ��A)�gU�
���1�L��q)����SP�0�X��!�,���~�R�T<��t�db���毕hQ ٥'4�p�Q6 �RR�/��ܝu½��K��D)�|�:��D��M�Z̒�H��JVi���ºKu��A<�̬�Ve�{�۸���3�r�ۍ���&+�����l@ߢ�v�p˧��p���"ez��+����'�j�� �-�>g�jE��u�#�_B6��k�q�$��R�2�גe`В>��o��R�M�h�0��.K��S�28&s�?�F���s-}x<ȶ��ܔJ��Z��[}Zl��� a��6-v�\o��'�0�[.L�� ������f��%�x뢟7 ڈ �h�*���A0b(� �d)V|r��K,�f�j�m�&�玔��*���N-ϕ�WM�����є�3�#�(���$����F28>���b�8��Hc6�w����:jR����v�]�|���f��t����	'~��\���?T�j�|r�y/�������ڕ��-b�ye?��'?����O���+�M&����JlV�辏�q*�^l�
�)���[.�����A7N���I���;����B�9�^���FH'�#&YNw����%< ]�b������Z�x���tL�D�a  �z��0E�WĪ��9�Y8�p,
���5ܕ	H�w�=��=7��j�]MYS@�ْ h�l�p�)�N�6�,��P�S'�|<�3;m�^�����*M(D�-g��)O�O����PL�X�Ɂ9����ĭ
�;e�)hݴX�iR�"CsX{�J��qJ��%��^.yl�����h(?~���u@v�,K�*�����zc��z�n�"�m)��99�Ws� �H8z�/�EE)Ξ�H(6�/��C��5m]�2O�i�~=��	�#��:ɫ5���u��c���F���>H���h+&�ƪ�.����<�ɹ�p�w:�_WV��IY�"֕����vm��$(��p5!e<Ñ2�9����i�~o���_9�J�Ն!��eK�d�v��td*<ǽ�´�SX���8�!tJ�\�x2�/{Z�ܛ��nhp�d������ �hd͆��f�pŧE�B���=}�|��|3�ݐy"𥟫ߧDVp�vmI��|�3��\BNk'-O[���&��!��)�0>MТZ���l�2��4��6���r+kݮ��:�ylqo��$�~}hw'��g.�JE;rh������{�| ���3�a)C�h1�z��q0��!��/��m�e��|�%w��;�����
SIɵ��Ն�,I�@c`8�F�Ӱ���gP��-5-=bP+4wZ�N��_���TG-����:_�W�j/�F�cQ�wT5}H(ĢU��o����-{��M�h���ŕwQi/��6,⢧S�/Y/������)}���&ߒ[�FO��Q�7�Roݧ�(S&�M�|�%�P���NW�[
~���q%,u9YH�C���mC�Ҳ��s๓��S@��X��p`5�mQ��z�y���!�\�.�:5��A��5��"��?W�v-l�\f�-(VU�\�}���r�5����`/So��H~��dt����W]u`F�E\�$`�`�!����\�I�$T"كViܟ%osX��?�R���x�Z��(u��F�]�P˳��8�J�K���7u4�w�r�m�!�6AGg�78�Z�X{dR���X&�T�6�VE��d��^15F�o�=HU&�/
n�o-�iSǢ�xҢ�Y��7��ǡɊ�w��|�v�=t��{�t/]��I)V!.4�I ���(����3zM�>�]�}�r�HD`����xc�6C������0[�����Ϗ��WB^�S-�c[�tMo/�0�L"�՘������q|0�R4 �	(-����~�*�H��KN�q���� ��i�����0�aQ~Bz�Cj��o��y���*��/��K��ս�)�_GΡ�v���"��u8��8O���#%�TP��D����fy������ ��aLC�]������ސ��k�N�F�>�]>�C�㞊����,��'�V�6۹�i��l�G��?�,�1�>��{-¾#0�	�2CQ�5�y*�(�']��w苮���������f:�r$A�p0&l�����{��X�r�ٛ�a*aE!β</��i�(�K*�79��C`�F�
uɡ��`3��=��-�
���
����m���/�� J�n���yH�D��?F%�l��e`��+���e=��-��jB��0fT�A*$�D(�J{O:\B�gҳ ��!�޾�V�&�D�A^����~�K�n��=T�n��� �0׏���d�N��ih�m�y�4�
�G���w��������������%!���(}^�[���I�� K��`T��|����(s�	GZ�m�z_� �|jJ� =�)�c�2����NX���A����Q!b� k)�V�p�P�iFj3�
���W���'s����k��hey>~st��~�oM�UCi���)p�g�I�;������J��b9E��l��g��6��
M�Z��`���@��ϙ��j���n���)�)�Ը?"@<��:��g��󾰲�:U�<��x��H|w*"�^�[��XT�^�^�p�C���^a�pd�ס�~��a쩇qwd��e{�'�	+k�U��{[�����g҆=;�%͙p<�[�}���Ks�h��?x���E*wr�W����+230�&��[��i���;��0�8Zk�JgJ���6]B�~~}��P�E4͌�6�K�]�8�ǁb2x��c���o`G)���Ҹ���0c����	�x�HT�*R.��ͅ3��7�@����|�w������ƹ�VE��J��6�����7Z�,�� ��7E2U?�C�{���鞕B�i
9?���[��'�5*�)C
��gh}�`oYH�w�3��k����g��hY�Z"��̝:���?��k��k��OK��`Kz @�T�I�e �����[1�ZLDĠ�~,�������P�R�?HcH��q��^�(�-=-w�o���H�)SC�W�P�hsq'ȮX�B�F�p�t���4mQH�K:�g�O�$&�Y��jS�Xߵ�A����(�q��a����B
������dA��i>."<��b��h�H�}�w��f.|���ˏq�K���L�ކ��|Y,#z�9Ö�p���F�>C@wL��Uro9��a��|�����Gl�Z(6� s�&�kM� 9Jy6TԶ�����;�`�Rه����n�T:��gr3݁uX���o ��Z�[�Q�F���wS���FX9�.�o�k?/��]��xp�� �!�:����4���_�$��K��y��`���v{4+%.��$�����i�6L���O�E���\��k+l.u���r�ў�qN�����z���v'-�\?�_�@b�ϯ���uV�.g:��II7��\�;�'���˟tcRm�Զ��~8��	4=�s.��6�뿽:֔�6B��"
�d�����3���f������(���Q���!�h����*n-dotQ������j��RN<H
�^�F���V������'k�K�3_R���<��L���%m�h�1��|�i�E�Akq<�K���5<\�x'[𙎔t�D虓�咈�P^ZT�P^�I0I��j��H4��}"e��ٷv5�:~znɶ�[�h'*��Q�c{N���=W �`���[#QF���dC&9F�#mr�,��r�:d[���WX���]B��o^�e<��"����NKe���	�Ow�Q7�L(C7��Ip'b�R�],�X�GABh�\vHi��?OcA�54�L��.��%a�V`�e��(�V>�
�D|���c)�����W;���=®6�t5���$B����
&S��?ɥ�L�m�(�v%uԻ�D����ﾵ���M� J3��q9A2�m�ՌѸ�|� W8l��n�������4�N�4�^≇~�������x3�E;�w�@�00-���w��=�JiM��	�"��r��0����6d&Ȕ-`�����ZZFf���5�������סV�(z�u?Oe�ˡ�$�B�I�^0��F���ݟ�"��Ȗ����Y 3+�z�����Ua�)���7����g����|�Jdr�
��d�vQNڋK�&�
�ƨ��V7�����W��͋�x�KJ)�#��Y)s�mr��j�b���Ԥ;}W��rE�T����3%_q�1|�q� ��s�T鸬��Z�c�~:&��>��f'9�ln�Дq�а3�aQ�fh�u
�-��肂�"��׹��{c}��F1�X��_�#�/�]�4�?���0��Ƣ�/*!C)�Uwy���9Y<zP������yZ,Fd`ڸǜ}��D,s<�l&0±��8V��j� ���{�>�A�0�5���>�4#��Y�:+ݣ'|~6����|-B�÷j��'*ƮN��'�&�_�n�E:
���7�|�'4c��g��Z��f|�[���X<qYDreyc���aR��
��8Y����#*�SX��F {�9M�I:(v�B����=[O�-��$�[^mJP�tZM%]������!c!j2��y8`�b�F���p����<�qs�RhM%~:iZ��x�Ư��
���)�� �F)f��\�ˇM@l�އ���|$.G��vA4^�֣��I�2�@��s�{\�8��]�ǩ�Կ��-��^�NZ��*�r��,�j5�5F��~b��k�[��h��������������}V�@�V׳ԣ[�XR��u�S���݌K>k?�	��ڇ��1|j�%��'���z*��jItzK�L��ɋ����|�h����'A��v�>R�'ti9�&�ic�=V8!�> ǜx�O�;�@��-����x�Asn�]�M�$�%ξW���H��Ѣ5a49]�Qw^�e0�����ֶqՏ��6S�,�S���M8�N�iHz|�r�T���l������O�>{�h���Āoő�� OBE2��B��(V���!���J���� ˶Z�q�+�5pO��/� r�&�����Z�*0��ù������Y`�u7di�!��Vɹ�<�w��ӧ"�M��A����]��;.Y߾�#�H�3<��L?M���m��	���rlX|�il�H/����a���Vi��ZR�t��Ȧd�]����4%�Y,�\�{*��r̀�=���1X�~����Xs����tL��mz�O�	̹���L8�/��rpt��Xk1�p%��m �i@��:s��j�R�Ob�jY
v�9w��%%	����ƻ�
���k�p`�zx:��fW��e~���*w!��p'$�mۅ��P-�S��i�����=a����$掇ɥ��<��� ��h�3�(,�%J�Qi���p`��r<���sZiq�2{3W,�r�x����B���|8���.�b�\�U����ȩ��R$��P�?�C��TYb���@Ɇ?����T'��'@�x������j��n��Ϊk-MS�=n�5֟�Y�g�g�6D��v��R���XWWW�����'�f���Ax��֩��D$#'��%��uDnF�U}2�(ZS##�.y��a�tf�~��A � �@&r\	�3a��|\6*nP�Ƀ��)�Rs�Ĭ�����t�0��{U�"š�SMEf��QJ� )��t��y�ӽ�/vu���]�Ke<�WUUrl�k����s��dL̹����]��c�Nh��	G迆����vOɆ�w�EL�6�5�_U}R�l�����h�Yu�sE���w����ňq��R'D���f���~���m�BI|D0qp�E������k���9�}f�Ѫ!A[(��>����ɭ��~.����^�#CQ�h�>曨�[[K0�Vq�{U��L�Ok*�
�ޥF�^��

R���	�����x~1v��/Oz�;�>��v�z!5�j~��j�M.t� +�qƗyE٘|B�b��Ԇz�Ó� �b����Y�7ܞ��ҝ��8�G�4��}�Y�l�{$,����o�^lv6Nj����͔�����_V9���c�V!��q�8��cg_��R��+}_K��n	�ͳ�����č�&����-�7�9�N'���������)]��~��GuY����a�hv\�br��4�B/�"z�R���	���9��~� oJ�g�*��'[�3!��ZQQ�g�mcx"���V���N�NE�y�n��gkqj�ňV;e����1�	�l�X��{���R�u!�������6��C�R$�7�ss?j���4�뵉�|:\[{����l�m�,\z��x��j�?@��e�lP����Z��X�Lԉ�њ��.��G,�T���>M�Z��|WLU�+s�m��3�n6D��
�[ٗ%_�vjF�0R4�⌧�yB�^�5�H\�7��Mϩ�XD5�����O�:X���޼x���s<��1����⟫�����5T�����`�*����S�C�Ƕr9$(qEv36h"�J<P�E�t���Ls��jC9!��s��_��[� �'MK�N}��mKA���0پo�f��D�b��V��8P,:�EX�����-���L"�q�g�z>���˧���`���)1�3!Ͼ�����7��Dz_��Ֆ���>tc�����<E���G�\0�T�t���Dn|zLу_�q�V+��!��ܗ*7���7ha__�KXR���H���ѓ�,/�ּ���'�S�~��"�����yX��n��x��D�/����ޭ�t����D��I�0�Q����.��sO���E8�6�?m��n8ߟ�����niѫ�ʮLB��6��n�MLL�P�yo��%�y'� �}�~�����SXx�&�?�wp�G��OM�����|<����4t���1��Z��p����L��5Go ��7���Pw��0(�9�C,Y6��n��ў<�ӯˣ�V^TblM^�12�m��n�Ԇ�(��[�ܛm�����J����C"6�����J�����t+�]l||D�3P���kL�-6�.q7�?�8WVy�5�����.��v�Y�S}�Ӻˢ����\&$��B�u��t�2�º:���K���^�3/�lI\�]��;r2���Ҋ#7�݁�}��� ������(Bލ�&frr�F��Q6�:�nl�6��}�[�/��u*�(M� 9�
�W˙�
��|�`��蜞�����rH�lD'��6� �|���*RXιf�W��@ҏ0.a�[-��1H��}[SF+�~�`��Va�'D�x�2��}�A�ߓ�Qi�7�Y)���e�f*�h�wZ�����p�-����Q���lq�l}q��*��˓���L�a�������ϗu�YMk�L�Ǌ[߹�<��|�z1�����h��8�c�Ǽ�op�d�ݶ弜-z���ߚ����� �K(1��~��������L�v�Jd'M}�MvR:ۈ�����$LG;�Ɩo������f0�O���UhĜ�"TA,`o�#��
�Z�
���K�'s�����)1�.�t�'9�] i\-F�����@|�4�Y���|�����עL��U�K������p|��`����%l48��w���k��4��:M�C���آ���J��Bn�|��f������o��޹ڵ˞m�����c��U�����+�nM��6�$X����m�^�Y$�朆��6�9�-!���jC&�,o^��I9���J�I��n���Ug�8*�UՏd�4�!�e��E
��k�f�����(��"B[��3����a~4m�f���8e��_|�Vsƕ�솘A�َ(�UG�e��h@����\�'豱*��?d`Q���.��^���~qߋ��G���E8�ъm�KL	RZ~�,.�u��Rs�E���eg,�(�-�?�M
�ϵ�	N�#	҂٬x�א�~�d@�XP��:^�v算��5  �?K�}�c���I�~��\��%?����~��iRb"���[뺂��4Xd�
g��`F�D�fx�r���T��kD�]x3M݁M���gSӝ�0r..�vV��r=:�g1�;�T�,�Ram_�[���C1��7y����~�����}3o^���hi��S23�Ŋ8���Na*0"\��H�xڂ��g����-��O��Z��qڶ�_N��>�4�X�(e��~,<{�M>�!�����.�(:��OT��IE�s��U���+]��̾E���Zkv�.*(k��+�ϟ�/Y<aQ�P�S�e��������@B"�y��/���U�Օ�,h�(���~��?�W�q�\��}ޞ��LZ�=:v�S,��J���&r��?�&��h������Wl�z�l���꯮g+��z�-�t��Zk�p&�]9d���q3d�C�#*�:n�	�W+ZZ�o�<_�#%)h�?LC��U�j��y�`c�յYm��,(裧�خ������'>s�M�{������Ĥ�a����O��ޖ����+��A!Z1���@U��d��5OPљ5��K�YIq)".+92�ʮ�$��i���''���J��h�X��Uon�&����9f�,>?��:�q/��ie_���W%�`?Vb����S�,��ÒIZ���G����>[m|=}�=�h���mŗ���0�C?����<O��]�]3%W��i�����+�����Խ��Z�ۮV[�U��r;�LH�ˋ��8���������6�j�w3�qY�3V=��BBP�L��Tv���(:'SC�ӭ�斫�<��dn��-�z}ў�k�Cկ�Ϗ?*�^�]�7y�9�X+!/�M[,3��g��i�Zpa�M�����f������J�]��yݤ�|�7<���NP�̛i�M�?�?/����B�(�/��/��<N��E<�:�i3�b )�AX%e�֒i�<�`�B��W���ޣ$'�a�T�:������3��c�ܐ�9��#S#��2~V��{��x^�s���و���8� s�\��Q��Nl�&��<DL��4�t#_�1�Zo��y��sPz-#�~�]�"��-"VɔEPݟ��NlW~8�����O,a�a�T_5l���Q�����q��!P�_T������􂜅g�e������54�Z�V�g�v�^�`�t���DV�!���zH�@��~�0b/.)�jhL�Ԃ�.T|��i��lT/Ո��$�wS�x'�."���$	f�`�v2eVT���8��g��(����q�@�T��QՐS�������"|�	�o��ئ�@6t�݀�e��vm�	���ÿ�h���N�檪�󶶗KA��b��{(+�z8�5-�����W�l��<��é�^���a\��:Jq����}���o����b�
Ȁ���a^��\S�=�����d��������o0a[��D���rl�q��?�2e�Un&B3��ģ��0��;��YI��u��M
	(�	�,Ӻ5�
s�ruu%������)�⎍S~���6AL����ȇ��;M�~��j�^�	P��<�hʗk�]�-F����6k-�)M?�9�6:kPw�A�2� ������zu^)�[ľ���6LT�����2�%�z��B���
�����C �o�ْmEY�T�,x.�M�Z!��o䚴�F���qn߉���3��ت�n���j�P�!��hcUR_9�o���� �U@�}*Ol���Y�=*Ѭ�"�ΗB��!{����jq9�f1��XJ�������[�ճrv/������¬Fd־�2D��Ze�Ƭ"	���~:�޸�tS7�#Ytk����u�������Q���<�F�HHrt��oő���"ɶ�s'k	��JJu��{�(lS�6��N��\@(=�u�M����A R]��>;���r$��H�����V MюNI9d>�8 Ν�#xuϝO"�m@�"&d"���ǭ7|�|'敋�+�wT�k��'��I5KM��}}}�D|u�������ճ��N��ܮ���}��ȥ���h���� �+��g���
p��cR�6�fL"���I+�]�af������Y?s�1n��S�x�.TH7��U�zf����nx�\���r��wu��*�F���R����ߚ$O�Z���$w\5��d��1�d���㒓���Ґ���:��M�y+)�:�: ܬ<(��i�1!���؊�">j�>��<C�p3e���}���8*�g��@��SBD���8 \���m��l˩����vѭo��j���*^  �:��������`��%F�Y���|xp'�&%�M5�E� Ď���%f��XmR�+�)A��R�����#��B^K7ǥv��oG��4P �]d��ceI��3��"�M&������z��)�]��n�y8~�
,��x�T�W�B����Z�H�b}Б�f`�=(�pn�Ť�*ԟ����*a�WFEK(�b
����C��Y$�TNuU��3� �8��z�߉�����O.̴֛��0�E�
��^�[|1�

(�y��G{qY�D^���\�{��}AI��}|��a+�����g���U�����s�
;'=���l`V�h()Ca�����fiWA��fff���0���l���P_�'������]�8�+�J�������k���oʦlI��DC:}��=�ꘘ{_�>��
O���p�^���!�8�E��1((�]�ז`���z��l����l
�͔����������f���q9V3�+M� �kwݝUvX�_4H/���|3ՆJw��ׂ�@���v4v������S����1K���,�"y�5fr�9"P���T�Y2�}'�1�^��c�V�^�~���WaA&���?��C|,�����o<#�	�VUM!�At��R�Z�z�*��\������M(��-��$w1v:��7Z�f��"���~x��*S�l��ﵙp!���v��M�Lȶq�qʒ�4wXd�˵ ~U���*�"�p|J[��u��J�J�}`P�1/��GaA����|l��߉_� ���m͵�ޏ�1|A8���r�?*O�!A:dg�B�CʟZ,�I�&ox^d����1�@��9�jf�(�LY���e7���]EG�{��)G{�E��e��l�,����+L��X�E����ϗ�ʎ'�[�l������Xs��R@u��߯�U�M�-KH�� U�!���h8���ڈ�"�+A���f��l^}C"�k�f���?��>�~���ܯv���L��ͩ�f��˚���go`Ё,��(�X���+���4��^���T��S�Rg!i�yV_�4~<�R���|E���<�0�Z)����Q�XK��p��R0�><<���|G��ͭ�6��|���J��;�Ü�3m٦��B����{f*��=�o$ܪ����پ��CF{{{3���߾}?[���-T�����q�	�/��/�aaW�+�3�NL'�Ō�c>��M��8��Gqyָ����������{O#�M:���?O��V�m�Ս��!oK����e�<_9����w��ۼ>�Q��W��� 8H0����uh?i��hj�x�]Otq6�v��rr�����#��&���^l�+i`�Y�~�mȯ���?�!���M��c�f���c$laj`��9,����ۓa"f�gB"~g�ǳ�w�S�2���d9��O��Ӎ/�]{��RY<��ek��^:yj^�oQ2���C������钽�Iؽ��CSƋ�n�s���0.�X��JL�+˩�W�wz�|�Ȭ�d�e[�,�f�OAt8��c$��ڴ���FD`FQ�2Ej�e
�6�z�'��$6l7$C�X!>������Bnz�럮�u<w̛ed;�,���`^ط /�֋L��~����I(ff������A�<V�����"r��w�d���v����drQm��OC�J��@�Kf�v�$�2|q�cHr`<������b�Wh1�N��Ìy��܁{�%��lQt�tsR)Eğ0aJ��%@@�@��)�����ÊM��?���8���N1^��.:8xǶul��6�F��z�ԨH8ل��������\ �?� �fi`�u��6w���X6�h�9��|ٵz�8�k�������8%��^o5ޯZonn���L�l���*�u�PH��l5���a+��_4)e�9����0QR,���PB��x�u�D(��VF&���r
�E!$$B��X�Ǘ�TC���۸)��Ǹ7���� o������\�����~PPP ��u)Q��n��X:e���4Sᬬ,�4��Q�΋������e(y\j����N�!��b0��[�-�v#�]R��ᓝj�' ���Åʎ�� �6�C��a��l9K��R��U)r�og�̵�4	i2���re�w�[
��ζ=c)�;9�����c4�uNZ������'k���RN5�~n[T,���epBf����u���4{�^����G$iw�����>��[���ʶ�n����m���w��.<0��
��W�4R�c�ɋ���_!�M�Gd�Lc��Y��Y��c`s�=�X��qle)���wZIII��%ㆲ����'��M�q.5��4}{�����Jl�F��u��D���I "x�oaf̌�wseʇ���sX�������%��ag�:�rџ���l�����o:iv_���k��r���IԽޠRɄOPEezai)E>S1ۢv99����c����X�"��|��e,�2c0�f���e����Yx�?�@sBRH��J��e8� `P}��q�(�om���Pc�覥�CSQ��hv;�Z�wӗT��>�3���wo({y9U�`����Qf���A2�l��Y�G�o�*���Fi�����UK��M7åX2������mo����� MFTX� &F{���*>�mFfFF���NßP��x0k?�q���Y���m��%3�h�Gp������@]�.xL�x��7�v�R$��.��=�ϡn�I�ώN3�#"�����k�	Y�� ��Kg����AӖ�d�>���>d���=R�%�~j~F����!Z]�Ɉ�6����Tk1L�5yun&���՗XL�G���yTID`�V�8�rC�������������`�� ��g�ڄ���Q�(F�6���B�D1�ֽ\��lt����?sp����m���TB�5���#gj�a�F�0e�֚�*�.4 ��ڏ�Δ����0ܢ-�ۨ���.c���b��~����Cu>�͍�`�~���oopE�P���Ў���k���R�h���D�����:5���Ҫ�?op7�KKM�t�ɽ������:�!���~���.����r�ˉr����������.�ZD��[i?�xH�O;6)�U�_��Y���9��Q?�-�&d^��Z�m��k�oSs���S��mT�	�&�����
ƴƗ��/�C1�_n���<~�����W5= �n��ƅ^ofkj�z�82���v���K�N�C���QhR�`���j������rΣ�9�2�I,�~��V�b�_��eJa��8�mL���g�:�J������%�F�'y%^�Q�C`I���������E'(���u�;�2�F)�B
9��Xdh��<�ߪ��� q�?��7����J,��'���dI��.6B-��]�$J��ĥ�U�"��r����l�
��>�z>�bN�8*�2_�R�<�l�\��6ȴy�����$'&�4�B�q"�I��P�'�P&��<Qa#%�:O���B��G\��>Q��M���Z������!:�(9;�jS ��S��uꚚq���S1��ⱋ8���b�:��'���5��98dͺ��ͅ|iI������� ��H�2�۹8'.#� ʹ󘱷��{�l���"=�׻d�d�m���R+7�Y׹���)n��}�d=1d@�_E
��n<��xmt�@J2�E&�"@`v#�i�D��x����ţ��5�4���jVr2&JJ*��ϔ�MM�0X88k/:Ұ>v,��s�-��v�:�+;��<�&���zM����?�UNDM�ָ�լ���?2fVl�d!���B@�'�RiEyV���s��v����
g����:��߿5�O��DCCwiU�!�`Pa'8�P���*�=�2e�/�I��y̖)�̭�#���/�^������ ��б�-����������H,֛�F
vzpv�nXJ]v455eW4��+	�.5�����+ϐ�^��U������»�!''�΋Ծ�Y�1L��}�{�J�*
�~�y72���#ǈηe�����Q.�ui��1�>���-���N��ѣ�q}�����p���c�݀��("�"|�����aN���������Huo���E�6zA�C�U ��ZQQS������&*���і��1���\��7�|FN���';R���~K4��nP�O=� c1)&~��>R�9�<��|��/��e��?��(���L~�~��I����C���;����ȓO� �fhH>8jd���p~mC�@JSݷ,�'(�2Jh���_��e'������>�qf�������.�jA����������������=6S��a����D%.�喉[z�E����൚�o�:�@�`��b�o��)#<ƻU趞3��+w�w��%4H�e�^�֮��^Bp9>Y���k�y.�.�U˗SUU]�Z�����L�D��J@0��&�g��7�aH���+U%�ix
B�a3�Τ��"Z����o���|�{��(;�{�*#��H�o����$v*�.f(�jE`����+Ld1P��y-�7_:t�t�sE>������x�5��X#Sr��nq��J�gy p|6�_�7^9����Eƍʓ���o?U"�D��(x�M�A��]{���,�5y� �̕X����g����_|f�I-Ų?}��I��<���C2�#>�ߑm���C;�uw7�7=5�d��5 �޸��x��/�L-E��KĠ%
��C�W��NDD��X#�p��[�u�8�W��]��E��\~�c~t 9���ę��U�|��W�ٵ55�����i����4��01��j�i{(�o:��O��n�q�o6]�n��o�3�e��2�J�Ėt�� ht��]�3R�?ݹ3HmI������$eI�#0K�؝�����9�q�(c	;J��NM����,Bk%rc	J\F���w�顐 ?����w�m2-�X>|I��귝8�����F]~_��k��%%��#����I?�m7�2H��)c�O�b���1�gpb����v�2�wRq��
$�y�dr'&�$����6�N�L>�}�С�v�"|����$s���S7�6rûy�J�H h���B�)S=)�q��`��\� g!$4�	q#�%/�KA�L���2��t�RI(��$��Fde�=���Ϟ��m���k�U(bX_d��j�b����^9"�>U��x�'����_@>���e��UI��=����u�����W��p�_�դp��Eֹ�����r���Ŧp�B�kd^�n_,�T(0��Ј��i����zYQ$]WQ����F.�U���Sd�����e�0����i��Fœ�jM�Z�4F,b���C��ܨj@لy��yj��PJ�ş�j8��G-s�*b{6�6�m/;�{�/��*�I"�T1�e32��j"W�9��u�īM)��?P�J��޵  ���]���<�&Y�꯯&Oh�#dR���NwEi{�X|�(��}�]$��mQ,:[�����bR43�/�>a������C�%<\���}ˢ;��_L����0%��i|���G��&�̓iy]&�5�U�xAwy��S�>bP�q�ɖ�i���bcH(t�~�3��`4N3��W���_Pq�ڸz$1���%m��a�k��]�25�e���z��Q���umWŶm�Êm۶:NǶ�a;�ضm����Η}���_�����c�k�k]�7c�̑ݰ��ݷ�ʗ�������Wwx���	/�a���+@m�a�>Pʵ[j��������:��~>���򽉘� ����G���@�Bg`��p����A|��b�a��E�J��s�� 3�B+>�0>�� �,�n�=ۭ<��Т���VHPz�B�����y��Üi�À�A��9��aO9Uɱ�d����N�d��dOo1�E�YiH�Ť'EI�U��� mR�ƅ��M�����V���j�Φ�R�Ő�����ۥ�u;�((���������i7��I�NW�/Q܁}��J�FC0S)��J��#b߻����;��U����x��V�XdŒtm"cb�P�w+œ,&C,1����`���pV�
q�6��mr� �8��^`}��y����ܜ��oԲ���}��]�j��Ь������3S�MAk��`��dY��n2��O`��w7s���,Q>s��D<����VctXI��oȕ+��`
��@�����ɫ��2�Xf"�����\8�/|�H=�����+۬��s�c��^>-�Y��&i�����3U��8��}�h/��J�?e��M_7_�z�@GG?_-��7�:m����l����p E�e��3���r����6Z��!2�G`�i/P��z����?�%D�5�O{D�(�� �����IX-�ԓ%�'�,�O�C!��_��]K��\`���!��y�Ō�n���-,h���B��FUd@p,��"\�u-k���������=P���	���an�d��������H����d:G�����������=��vi!��4�����^����p߼2�f�K�Jb�J�v_U�����aIP�?
����::��W�����<4	�����"j(_����U!�@2^�d�����]RLk ���i��P�w}�)���9�x�:U�>m����Pz��D��3+���0�����"!�;%e�Ib�@��y�2��K��tOW��I�Z2o��DI��B���]��Z�a�:�a7��a���y�;	��n�`��!����k1ssh�_tex]���>���9==mx�h�E���m�<�O��^�?��lF���=#�8S����a[4�a�s�T���;�{�b���͎��_���� K�J4@B�@<:5��G��K��#&�s�����wVh�/"�gl����o<i��rL95
@[0R�H��8�	�v���Q��Ixs2����:|�ج�Q㩌�����Dp/$]3rpI$I����?P��98���:��4������C�A�NON��`�@��6ғ����欭�ك�����Л�@����%���d����n��U��Ϸj��PAZ�w!�Q$)&��N�&@Iz �S�Z2�z����*���u���犱�lZBR�K"aHB�k�B3�+WWHH��[�9m��1t�Q��j ���&T����e���(.���_��������76dP�{X�[��^�}/���C��F/ˢ>���v'4Tz���/}�����g�aA�K3-6c�=�j�-4	`�ט��Y��Ƚ/�WH���HG�H��Wт�ğ}M�K�;��"!@������D��R��y��q!�}ZP*54(�C(�o	A$���>6氲*�sd&
�%�t��U5'^Ġ'�q�g>�R��./e���q�W�����@(B��T�Tv��'D�w20�0j�T�y�p�/�#��dq��LO�Aq\t�^ϟnf�[)-�k�H��_��,��<h�BМc��ї6��\�s-4#10��:�V�HAWv�A��b��r`�Y�B3�{.�9�øz<�%��� ��L��M��®x������q#S�u;ո>�Ə���*�ܮ��<�'�D����C�Fez��
�%j����}'O$x^�L�4�=P/��|���¿}%�*%-m}�]����GM4!�6drF�ʩ�@�\Ǜ�����C�gTo�dxw�˙^'��"��گ5�"�s�����CGZ�(�~	���:�*X@�Jb��@⛇�
sj�I�������Αe�sx0� ��(���������z�6��pF̮� \��a�u�����β9;!�\6�H���(�饀�TV���&��RL��d�y�p�*�Ȋꮌ��O����у��"�v7�(|��,� ��h�������.>�!i��V�Ek������W�݋������$�~1-�
��:7��Ō �>ݾ�������|�i���X��O��	`�K��=!�����ɜ6�����jr��VN;<N������/N�Hh"E���F��a�Z�"6�;����&hIg aᄰw��nURY>T#��H[V��/*N�����%��ȴ�1W8ް���hS�0�n�W����F/�l|6�+���e�����6��]W���Ӥ=y3
��3��O�-]i��?�LH �iC�(���%���trF��t�ʉ��4��ᆌ��D����|�	~$�!�geb���wY����dn��e9S���:����ƌ'G��)�l�LU�ͅ
������xi�Y̸�H~L���Џ���6��b��YfR[,A^��&��A�
C NՋ3��b��q5�8���ZsO���z5���I�9	3��ʕ�R�>���֞�ͦ��C��Ś3�X���UIp�1��Ǥ��q���=_�$i��R�:��)���(���I(:�WR,>ZjO�g�:�n��P�P�z��)�v��ؔ%:'.�bi{H1p�c�������>��/�;�?�C�f��oq��kw��>Ul�ypp�x�LH2��%X�x'�">2�Lx�z�B����7�g�e\�vt�Y���#�j?)M|H*M��&A�l0!�t���w�D�y�r�J�������'��RŶxX�5f� i���#t�n�B!��
*�(]*Q�g�	�^��1t3'���h���Pɳ��)�K콈+/}��P{�l>��swI2�~�VbV�� ���q�2�3����H�i�#��#o��X���bmQѲ���G�*�r����(�fl{&�]���m��Y�w� ��*�Ė��y6�;$�߫)2����x*�;q1`IT�'�|md��wȟ����	�6�)��	�R�.��B()HiunjM�cS(oD�¦u��0-�У��^<�{����/�"��UH����|!6�-ꘗG�a���o��z_�����'hF��6u���cE��m�\
���k��ll�ww�s<v~��P�����"f~�}��`�?f��0?@O�:�=�)Iӧ�phw?h����������I��lY�g��� ��������q�y>����S^���3x��ﴰl�O;9<44%��"��'�I�ŕD�
�.2ң��~aDN{̜�+�bh��S犊�Cģ)�e��8
e��CA�d����B�.Uz����b�2N�6.�x�f�
.�/�xcj�=ҵ�[�F����*���
��p+�@��!�h��2��kF����¶|M�a�)�"���+9��)�z;�����Fz�/�� ��Ƒ��Y�J�n������Й�$��c{o�ʹ�K
HY_��2�K�һ4d0`�U�mQ)����L@�B�7��6�uWc3��\��UpaDJ����5�����`ƍAQo�uU��=藔��B�G�$d�zl�V����� �kN{�!v�Ie,R^{Ҡ-짟�	+XmPȿaN{li�w|=��Q�*�Javh��D�ە���ء��4v��icX<���������s2�IJBŕ`KKs�n�=���N)*,�p^x�B���
_����/0-+N8��B��s���ĐSv ��&U'k ��t4V�YR)%ˁ��.�j��=�)ɭ��M��Ii?�\��!���zb|`�Zɿ0KC,x}���'��� 2�1w+B�AٰY(�C�0Kf2"�u��E&	�S�N�p�x�|�+��H�"���6d��4C
28((?׍3��jFB̒`(����4܇��
�*	$$"�		@ ���aX��hT�|�ڵ0� �An+b!�*�`E�f.$����3�};U�D�15n6�/pيaޭ�29�&�B���;���T��d��9{�>�'�����r����I����m��X���I���mI��1�f���w�l}�y}w���`����S�6��j8+i�'?-��L^�����������rсI�r&&{R���@��>����_�xX��@aj"ңh���@<2B6�'Rǽ��k'��-������B������O���s\F�5��!��5�
�J��-��<H$�ߨ�]�ZLUFIhi����J�5X��;p�&��h�g�w���D�5�n\��=�񝷀�򶵏�N9S�c�dTq�3�H����ځ��o�g��j(�4*J'p*ayS,,�K]����ho�~?_�n'&:K�:�Z-;���u��{*�_�A����	�m89#Aђ{e�s��b�K�d�^k]i]��;����N�:	��X߮^JLՉ����'�	��R���{q��	zI���!�Q������V��
���N��ߖ�hf�Geuuu��p�h�FEz2Ի��֊f �N}ۡ�[��9*B�W�2T��mc4$IJ��*]l۞  ���;(�O͍�.��3��tB�ҥ7�>�l$�A���]�C9B�Q�v b�ڠu��7�ť?�k�%�����
�x���lAZ#��n��F����<xo�_�:`��~��G6��\7��|��s�~�d��qi*��*뜳��s�c��w��<�4/�O� ��7��A���nW;�K��fE��&c�U2y苁Q��H�d��VO���<'Q���nD7�8G��������`�_�����r8��U`
i��C@Y�Ґ�P6}��Ju*a��л�f����8o�)�
�ñ�y��,�<A�c�X�L�d���D9&�4�i��ΐ�
v��M��V���K`�{�H��.��l���g;~!�#`�_�)Cњ���{F��jz���V��Xk�g̊RjQk ��Tdj}������{�V�Z��y�;l���揚Κȡ9��R����$`U[�����~�<��P�!�F3�v����5Y��#s�h,Ivvv��*m�[�W��TDtϼ/�;å�Su��.�'3�+�����d�Z�^��x�I��k�}�����7FǹȒ.�x��]'#��G| �2���g0
sI�ؗb���*���Α�U,�AkIgF��,���ow���Hh������Կ��'(�ܻ�?�]�!���B+e~C�Qt������K%O�E��#�9��\lQh�h>f�CO��[/�:ꢭ���;�a���ir������a+A��V�2�s?�k1��^�����a*�9AO�کO�G�� �(�*��H����}���������l����<�A�*Uk[����4�l:hC�e]yq��ӥG�w��L��^��Ǧ��}l������� ����?������klll��(�-}I_��q�VK���D$7���r����I�����'����a
�x���XJ§n�ZZC�l�=�|�̧=#�v:H�E��  8@0��}&@��E����M�miب8�^�K3���J��\���HEN'��w0�_	���1�I�LN��W�Ww{*���G��&�O0|�pz�dn��+�Z�p �#]�yI��0ɺ\�_�й���tH��� ��]]���cl�Y��d0�sV@�E�{{�jE�|�*�����&�����7�4.�q�2m�I����+�����S�j��{���b?�u���k{��I�)�7ۿaC7��I[�@�@�(���&�x�8���"�k̈�>�sN�[���4�E6��s�H4TH��gA�ɖ�\_	0� =�sP�	���\_��W[�J	���Dg0�Q@�E�L�iǅ�1�U�x�6��u9����B�<�XZ��}�@WZ͐�r���u�A`)�]�h�zEW]~�1���u����i����rU{�-J��k �N |�W��b��$��5�6�A��R���ۢ��/W���~ش	����ˌH,����(#-�3�Y;<)��Z}��˸/���F��M���"�28����m(y�Uhg!�A���!H����~��Z�8]�O�J��0�ǌ���v�JP��B��7�9.��b����̨TR{��-������i�e�o,�o!��$K�_��o#L��S�%� �7����\Wcn=W� cmW/�&��v��`S�9Zn�zV\rSM����//b�8ѮZ������%�.C��ĮJ\ջɴ��o��9�^��V�s��'�� R#�W�NZ[e��L�.���Mxb�7��Qꜷ��܏�p�
�r�/�5����78n�~ &��@���vM���Swt��K�\֬��^�7>�d[kr���D^M]�J��y�~q�(%%��Q#�}��xF� 7M���Y��k�+�/�iր�:q-�ڈ�H*YʍoYJ�<G�"��� \F��r��}-
���洂��@��v82�y[I��Y�!��ROR��Y5���u�98Vǧ�(�KnF�<���,�����Jj鯺*�E ��m�ȵJ���4� �^����(��^��hc�e'��<��N�G���az�V�e����P�B�(�e�"T��P��`�߀Z��K];��1�\�2��1tZZ��2�?M�{Aw��<��_��6�~w���v u����:�X6*j`24�S��ss�?��O���gma�773��4�(.��.U��\S*�s�(��"g���(�[����S��\�F#�����\A�2��|��ZgǍ���*��;I���*9b�|�P**j���f\�c�1��}���2O�$tKv%-��8�E��F\��xI'g�QV`.>!�L��HQ�|gE<H �r�)D��+`�ͽU�j�_WRcQ���nź�
?W��/�&������
���l�]uv�6�ZO�����SQ�wz�D(��@�I��P��0~�2Omq
���k��Kɛ?S���c��X�
#���%��G� �E�����y�t�,^�Q�@�j9���d�U��Ӫ���4o�g�Ĕ���⳪��9u�XLz+{K����mn��'��L^��%аdZ�u"A��H�!�І��#��6rR��(�IO��Ȗ�:%��!�۝�"#z6{N���dK�ZU���I�ŧ>���q���(1U�bܮ�Z-�����J�&�>�FТ��3�/z�n���C�V
�f.�sz�_P}�Is�֧-9����9vo��cR��<_k��S����]yX�h!Ȓ�(n͒H�J���/4��p[�?�Y��0K�e����Z�HVv�0�L�QS*��t�`�2��Oǧ3wo<d���D���.�A���^^ �i���_���*�M�!�$p�=�~v����$��Fx�[mjg����������B;0����{f�)W�F Ifp��X|����^��`�B-���s&��u�ad��:B�$\ˎG |��Tۚ�( m�ԨD[���J���}�h���Ny�[� Rg��.����a��ꮏ��tC
��Ť�̈́��9���,�
喫�}e?o�n G�i��x�^��⽍Ξj����z�i%������D ��'�2���U"h,Έ #d������_��v�)�������p�[����n�ؾ3
 lN� gAN������7��Iޠ�!x={�eS�P[��8**�>%E�������cK�+��n�<� ���&V�� v��=H�d�&'��u�ب�{�2�g��t�s�2��nK�����)���Rw�A�+>~f\�qOd��Ī%��_��kB�#sE��'\�ar 1KR{Uϲ�d5ږ���hTX���2̉�w9i��}�BI��D�%S�?]�Vc��N��7�G
������(�	WH��������ݙ����$����v��㛊���4�lڬ�#{5[Nwe~�M����ڷ-ϒM�eyO��ġ����f���t�x���H�%���������y6�aQU��v+-�#��؈�C���1�'�,B�P�V�͍�]M/���vv1^�D��ʉ��N���b}�[w��舨	����-,'!1� s���i���aŦ4�G�E������������`������ό6�m~i����B~���}y�/߆����܅Q���v����n��X ���m�KQ�C$0�;=��;E�W�����~�K�Y-�Ԅ��Ic7Qʬ~�T�s$]��c?.�����������X�Yeuұ8���U!Ɲ���X'+��z�0=Y�զ6�u���f���`"���kdB�;h{(��/�ۭF�%I ]��!�8��}DKj�*����YC]�>^�<)���({��K	�(�h����������	��N�4M�,�A[��s���9L�� �̈[���qX<���qU���wg���wׁ*��$E�����{��Z^�����,p�O�d�&U�ϟ��8�g	;hn�_��S���VTw}��EE�B�&R�pQ�\ig��WN�J�)���|�&B3(�!̖r��ȸ�]�"��s:����Ee/4�/��ؓsb�+����H1 ̞��䢱Y�>�٤�J>uq�-Y�/�S硑���-G��ۨ��xI��]i��[~�����ޅ����$��ӎqA�5�8{�A�$v�6�f](�j];��M~saɵ��Ġ����]�V?<�Z����+#��d�[Ǻ�
$Ϡ[k��wQ����-��/�իJ:I��]dל�~AU��LzH��j�Μ>�'�<qm?��p�vZ����.��oJ����qD}��C�����5=5>��_o{�YtK1�����鮄cHzKFE��!�#G���.u��Q8���:Au�JW�X�=��t�����\��$S�]��-��������̌����T���Ӵwnf��m f�"�U���������k��<.��.�!"�;{�x~�]A��7R�S�$�oC��TEyD9 �p��<]�BI7����	���d�Y�X�/��Jd�	�{s���"2
�̹�p��!`�`TT4�frڣ)�K3㦨�d.�q#f���9�FPl��U��Z�v��i(EIQz��6a�{]�U��xW���(���/���x5�{y׶��Mt���/�m�$��8G!|�Y:	_Y[�(ڊY�ęV���8%���OJ��L�]��͈B�0v�0ՁM�@��\�
ڝ�boy�"��L���	'n�X
��u��gfT<x�Y=��=ШVLpT:�jJ�*:����7,x����a"�c����idI�-]���ھ#Q���]�����c�jkz�P:Ba���ET��i[h�J�_� ���pW¹�/ �b$R�vkz��ʊ&VWL+�
-
�����ʨ���X6�����_�#�wÉu�S�B��ՙii1���*.W�׿�|��d�%���+z�Z;����?󴀁��e�g�I��!BP�x0��d�:���N��{u��� y�j�K�2�n_��]�Z���>U�o�@�5h�'�B��v��9�r�զ��s7�#�Ďڀc���8p�q!���Ʌ�!� �3�S���qnͪG�󝹜�>��}�$~���X��*�����W�����_=�R�,��5���x��؋UJ��D�&��]�v����Mt��4ƌ�φ����5IԢ�Gƴ.��h&K��śu�T�l���H$��ث9wZD�	�QB��~��Ѭ7Y������ ��ǀ���ݏO�����ž����~��lA?7]�w#�A�@�����|���i��3Tw89@��d�_,�;P+��ǌ��ӻ���	�d+(aƓ���0wz�~Y��|�q=N�	�'�w9_���s�Do���5x޼u�D�c�7[��r;�XI�l'���ɨ����{f��yD(�.IƼI���d ��뢔������>�wYL�+��J#>]�#+n�8�
5���@��WT|�S�� !�;�B�4�����W.�l|�����~ր3�@�_����A� ��;`$H���b ]�����߇��`���늏"F�����)��k�q�XgS����X�a���� #+[��g�x9s�=���r�����w�
|i�S.����{���� �F�y�Q�頼9��j���K��/Uq�`.��l=F���ɵt��,쎗 �7�׬k��T��3����v��ܼ_�����������*/?���^
�AdHJ1|�y9���*.|�,�H�c��i�G~��N�Ҁ�(�e�Cs8�ݏ��y����`R�Ӂ��Ә/o����+*Nsj	�Aq"N�u
*b�a#�uG2��T��iֲ�f���֚LQ�r�Ր!��%"��$�ĥ*�
+��'w�ҭ��C$aO"
�Н2"����è�ϙ����ZNvp�ԧ�����5�e(k,�����k�TwF<�Zgl�ŧ}��"�k�"��xى���?��������3��B!�	�v�`��>_�&��J�������:A�eف�Uŀ��j�J	���F�I�G?c�a��6�����n����-�H����-���9�J)"�#��YFsԹd����B�EY�``����~���Gz\6�'aU�ðMep����}{��d��&�u΁�,��f�h
�D��
^���&�s��&{��6Ҍx�k��Par�� �J�+�"��&�Q�S����rBZ�(��S	e��J�]2�\}�;		̈R�JO�,]� ��!��J���2�Y�S��&��@�'VT}�nR��)��H�tܸ��aC���!����	i��5�w{ƆyP����n�<S$�I��C������w.���`}dΎ���ktŭ��E��2�Q���i�j�8�z���t�T63e�����g�;Λ��m��?�ҭJ���Z�[�ah�Ǖ����5�Ai�qXP��*��#�|i6�z�BǴ�"�
<�qm�ԯ�uO^4���.9�n��ޞ� CD�F����Շ�B<@���2/M���|�=ҍu�7aS�-�3��l���ކ7B"�'*������C����e�+SG��5�nL���Ku`>f^Ɛ�9 �.m�9����Ɓ�q�'�P�_�<�<@��
�=>((w�}�����|TS��d��ŝb�u����̬e4�L[p4�jV>}t�io�ʒ�𭌊J�AY'�(��ҳFXG��b��z�)%�Y��J��X�w��e�q�ʰz �ĭ��|�ˢI��g�]�ϟp�[��_X��/NR\x�Q+RM�O�8z��U��Yk�JJH��jL�,�#��qݶ���ކg�D,+������7��L��GlC����L�P�<$`Nw��r#�� 8�Z�Wj�/┃��pcB��B4���� ���$\'�
�9�D(��()��5�w�_�Q��wr�a� d8��pGV�Ě����V�%���&�Z@�����U ���L &-���	���F!/�3�@���\6y �jl����+t��P;���[��?��?��,�c.=
�2����n�@�$��&�ݾu^�������$�\@l�<~Q����Cʜ���J��DPLbu֨�S�:�� r�k[�P����Y�8 ʕW�������ɉ�������b��࠽���{952�2���FY�B\DY�>��8�]���wy�h*��M��W�Ca�̆����������/�k�:ݯ����?���V����5��\82f��"����#���Z�~)H2Y��LIeOZ&@���E���'&#�SFK��+<h��Nd�O�>(b����"	���<�rBR�ӱ�1��P�>�I��$F���#*9g6�414w|-��s�P<c3�n'j9��l��r~�#��H�0�EQ2+TԀ�m�/(�Z5��m|���|<��	��-�>v̪��EIK��l��k������t��ZN��� ��
0�MD�����|a�2T�D S1���!�@x�H�e2��&���R��X�o����ç���<�S΢B�����w��e)�f� �B��zG�]��ίyy~����m��O7ۿ�pɛu>ny�oy_Dc�z����Gz wo_�t�&���@�����Ci��;j����|a�p���J9����J2�8 P���ykd�N <� �6�DT�k���bج(OZ�,{xdT!C��e���Aw^��]�i��3Pa<��|H[oaN���	�����<�T��Y��PS[��EG�7�[~G��!"��*}Y�����=���8����Ӡ�	pE�����1(�v���f�.�m���FUu�ي%j_R�2H�����lW5E+�{�Li�"�Z7��g�P�"6/�CA�,>�� �E�_�<L��>��}q�A[��:N_�q\eĲ2_W	'�c�lىqj�1��"�\�e�58N�j1F��L�O�?���7�⎭�}�n@<�~D���ǴL�P2_qB$�
�`�|���a'���L�`�(˪iPNn"#%��A��Dw��*�ܨ�� @��*S�n� d�/�����S���~���+\� �/�y��y����$H�H����!�>��=� y�D<j:��ｺc�=g�B�ţ k�$���l��b�|�@��P������@��1Hk������a@IX_Qs�����k��x�7;�ҷu0���lh�я��ڿ��;Rl��J;�΄jM��"7�5�2��L&�����2N5���K�+�Q}۠v9d��T���II��L@��[�`�E�����o�����������ҞV,��V/R���F����
C�k&<\N�U�����~�Ǐg�1�K��8m��)�5|Z��XW�����4�cX- �)-C|N5�#?�_>�
c�ĝt6��1ë�)~����B�tf �7����W��OX��V�輼~���J�NP��=.�0x.���Y
�	�)����.�;6`�-�4���*M�����&�Q9R!|ܞ[��$N6��b0TC\��8� Y�O�4��`,���-j���-X�E�p��c7%7�Y���NY���<��������Q�����k���|��6��C��S�{�r��W��8=���	p��4{����L�$�R*���B@595%�jg{����,0��V�Ӆ�O=�	�@���1��P�R]�5T
x��@�{*��b(�<qd��y�������EH���u|���Ů�'�ˑ� 2ю�QI7�r�*y���;�� 8��f�"�����#Q����"��=�����ޏ���L��O��xxk�8����A�p�9�op�se�b� ���n)����t:z�n�l\"y �XN���<� <��nr�Ӕv	��Y��w��E��e����f�j{y���{��0[)�'v�%{ޗ���%��q(����vU�IL}o'��6ۊ���H��M����;40��?�U�Ŷ�0��:�B�ЄRtT��kl��|�v�e�B�00)�)����)��bb��7�`Fp�+�	�c.M��*�	�f���~K��-o7��oM���#Y��,�I���M�nfY� 	�D���M����Zy'��5;�vJʩ�	;�Mr�2e�	2㦺�����<�n�U�C��r0��Gb�b��1ųZ�U��<��;�e���B*�&a��Q�v��f�u��&G�����E�p��,��S���_�#j�^����e!�>��U�9_bL_~��Z�jF����ӡ���Oтf��Oc$nw��VKSڋ�:I��"]y�u�$�o7���lW��yJ�;3�G��n�zx/;�/R3�kdӘ$������U���(�S�[���h�T�Tz��٘,hv�����$���X �~ �c��|�e���x��j��!�!B��e^!B�_2pTLo�{�'���!����������w�����q��`ݭ���k���׉��[-��4)��H�������J��Z��5]��Ҫz��#�]	Ԟ !Z*eDX�.�6t���)	9�j�s� ��Úɒ��}#�8Zet1Yv��{�_z��8+JB��'�}���t4�N�7�?����>i�Q�d�$}a�D]��e�'�G�Ig��[�������(���ǎZ��t�r�X=^l�}@�~���Ӳ���ɟ?x@�3��n�W4�J�_'\
�O[��\�Ո�~[�_���� �x5'����*Y��#?2�
j��2LOb-+�^�~�Bz��D�mMvm���G5h�y8���1�
�b"=1i|JQtG��3�v�"Bz�����|3-�*�K =U�?,iC�-nZ;r���qQ��w�	A�0�q?�=�b�CC@�=b���G ~��� ��h�S!�uˑ�Q�OȸlOp畴锁2��3����a!�5 �\���ġ-g.w�T��X�0�DJ�Fw�k@��J�`���`"�+z>9��� ?T�� k$on�܍�g���t� ��^|�2�z4\S'�H�-�����ҁ,jk���>������yz���$�CF�����6��'�t�S~����0�	� *+դr��y�ۮ�f%�}KKk�H�%�j���٢�^�������L��:�q����肯�m��$Vr��f�rpdHG-��_sV��jwfwTn(;%���� #�P#xHm2Mw���d�y��v�,��w��F�)SC�{�+�%���MMX*;���/��4��^?ݵ�?t�͠��v�F�(��b��[�^:tb⯀����X+����~&)���3���sq���}����w�#����RO��q���h���W���W$��e0� J �1��#��X{cr0�Uõ�����J��&��
6B�@���4&;��ݯ5�<��&:��7IywFz+�Kw�
"j%ns=���GVxo����g�~��m�e�&V�Rj'b)Z���d�4c�8LFn���}C�e������+�?�0̬�p���ʅ�V����֦,�Rr��!��?���g34�	6c @�lh�סi�Y�|SR!#��R.Xݫ�F���GJ�dsޏ�|6����ý������9	�?�γ�
���A�%�tttT���R��Ș��S�A��b����t��U7��X�!����0γi֖Յ���?�ONwц�G |F���R�ޮ�_	۪' ��V��z�V�*��N~�$:]Vڢ��k��(������[�����A둈'��ݑ  1@���`'�E��C�;-� ��q!FA�8q�f����￯q?�<o��8���4�8�&F���Zu��WI�p��[�j�C!�\7�:��~��2�7�"���b�7`X�}{�����]2YP�=  xߎe�/)�,R$�%����f�b�mN��J��uiP��dYSc��U�/�}0PtP��B!���'�82�̟��
���t�/.�&!G����|��(u�Nc��ޠ,RT��>���x���`�#4��v��M
d�F���3�]�24$,^�3�nmees�J��X\�>F��J�sc$�I�[%2�q����㙼솶a� �_�w1�R��dkݙ�gb�6M�^cV�����4��f�*dhz����Sd�\绂�g��0i��W���?`�v������D*|���W��*�15�<'���B_Y�bǻNb�K�#��+�NLU�*�&�r>��|����ُ�+���zF�s�T}}ߋ�y��H�������\��M>s��� ��\�iRF`��E%\OM)}���m�~7_eϱ��
�����_��� ~;��2=��n��x
�0�ġ1?7�7is��s��F08(�m[�&�x��KB��%����b�T����G�W͠�b����d?��pЄ?��C�w��哺4��^�{��]�0���Eb{�V]���o���ib�E� vX�G�"M�/�ռL"9z$�.���=�;�n
,?IXL�:>2�e���p;��^��6 ���<|��C����hj��y�!�d���.�0�L���U	����ψ�"Y���333�d�_��.�%�|��p�{�oɻ��p����8�ˑ�����@�tv���*>�E*�=4W"��0߈NH��B��BԼ�9�#�3&E[F\H��S��M囁�ق�"o �㚹!Rg�GR>�Fz�q���	��}��k�o�V���M�D7�%l�i
�������ƪG�h�M�"�����"���t"��9tT2�t���w������/���J8��L}ePM���{p�`�����9�!������݂���=�sy������[5�=���L�*�87C�rR�s���IDb�\,iY��J�&�9���ŋ���+�Q/��y=UV�'B����^�?�e'�?3���q�n������C�jjXQk�����%q��d���Inv�۟�=m;>ֻ��u?�}�ny_�e񸾀uȧ�K�d�O�/UjV���ג��/՝�q�U�B��gi������-�ms�����
-��� �՟\�W]��# Bb�
�����y�u9��hY���Qj��j��2�p�H7�h �ܽ,׭�fu;���Y�̔�'C�J|�����`K{ޟ.�1�jx�\��0b����K�]��2�?����Tm	t���v�/Fl�O�w���ސ�)���A\[��n�&*�6<ޜ����*�8�Ñ��&���(Jaٜ���f�~�L=�W���Q5�+�4�b���!>*�˓WpV�DU@���8�QA���Bi�#�����YA}2�^2::K�A�X�8s-��H��|��y(���rO��a����~���cr���\�y�������x� �_ �C]Ex\�������"�,4��D�_q\�<�A"�z�����w�K��M�SH/���^�ρ���` {�qXb5�Q�VD������#V�*��5K�:�Lrj�|���Y�P�)�3�8RdN�r�/���-O�kc���c��OFcZE��O0�m�;!%��L����5.����;�Gko�=ޱ�J<A9�B%!�iVw^�^�b���l�֫E|�Y�$/y�/�+j'�9xQ�!��W�(�Gs�[�)YgN��[]U�É�d* fD��5[�.��I]:~�f�=��A��Dbl������lWSG���@��ȫo-rB�>�`��]@7�'������o'�L"f��`"���#�x�㦂�uLR�l�!�0T �����~����R��/
.X%��6�Y��7���0֛�W�=R?�K��W�Q�Ĝ��j���K��#��PCB�iK�7��u��J�S��<�%�d�7;;_���BC�)�C\��%��8��rr�4ʔ7{y5z���a0�Z�q��{E;��}��C�$v���{����1���#���{������:�r�E0�"̏^1䏰�A���1�GF�"yˆf����![��>�i��Y�ƥ��c
��Tj5T�'��:��2qq�=W���`&a,�W�"������ā���[����U��U�?�@'3y]��/�4/]�μ��M�]]a �*P(�iw$O��u�DZk�^t��y����~]�C�j>�?�\=>�b����oE��;c�7B��������g���AH��Ǘ����Le*���b�������w���Ï9��ΣlO"ǎN�Z�?��;��І;�TJCL�?���c���+
e_Hm�B*e���y� ��w�Le0 _����GR`�x�Pcs�`}:��U1�|�a)G�`���,���,(��9�c��Y�O'��-��Ԉ���!��(�.��)I��=�uS
Wl.��xx���Ef��UT�ᆻ��	|�]T��@���S����B��/7-'�֊m?����aYZE^]hZY��ͩ�j��h+ދ���ם>���,s����%�)�d�r��:C�DI��,���)���愆�:�x��.o;,Wq|\�P$����xn���dL�����2�{K��J�}�v�n��^��/��<���>&0S�����'��y�����W����Y���9!�U2m�\MS�j���|k��%2�>＊ �Tf8��C��UJ��?"U�2T�ϕ�W9y�S�4��`7���L�a�$�f���l>f�����
\�l�(�G�G�_X iqk���+ɱ��DD��K���l��"���=��-W�?{k^�8�DT׋9)d��Ɩ���O�Dd6�thT�0ӛ��tg�y2�Q�סbW�ry �f�z�0.Hc1�Sw�U55�@|�����Kw�xRK���L0[I��켔K��@�R�@e\� LJ_����&�J[{�9�+��.#�����צO��0dL�������r��"����Oߺӥ�E����Z��-'N�o+���ޡ�V�\�.���V�+�?�^5�}Vy�B��ۓ��nX��f�B��q9���ج�32g��|���[/�J�unn�p$:kp�� @�d�N�.�"����k���C��LC�� r�:f�Y(J��n&���d��ʩ��=��D_-Խ��	��h�j��:Ć�H �'˯� �$$����_��gG���I��A2t<�Ѹ�+j�~hNj��ġ\屘�N��<5rQ��&+�8�F�B�v2'i���b���R����ل�"���6�B�t:�a�^��T�	`�(� b�2C�g�Ht�[e����I��u0�:< �4=-��2Ī$1�zy6.9�����(����F�2��d���
?�M v��h�IrJ�/��M2��J̾1S�gr^$(�� �c!2I�`Hpo�+7����s�Z�^'��֏X��P���R�xO
��,k������x���)��er>�8�ڜ����rl�p�s?=?O���z5��e�h�4Ň�7U쩬RVxÞYuA
��g䨊8>ee�;F@�PZ�8�q��"��A!7�Դ����J��s��#��$Dɟ��9U||�8�)��@(�R}h�$��x�S콝����#�2]_ҳi��j�b���X�)�
�����JN��0�ʄ��$'���
ؼ̟�ZNkRn rh�3���j�Q(_���ʋˎ*=��9{�$�|���d8u���:n�s��&555S_� f�(e&(=�M����h51n�C�B�LV�q�q)��X���]�`��{���n�B
�TF��|1腥�D
�I��*������{D���*����������|���*���!,��/���0��L�JI9��U���q����½�����9���r���㺥�r�kB�7Y�}t+�^"��?��A<�ҁ��զ z��F�0�����$5�s�D�������^����֯o��!�0����"o#��a]A^&�.I�-��h��ZT����ɛK^6|�L�?�[����5��� ��G��*�I�<ʲ\������o���~��ݥ}^�$Y��U�|�!E�C�O�;�����7��|a�(c�`��ݝӭm��8��Jh�j?��n�%"�g�󭖫ö�<)�,-é!�����Z	�Ƴ��)�Qx�����J�w�$�}�B	�8�e'�ښ�]X����lE�(�Z���v����O���U�f�L�����,�O{y�X�B0N�Ó��?v�8�b�>췻\����9�	�%6��@L�/O���~��SQS#�v�����l���T	Z��� E��I��������f"y׾����u�B��ꋔ�S��r|�'�x]���|�����k�t롷yj<��_"��
���y���c��%)vLZ5�^=��@�|�R�`�\)_��CO�;Vq,�l�Y2���`4�<�z9���ɴ�Sm��0)\d�d��G�E�>]�6�PYd~�W!"K �Z*�V5�������(\,��8�^��Sr�X��>�U����	��AaSC���nL��Cˋ'Snê�
_ִכqt��4,쫩���-T[l��ƒ�l��̙NЧ�{�Z�w{Kp��I���촟ɐ�f⡲�/��*���Dڼ�4���\3Jv8�ʵ�v�����a���jE
���cUyy����p(����$�F_�`�a5��dh��y�zᚲB2�Z���ϳ�f@IҼ��a |�wc�ر�P9���p�F��p5��.ߍ�sVղ6��w�����������Pq��� �[l�/��!z؈M���½:����zo����_�����WO���k�D6��̆n���9��)W��^���T��"�������G(~G2=�? W�w�T�k���1���[���]�|�q�<1c�����F���*ܢ��ۚ�E1ؒr����� ���~��R�Lf��'��',U��閛°��?��e"&��{ PjE���V��ʐ��o4��P)I)� �(T(ґ����ۓ10r��~�ϙ>�'������ThT�F�b�ҵ~�a�;��|�--ۆ%����MAZdgs�%m�8�d�>12n���#�HFb}�s���h�S����|��9�{�vg��/q�3�ž��[���~�.Ot�&��C &�OT�����
�������-�~������Ƿ�q��j[�-��qp@��w��R��u+2��}�?o����n3L�kL|G�xQ�
I�`9�����Le����t�N�O�,��NXd���&�����<;�q\5@6���t���� �b0ğm���Ǔ�v[�"N]r��H�O\X ��w{Q�8������=>��C+ �B�;��.���R�m��Be\˗ st�CI(�s�w/~�p���<��0�R���8��&MS�pT߀}8*c��VG˴��3y�� �u�^�q����;	n�l��h�ܼ�!���o:�W�_����KS;yED���_��'t�����1j@�D�j�S8k�gi�W}8�=ݸ�Qِy���׺u\�H4:;��\T�iQ�ﭮ��_(��z���,�7�k~Z���m�I��t�_af��Y��Hm�w�b��o���ܓ��W���~3���e�N(S�����|����g"��g�f("E����Wrb\���j�3�i���� 2~!}�/���H�<=���=1}�MM��!�D��p���5&���ɈC=~F�3�X˯M���e/�/�_I�Q�R&ډ+�$�}0�ϊ�BaY��<'!{fߐ��+�_���C
4f��5�5wCX5��T2��Ƙ�_(�T�cyU�#��sƈ�9���͢i�����O�AEb��*�7��G
M���:�K���>�g׊�)�pR�jW{:���'^9�fS���c]��5���OE�$JW�z&p��0���uD�u�7�������C����ǎ����0��U�~��ؐ���u��#�x�2���ؼ��=Ϗ����V`UY��*U�@�4�M��FS(����C%�0A�N��[\���-��*���&7�L��O�f%�3��o���M#?{!&���77;��#�σ,�7S�K<j�ƃ[��N�+|��Wj�7��,C�� �ï���gvsNE!\Mg���A��BE5���Hn��,��{>�Ւk�Z꿝H�K(��+�O s@����U�
	F�1�6��A����?67������k��.�*�a<[���������h�Q�AAe�	��]��ZJ��,ߏ��NK�3��}ˌY���7�㖰������%��lT�)��***�/a)	˛E>P��e1\N4��˘�clF���� ��y�����o���(�9U���B���dY� �1.�?^���o�.M�2,���.잝�7М2�0��:���?,a;[����pR���l�i���nc6��7a#������t�9����Q�����v��}�h�C��f%ߢӍ������h��<K���(�"4|���5�[~�Be{݌}L|��455�j�h@@ 9p8��_����6W�P�FK���oyU��N�H>�ᐈAv�L��U��ro�e�J��\uF�v������"_�\Aw���E��Ze-E�hNc,Px����."���H���6c(������#��?Eha-|+,����' ��5�Qh9/6 Z�"��Pw�C�-<�����S ~*�4�d��0���bt.�a��sÓ�����6=�ou'�a�U�7�5�-aX��T�s��� Hd]6����b������j����3���y;���|A�O�6�h�DrU,��"����׽`*�c�6%��M�*P���!��݄�Z����I q�Oɼ��n�a����[Z�0�����d��X�,����l����$vPW��A���2W�xpc�:��������J_ �]���V�����m��w<�{���Z=�[-�w �=4Lq[M=����<��gHf`Xo5y��iF����c��uQ�zu��A8R{�22N�	��cfV�""Ϝ7}������C?LjD���?k<�q�d"��{��=��W93j6��<�a��HEy��K�=:�WN��F��H5��~�����<j�H>���;O�dY/�/��_�:�Eߙ�Ԍ)%ev�$Y9���{�t�Y�`s���a`T������~ȸ�L&-��j#zTO�]N�_-�ɤ�i���ϿS�f�Hx�+�CCbպ>��mF�_)//_2?_oJ#5m�]J
~�G�_jl��>\8^4���͏�yI�P0ɇ�py�P6o����aɉO�~xb�����.<!��e�:���9gK�#ʴc�h;�����K����wc�J�"�!��wi�ˇ�����2�س����`x��&Â������,0r���+����c��Jd�����������mdp̷�]����{��y׶�T���o:b�ْw���ߌ���Y�����E�tQ��8Rp����ec]5��ڐ�X�.�T�uKrf��pHj��ã�ɰ�!�N25�,l�����p����ȿw��^4�ځ{�っ�;���(	mT
���tU�[o���k�G���8�L(�)G��A���e��W�]n���r�ݗ����\��X5���m�,JF�䴏nL���HGh=�;2զu��:��f�X��eϕ��75�	0�S=��}HJ��k��gjj�$�B�E��0c��՟gεv�� ��m&y������� 95����q/�E�9T��L�lB�4�	k2�/���\�|���n�7��<�K�����+�ɚ�M��=������ik�����~��v�k�����:Ǧ�m����������.)qR����T����m/�S"���~���_����ښV=7/�o~ff����.d�(f���r��07i�"k�?�k�`jvy4]=�_u�@��F�PF���~C$�OF{8�ƒ,:�[��-�Z��B�Wp@�^Z[79 �b��ۻ��].��D�SJ���BvSj}�	���d�{�^D�q��+�(䱏r�+�����[W�$~�V���+����r�Mca(q ��vL�U�p�oTU�a'��󒴈�"^��L^�.�լ�	�6���̕�{V�g��-�J���X�K��r�4$��~�*�¼'�b�hM��O08E� ��~������α+y��F�P�  ;B�PفQ���.�� �9`���1�2R�9�1G�cs�������T���uu݆GS��?���w�*�$�ݦ?��h�p$��������x!L�g;��:l ���	����Ҧ��>�����	�`��'ׂ%,�\v\���L�,��e�l��j�t�`�����.��J��j�{m9_\�w��v��/H�@��[L��2��2>�qqqɛ>�������ia�D`�0�4h�^܁��n6���J�F�(9��8�����R2�!Y��e���μ��G��sZd���EQQ�������@�_".��S"��#k����^t^�����W<<<�=����ݖ�����>=���0A�����z�)]��P�b� ��,�����~����T�-2M���ӟ�ӵi�����8ts�$EX��&Y���ssr.{A�a�;&�y*�¤o	
�G�X�QQ��>���;�(]���c�7Y���<1�W�H�5#�@J��>o۸q���2�>~����4���倌|nhd�[�貚��fR �qq��"JDˑkǪ��B���f�8A ��Ph7F@�� }�(9���A��b�xw������ v|>�f�[X���9U15r�Y�� <�z{�� R�w�o#���.�� H���f1En����.���Ѳ��+xѱ%c�W&�4�".��/M�4�ǲ�۬7v��(	?R�u��4u}��>^�[l�ڋ����tw��mu�S��ص�/*a͈<��F|�&��al��7S�Lx�G�#�xw�W���f�o����JW��iqS�N��ml[6�t�k>�?�c̐�n=\�q��E0��� c�xeR�mo�37�7���`t�A�����l��ܖ ��޿t�R�rv�����j�磞�� Z�Pu�ݸ@y�~�m����7�� �$i�N}����&�&��e���Ɛv���&�ev�"e(999���{r666��`EF�(̅�%LvV���;s�?�Y�>H!���+7��ϗ�5��
N������'����)#6mY�<)WĂ��ť�/7Y�9~�? �3�{Ǩ��B�L%�[ �e�<;i<�a���Hy(mi���yޞt'�6A^X3�E�iԻ�;�״$�J=gi�P�9����}iH�����汩����������͙k�f�N)�x_z��q�F�bT�
��T��<��nU�afz�B�}�H�t
�v�~E��HV���~H#��G�K}`EK�Zޱ@����H
�;�^㶚X�s|�I�����z����΅Ldbeǽ��$|�Y�Lo#���+9�89 ى����HF�(CQ�.�r�ә�����:P��� ����wu�y9���8�c�I�"��$��l�L����	�?2�5������H"O�Ct���������N rO��l�O�=����2�����{��9yD�ӅK�Eϲ�^�Ǵ3 �+�݊T�n��_��Z#�!��C�&����>Qf}���~+�L����4��Y0��8���o�)�?pѨ�NSZ��2���q�(Φ*�0u)*6_ae��%��e� �3QTAejo�=u�`��5 o\;��U�ЗLl~L���!��g �VSS�cI�u��~�|����O�X���m ����p��yZ&q�}Fx��~�����5������T�<H?�{>�/̦r>3%���8{̦���ɶ*�l�v���T��5Y�?�u�ƌ�o�̚7������t��i+���L�O���XZZz��՜`"J&ܘV&n8����>	Q$�^�-\����Qi���9ľ�U"d�~J�\@%�ӥ�����p�q�X�T>�x̹EZ�^�k��vrbt��?ӽEY���� �y�K���-W��Y����s��Eٕ0\��;zj\�@\�8[&�F�e�'x���^�i�C`ڳ�, ������Z9.NX}���I�-A-I�%W9�P]�z�ߊ�-z�b��N��sQ-'�y��LLXT�[
 &����!�"��zǬH�*n�ssܩ�q��$��8�y����ݱ���Z�r��bb�KSYM�?0���>���ߓ����FG"-p9j��ö%�2��B��ie8���c�x&����e�(+S��3��V��W�q�R�"�Q�?�i?��s2�b�u+~���t��W�5Es�
���)-+�eN�����-�g�ǯ�(c�5�Eh/9��\�〽�S�Q@��T߂���l�o���z�#;4��*�w�]���n{�-a�I]̶d$C���wcњ4��I"��wN��=YnY3f��]7�-�ׇ��IW��H��EW�c|�&^[K}^ n:��ƅ�-w,=�H_�>�x[^6CF���X��+5Û�U�k*�Wv�b�@.5ZmD<\��d�R��8��s�g���̯��1� �</������	9�vX(�������/���|ۏ�y�f+�G����*��"||vk�?.����˜;�Ql׫7�)s�
�VK�m;?��>ߎ8.e�U��;���b�_F��#Q1�dR~g�>�P&�u�k/`�9�͗(l��yf}���󟞝���w^��N��&�u�R)+�I��� E����:"����M� e����#9�!F*GnM�"c\���)Z6gΊ)�`�+��#�c�Dv�Ȟ�2R�\Ǘ�̒�@L�ǵ�I�@���z�Sv�×@s�a�?.̺��w]�R�5�A�����Aj���5�O|���Nl������p��O�S[�i���Z����!������_i��f����F�#��_<��ݴ2��\���"m�D���Ҡ�^�d�h/vFݾ��٧J}�,��眑�D�9��]`4q���E���Y�☦�J.M`� �T�ӟ/�2Kg~�Ōx���c�'��S����/�E��̈́�	��g2�6����=������iO/S�{h莑���Io��0�)����t�v�MK�Ҿ�~'��E�U̲ܪ�Z�ÌL��M�%$,���'�Z�J)N��2u�ѽ�����:��
�\�l��{]���t�WȻ�F��U�Q�!f�e����>$�2�
�=b>*8�%ꖬ��{ޒ��t�s%�j)��ts�^�A��FX��6�<�7��S��r�,�,����>�����v��ؽ��R�Uo>=��|ZE&��Ϩ`z��m!�����B ��>4���Gp���?��D���S�m�T8KH�������[��rѲ��H㣅D�s,�&��Wԅ��[0b�Eݫ��ժ�Ai>gWW�զ�tXo{
5Z()�j�<�'�O_�y
E}��3���㨨+sh%;@q�t�H���2��e���D �|��<+.���~�b��zp���YeXO��ٰۡ�����%6���b�¶�Ht�|�y}$u��C[�����x~�\n�Q���2�4/(1<<�35�����L��� o�>rZ\^��G
!ˠ�GQ�v��U�r�>�-z��=l�D	�k�y12�I�/]���|0G��OT���!Z��@L� M� g� �;U8O�=*��$_�y�:�%]ć���9�k�K�2r���&�|�8R����d�/&^s�F��y��jK>�� �h�qU����=��a��Va�i��6�*!�QF�8Rv1�c/�7KF�����{�Rz�	-o��ǎ9'��r�Hq5�|kk���J�]�܏��U,�:�&Nf�Z��hŠ#�nn�x���D�]�E�>��,n5H�a��kkG&�kC��PKf�$-n��c��)�rOb���4U�t��#Xt���z�C��J��Q���n�~yAQhF�����3�ψ= G��ci:**"H?,�)�a����G����Y��7�V���$E�Ң&Q�v�*E��y���*z�P��V���q@�r:�������L�F�Sj[�m�>�]�[W�/�v�P�Ľ<Q%$�����a���ڣ���\<�<VD��v-f��#Aq�}����T��^#��-E� �.mﲹ�.0]u�^�Y-U�F �`յE.��`���b�8�o��*M��4���8�=�� ���:Ler�peM��ˌ����`'��rD��|7�"
�ȅ�}��.����1I_���M����(F�^b$����ˈ4O���f�k�M�N�Z0l:a,h���w�����b`��Pl�Q��Y26���U�D��K$˰ ^��8�)���Zs���������?2��w�����Hs�+��?r�_�.\7|N+����n"^}��Sa�#Y��|�'A�m^O���E��"n�:׹sEQ��v;�ǻD��Q��k�7�؂�t�5�k�^	8����w�?[l�1�8ao�(b�+Nr0
������1bhK�v?Z4�)��A�voΩ�,C�goA�fI&*?��A��NKs!��	�䙧�H���3Y���!2�P�LOr֊���Ĳ�"�-9��A������1a�*Rʫ:�~�4�-���8� i,Q�$��/���/�N"�Qse��q;N����?p��.�{�O��*��9e7�_�p��<{uY���U�ܐCUXɋp�B��bUE�*����L��`]�q%��,��n��0���J�X���\}���I!��N���T��Γ��mG-v�$��d���:�lCE�7�P�(�#uu��̯��t�ЇF)ngƿc����C�����FSO�W>%�SŌ�,dǣ�[�i���7�A�g��i'�M�[��=�4��O�e�RB5���Vl<�����y��7T��PJ#x[Q3�~dJ��_0O3d����]?��L�1�(BI�]�kT��]��Jx����Q���C���%:[vk��B��ai��6p�����^9��⁔�s�%��MW�wS��e62 ̾V�5'0Z:}�&W�P3<�0���$��H:�ڄ�of�\�eca���Z���L>�bD�iC���}y8s=�@�����Q&�˻�Q{5V���	�K+*��}�4h�yu�5�J�>�
A���(���tg�K����(�A����gL�54�eL��C�6Z7��z����'f�,8�A�u���F�$㓺���1۾�7Z�o���|;�i�|�H��=��b6�2t;-��U�v���@漽s�~2�w5����f9���r��; �>�e
�������#T��e<G�-�Y��F"�Y$��9�{ݎ'�s'���<�L�GF;�<)ir�PQ�>y�r}�v
���ޗ�Y�E��W�@\�ւ٬���T�4w<\Ҡ�/i)jD��40[�I����5��k׾�*)�$A�1I�2� �-Hqq]�"�3�/����e�A0��_X�k������a�Ģ��76i<)�q�������5�l*�s`T�V��e�ej'�W0��i�l �e��W��ғN�d�ӽG�H�X���+	�4���Λ����T=���c�4�/BY� &c��x�P�:��D�^3�3�A��ppm:�P�B�P(T��4 l!����ו6�
�|����8�6Q�y^�����ru�2�<��%�TXj��^��0�r҃"�]_��� ‷�l�R{L	�<i=U4q9S������'������ݞbݳ�fw�yN��f�wmt\68&mT���u� G�3�<ۥ@�_����J�
|���v�����b�XZ�&�.����g6�۲5�  ����B�|�I�T{fgT�办T61���E��i����1�Պ���������p���9\��&���lb��xrc���b ��r�*��}��l�u1��I�Ȯ���5���?��'b�k�|_��*�_���6��̲^�D����F�F4�u���ہ 2���A����J��Fx-���r��!UB���BF��Ńgcc5���M�4������t-"��ۮ�����{_�9$�ź������a��,��VΝ8o��d:�k�e9\M��l8��<��lj�T{�d B'�� z��z�������'�-p�F�~:��ö�2�F	�5���� �;s���w��C1П��y��V2W�Ư85y���v*@�<��G~*�iC���D�Lu&=�s��ɜ���#�<��J��f@H�����-ϫ���IN���h��ƿ��28�̟a);}�O?�O�0������M���v� �.�_m5[~[�}�,�4kҲ�_݅l(��C��7!s_�*�m]*46��n�w9 <}?��/�[__C��%$�����_^^����x��WV4�E�ENC�\:U����rEs���Yr?��,���co�Ji��"���!e��.�p�\a�ԡ�͌�����6k�<m�=�m��������X���G�I.8�GG��+�B��(BݻS�_��Y��
����&#d��cB�������G�!�˛!d���3��7��^1ګ������qua%m�b�
ހ��0��.���ު���c<���^���zWU�q��O�~�\]l�C�O�G_1{|��N�>v�b�i���q^.���Cf����X
��@�2}֠���H��|�-)w��J��l>�-���3��$f0��󮗡�M�#uw$����Tg���,���M��z21u�X&F��k���.w��Oo��q ��0«�kzP5�ZZx�Q� lmb~J8s�z��`5]r��Q���QI��[�q���˜��ﻮϻ-�<�!���[����}*Ͷ�ɷG�+SL��8��96� DkU�>���O��x^���<���,����x�Y��-"���/Н�1Ƙ4Lf�D�uO%�F�e������/|^/8��!q�??��u�����ܓK��{)x5;�Qg� �ya��|���ַ>E�%�;�A�����p >�����
���+�&,L%e<�l��I��l�!M���0De��p�ѳ�na�(G���Kˈ9�X�Ia��ǥ�ۘ0y�9ї�=�[9�b:*#��<�7���dZ�o:݁#��-�3�\�16�q���TVG�ru����v�Ru�<:t,�����&�W}����7����嫄$9�Rڢ���������{A>0hX%�R&XFlB� H�U��鞜7O\ȟ�����g����j��`Z3��ׄ�0�ǆ�eX/�/4�*"��>� b� w�v&�@��6#6�ܐCv����֜vP���a��[#����+nj(��)���;:�|�ߊ���,�����f(H�P���+>Z���h���\�Ξ��+֥�L�/�v�v�-��Z}���<���xR���r�$|�U}��7�,0,˓7Q��Fw8���.��t�ZiAm���Q��%!p�TY��l'�ڶ��AS�e6x��Qa��2��nrf\�Qz�t��p�ә��lM���Ɵ�+C�s��(���=B�e�z�Hwot_���e��<v��r6h�ԗ�H3G~B���a����f�D�4#&nS p		���l�G���G�e��e���er��嘘�nT���k�Ă�3��j)�He�/�3}�k�����BC� ������χӕ2�};i+@�;��V�"�(�J#R�Õ�χ�[~��}�.����2u]fn���Һ:�b;^n|���_(b*'ش�o6^ٓp��sB��ΣMϕb`c�,����^\��! )`��z9v�n��A.,^qVy�^Ƿ����2t�'NYQV9MU�me�TD��*81�G�,��~��Qg}� s�V��Ia�6G>-R��Z��$�E%Y����(�
:P(�����b~7|W��[��	�L u?]�~s���e����|�hf�}�dG�?�p����Mߓd�<%�WIAj���Nv@qR��O%��������}ā���JKG���y�Bᆺ �a��X�r�/'���]�*�(���!��H4�2��Rc��L_��5�^2O"�tё�~��~�x�������V`�O0@�5�Gv&��^�Z2��(#a!�Is����Z����0٠ �Ag�Պ<	)��Ve��3���n�E��b��2��_�Xl?��K�[����j��Lt\΢[�G�H}�Щ#�ԣ�bK7���
e�!�����p�hD=���J��U�;��¨�XШ ƈ�C4��I���c-2#��f�}�d�?�Y ���i2`���i�Ƭґ249$(�D���/ҍ!2��=?;k�m�/��F�)��?ކɹ&p���y���c��L�pt�v����2����%D�Ss��jCf��JDB^�{"x�cɱ�N����7`x>�������y|�I�q�O�x��6���N��p���&,�+�,w�y�� T`���g��u[e�é�a�)�}�8!���vr��ۙ5M#���g��`��W��p6���I�F/OnyV�����jK���}u}�.�=4�</)�dp�(���Е�y��M0F������V�	�����	B}�0C�uZĺ�C��L��S��|�4J����BM�<���D0�u=�jb����Mj�p�F���f[�%�A ���lP�:mJ�\�J�����l��5�u��N�J՛ſ�d�2 �D�Dv�>����/�Nr��Eǐ��25u~i,m��h��V!�i�cL0S����-�Ae-�����B�~�TXmW��.-zߠ��Y��e(����tu��B�%���w�d��?LZm�* '���U�BٻH��; �v{��f�W�ᨨI؀��E��]��U�>EP�PJqp���=]������@���ռf�1d��d�W�Vp�����b������w��X0�M�i��)H����$���&:�Inp�QFE6)?ȑx=�JK��bO�m�&#7�A���I]��Րn4����xbV-l����~x�;'��7�53~�9���Td�xTޡ9r�Q�#=jew�G�KY?��=RH\+ŋ�)l�TÌV�Y�G�#����zx�Z����^#O�(Jd�]�:;D	[E��LOX���q�L�٬��R���n��f	,䇞?�@��dC͐��m���Ċ�c@�F��b��%C�2J��4"p�R���B��n�6���>�m��~�
&mJF�7��'+��,&��-�����|��ӤQ�#��D@�����?���GV�#n<7�s�`̝;ߞݶ�4�,��G�X��.���^��פ�}�ݗپu���CC����9cڔ�L&�X�V�
�|5�(��yK&	�K���,�pF�(U���j���D��+�L�ZMU�<�J�t<��\�V��J)K�&K�+�3�ؤ��E�\�l-��#w�s�V�=��deT\��mlEqI�1�D��`	���Nd �~�@xa�XH�$r�уx�����kAV�Ae�5\YxZ�,u�	����`��rZ��OzeA뺜׷}[4<0hE_j��T,{���bKx��H�%-��M�V���)�ɖ�����w)'ц�|<�\8�7�ֆD��sow�B�e&A�@���x��P�Ld�qm���(ݕ�s���&�הZ 2��W��*C�9<O�� �u��7X��C�]WJ�>ҵm����m�~�`�1ߕ�(@ӡ���ݭ����''�.���N�3'Ė�L�LL����Pٙ?�Us���N�:��\�"C(���z��b>�NY��]�9¼c��&ܰ~�����x��H�*k�{b��i7�18�����,V��Y�X�\����K����j�y"X����Z�����!�4�&�F̆�R�fUc����ѽ�W�N�ʗ�X��$�'<����P��Z(�3H*�q�Q���7k
�j(?Š(��*��*����i�݈oz��c )Ì�����hc��ڸF+�a����D�u����^���dr{GG��?��O^r�Ǯ��������^{�;�<������g�<n�T��3V�j�2��hi��|;�ܶx��ξ��O���h���\p܏���׬yv��|�����6���@�Z<S25�6?��s?z�QG�vAG[��G>��~��66<83��d[zH��n졶�n5����l���r�9>|ɂ$�bL��B�~�Z�YEV�䈺TݏF�y�/<�EI�Uƕw!�"��,$	)YYL(����6��FB�LX��y,��\���6���|��,��#�������LD�1,�u4N��F�����5Ȑ�6�v�3E<6f@VGa�R�d��#a�8�i�r�����	. T.w���pM1��3tWȒ�У!k$��=�̞mm�����\j,Rzq���X�7 �8ĩ�R6V�$K�����`��A���@�����|� ��n&B �3 �cYna&�ÅVݕ�ݎ ��0T(�ͼC�YU­d�8��x!`'�|��pZ�ڊ�)xI�	�MTj�e
h���q>֢ ���	����缳#|vE�������n�C�'����z�tc�u�z�f(�B=��<,x:+̖��]m@���.���!� ���=Tx$�u�e�a.��%!��9��x�p6��,��wp奶��B��o
���XS�h�>�Ok�]��>�EcY4�d��S	���O����5����M�g�<�kĴ�Έ^�%�����s����-���L ��� s7 )j�q<��{�Ⱦcl��QB���%K�.{��N�{����+��k�o�uǯ�4y���߼���W�~��?p�	�F�2���J{'��y�!����=�d���ϟ��K.���Z�/⋛o�y�W���_�j�U�$���r�a����?n1?�+[�h��]����ne c�ƍ�o��U)Q����5z�_���S\(5|���~k��B�;��B+G �A"��;3Y�R�l�\,y��ŗ~3��o� 1��rC���9O�`P28��� �K��T��I�5�֤ѵ䯗eC�2!m��R� Kq�`�	�������(����L������}���li��"�F�����\$�6�,H�MC�ٙ��/Γ�5�DlX���R �-�bѢ���"������9^�B>T���6�"�M�4�|R�cHǆkL$Hi�	��P�H��{���S�Ł��%}�ϥ�5.���o��3��1;�w;[�aN>߁�Ĳړ�	?���6�
��Ϭ��9�;sO�ya�-o��a���IO5������`eHp!�אE�[L헂�5m`���D�F�v��q����>ge�����w�$��BKdx �6m�ʒ(%�#�pZp��E� zjJ��b������㼲5������Cv,�1��hr�N��i��@�TT.zIm�K�&a!K+ �O�Vp�q�7&e0�(q��$T<CE�_e���c�3ӐE��K�����_F��,��y��1�\W�� ��
r�#wPȨ!c��"���k���Q���U/��۰� �b��Iމ����8��Rd���4���x�g?��O<��뮻n׋/��[�|�w���M�.��q���W7�=|�������lj�!��������/O�֡�>������[o{�E��.z�$�nB��uR:j�h���w���'.�m91��*���kN��o���996<by�=�-Pk ���-h�TI�`(�~L�:�d��k#N�7���U@Ȭ�T"*Sf7��吡�����lW�B!����%��(� ���b�b�3�W�WJ��H{��E׆q���uM&4� �� a�] ��У�e��B���dE��R��J�7@
�B4q�T��^�B
S����B�	�88�>2�y!Y�����v��\���z�٧p�d�)hU�E��8F�Pћ �]<�ߐ���\�&2�D�e��Ȫ�:�:F���bA�.������>=�~>�
�)��w������������ޝ����"�)�5y�$T�%��:F��)3>1(}�3}�P���h��/&��B2��V���Je�Z�$��p2��d��R�X�76�45wtu���c��֖}6nܸ�;�kB�|�9���@M�Z��)��[���a���UsiP4�g�z���G
)B��N�#	�#��ì�a/�$:<Cp^��W�����@��U����k}�[�c�ю���O�K�������NZ�?,��j�����}&bW����O�(sE�nf(Z��\S��@��%X_��u��GfI6غ���Be���c�����'e���Rc!0ó�������y�8�L�c�#15���I`'��dhd���nʔ����|�!�s�:�:���o\��%K���b�(:�~�]�9/�HE����۱�ߞ��U�Z�0/����H��)������?�|����y���9���֭[���3fڳ �q��X�"�{3��|n�U����~���;�s�d���|dp��ӧN��FG�]�ω�8㌨Z.�hQ�hhk�"���J��c��p0��G��w!Ȉ����	�X���&lwC���@F1:����R9��qMȗ�T+���BNQ�N�r��-�NR��и�%VאxPT�Ѯ��MV����mv/ ����L�d��/�1�W����.f��{W��-a��Yh�P�
6�����i`7I�^�	_�Y]i�9��V4������N����h'm�ri
�s�y�/�EV�E�����S�x	 Yi&����o�B��������&��3@0Y�K���� ` �I;wR����	����L�6jLCp�k��SB��c�g�w7��'�ɱl6;�N��Qu�%F��:�J�G�#m-m=M-M���;�7�����ڶ����L�6�0u���S�����&���u�?8����p����?��H�[� 5?,�l�8�D�3��/��Ր�=N կ�=��
`�^��6l��$z�	�&��h��|�c-��!X�AD#��ِ�PB���7 �����S9�X���T)�]0|��q��L���E�+�%@H?(�A���uƩ}��??�0Ͻ���^k�b�u!�y -Z��E��ǲ�b��yi�4�5ZW�-����}�xq���!H�nW����9�#�"��N0/<@�*&[��6�7��Y7��\��K �\�1P��޳�!�p�����|���P��_��������-����T*��a�-1�#�ĀE�y�*<�@�͵\ƞ�\.���'��oy׻����R�/�/|�G\��}���w6s���= 2�1�d)nٲ���c���v[��|�۵��~'�x�9�����qx{ks��d���fG�s�����x4Za,油&���c5�M���rD�P��g�%�Pڗ�u� 4���� 80�Dі�=ѻ�uN4R��-�	�Q���)Ċ[�ࠈ� �Z#����곔��-�d��g1��,<~�~�%��X1�e
.]������B��k�$s��0Z���+ȷ���uV��j���Z R�*�%�2��|����o�����ch!K�	 H��8���8�1Ƅ6mڰq�"a!a%�$�����ٙ��w$R�R�j�x�E�\ C²6��쇝)�}����\�!l�ͫ���-��_ֿ��u��n*���es뒩�p5J��t!ߘI%��[��NY��Ҳ~֬�[[�����;�M�]�F����lv|ٲe�__��K���;�w��M�J�s3�>�E�m����y��;�v9 c�y�@nn��ƙ9�y���6?�CL�Q�Io�v��nI����,�&��a������Ĕ >Xg(�[)S�g�G#����"C���}�o�h�G����n���a�/��ӸRqXkDl"�B� ���'AaE+�řOg�m�����/�Ř�R�.1��O#9"&�1H�|�/��������C��4�3�����s�_,�g_l����.ne��\-�;{���l�?c���L�Ĉ�;���N��l�:88������ꫯ�P'���O~�ӧ<����388x�����g�q<6n�زbn�p�(�U��gm�_�1ܷ���G�����w<��Z�O����~p������%�n����F��gk�>sw�=v�o��N;�Z��j�Qg����.�s�%�4�s�3�Yg�=ںus\ˠ�)��V��	6�E�B(7DH���N�s��U(ᄬ�c ���ڳ-����s�Ic2x�J��"�>>�+	4橇���a��\���ڧ���P&m�#K�I �B�?��p_,,����en����a��H
]@ŭ\
@U��|br�P=������!��W���[1R��������S�F2��ey��P���YN6z��>�w�ж`c��YIh�.;jF	τ�?�{ɋZԶ�+���P��Ki��?T����5^Ȃ�ٵ��vv���A�kxl���h��]��wn��ᜐ�Pf�=s���\����~��W-[�,�{�B���?��[o�s��?=��[o?������y����`�c#=v�g
��ոHTM�0g�JU��Rr��K0��uμ9$8�x�M�6���}��^-�+���g]�M׫e���E�r�X���ce�Ŝ�f�߸ق�P�blĸ��(b�X�%C�1������h�1�M�-�=#���Ͻֈ�1�������ݙ3��JY&xQ�2dh=��X,14�:̽�2/p(���%WS���s+�ƻb�(�%���&�8�L*i�BL�2ڸ'�lt}�2[�bf��tbUgGǯ���|������iE��䷾u��o��?�C�(�!`����a*6���EB?)A��Pjm����)S��|�Iǟ��'o�}W�'>�W��.ٸq�b����-&�����r��c�� c���u`�҃O���?}�iC������~�=�������Jw'�1-&4384���"�̊�SXt|kKK-V���"�S{��FΕ�E�{[Zf���J�mں�����ef�����!IE���J�a%ES��z����S��W�YRR&�cT�E-j�gb`ZZ[�ѱa˾�oVV�'�C%����ajK���(Y�b:�w��|��W����6�AV�O\�Q|�����r�$� �EA�z�c:���D2G���	t,����S:m���L�5����,�R)���q^��z(�U#,;�+E���2ꯝ)�X�X�2j@1�]-je�c��Q;B�*}g�\xq�" Kܓ��P�J�)���	��ٌ ����/s����cMQ~�� ���X��2�H>���~T7��    IDAT���;p�ś�ϟ�{��N(�B�������^{�>����7=�fݡ�ju~�u� ��ܲ��^�F8��E_��:|����,U���uW�8��`�z`�h������݇#X�._X/nI0<ս&���6�'��6�jw��e�	���R�'cŘA���Ɇ�����1�X�q����]b@8+�?�|k��F4j�ش5:��4�jU��x��}-����-�f���Z_<2�~S�)ǋ��M\�@S�*P-�##��	׳J�3�qf�y�jq�����XW���0r�M ����VĆ��\�2Ɗ��-�{�����ξ��3N�����_��߽��GYuj�PX����b����XX�m޲(GFH�wYO��c��`�ZrWw�ڮ��O|�[�|������ξ(��yo[�f��6m�2��3��G@,k�祢'�=r����i�ϻ�ҋ?�|��+Wf�>�{J��~,�J�͝5�6]����ˣg֭5?%�rd�7�I�2vtU�^Ԉ�(q��y����*�%*�=��
�sgy�J�9&�� 7��x�Z�9��+�|#���	^���Cj�a����*)���:����Z��oRR���`[޷p�Q�j�,T-�
���H~��	J>{0�oP��Q฿��9D�Q����P���-:(^v��L?�[�V7 �V��k�"�%%� �l���0���R����
��sE	;�IG�x\C+Fּ[;N�K�j����w��{�+Yz��e݄�t�#C�'0�6L5b��_���l>$|<��t4�X+fѧ��+��;��Dq�_=����ƦMЈ��^��D"�֖ۢj��E��db�T(���^+����[^��~� �;Ｓ��˯��_��3564O����▵���<�˜3�;Qŀ`�x�`%���ZV�T�j*UVc�]�uF�Է~�Z[l<��&��c#`G�tx�׶�-c�����%�[[��ł(�kr�Q���`.<.Ak2���=ϥy�ZP�&
��U,$�d
�T,��6�����'W2,���ܔ" �~���������k�F*ώ�el��[�Of-a�M�� .�Cj��˳S`� \�.�l�1|'v
y&i�0r�>2R��r����s?�O�~�𥉉���K�����L������7��0�5*��L���G�k�f#��-�����������>���k`�*���yᯏzݺ�o۴is3�����l>����2N�	�tt����s����m|����pν�Ry?A�/����2�8�Љ����w���y����E��Z!Z{>�{3X��J9�1m�Ł��hll��pO^�w�)�X-�i�Q֎�)^�R�`]),u��k�](k�+����cB-N��'�:ߨ��P�\u��ФRD���e��<�ҥd���xcS*,"�W�9/�]��9�ܹ.��@Yl��9>����B��L��.�1�>;H�W���k�`��5���5��
dU���� ����{�lY�r9	:��f�2�@$E� �I� \�w�t���|g�q�{�����_sQ��ΰ��H�h� B��z2F�z����g\�F�!�,#��ռ	�l��j<�u�U�x��޿\.����ON�6���-��zj��Y�/Z�h�w	<
�}�[��ӟް��'�<zlllI*�J�6�r^�W�e�p]r��9!e�8ᚴ��Q\i2�`
�sP�Rb�;�.����:�9���> �cx8b#<�b.+ 7E}}�k��>�Kڀ�d��+]q]�̩�KƊ㑭�H�q�p�d	s>�g4�'N+�@�[��)@���ڗ�@Q3�3�6>^c�47k "p;��B�L�PYk
2�����Xj�3��h�� =m�� ��arqgn�J1���k�!��AN1&�D�h�i����:P! �]v#���)��3)d3镯}����o\t����?�{�Ϳ���[o?qKO�!�Ba�����6�g|y1����˵T������d ��[Hu�Z)Μ1�;'�~���-�_*�������ꪫ?�z��'��\�fm� .ȜdsC\$*� ��������ǿ��3�|Q��	�cO}�[348��B�P0���)���X(=��ݒ����P��*�TI�L���K��l��F�)]���U���oΔ�0�������Q��N��UըXq�l���n���F5��z$ȵ�B���,�*��'�3�����[����T2jK<3&���:�迩lp}+�}�zn�z�>�
�,�!�wL�yR�1B �e�r~m��ؒN%�=*\PK�A�*I��C���Wʷ�B�K�{e<��(vG1'܃bGs�po����<�@�-�:xյP�r�B��Rh<��`-�r�P�$�J*�����*���M:��g��V�J��҆iT��!X�m��<a��؍���у��8��1D�˰ߎWT`��}P'
����i�����uc;R��/��]�@���	?2X뢙e
HKIp�g[l&����}�Y|��^u���{��P ~��;�?��́�������:��)����YG,�F������A?55c�57z ��D)�3�Y�����2G�h��������u�cz���>Ykb�$Kh'm�2��P�^�J�׷���>��a<,8�W0���^��?c��h̎g������֑�o����p�L�d�e�1s���	���B\H��hm3P�U�}�]����`,p�9�s���?��(���$d81�S�:���X�z�������sz�2�w�,�Ƕ�:�[/���wu�Q�_��W����_����AJ�7������Θ���-��.c�&�x��Vg؝i��&&��jii����������89륀�������馛>322��鹘1$U� O�E�NV�Zi}��esݴ�6�uԫ���G>rϋ��'�ȝz�[�<�\�j���n7�=s�Mh����,H�ֆ5�ސE�`�V���:��M���ζ�Z���a��X�<aY-�#�Ԓ�Zx�o�5\L��LU��J�k�!��
�W��q���w�5�?]�x�3K �
Q�Ъ�Y�M,�,�h�G�΀�P=��]Fc�������1.�î�Pb�0�=����\J��a<�J~_S`�U �U
N�K)c0T�<~),�in��&C�Z���'�����5i���G�A섁�,� � �LV(�L&����P.�L�Ӄ�tj$�Ύdҩ�\6���Ը���ms�)?�I$�S�T!�L�3��T
��K�"݌]e����H��)����J�|�<�444�P,�w�JӋ�Bw�T�*WJ�b��R�t���r��V(Ӟ)���gg�{�[���0L�R�������\x���d�M��,�T���_J��0�cB
J{;p-����!+1�˭�m���Y���[6�[�~뭷۷c��a�*�t����k�57aJg�䎐�l�$X�� fڗ�T��ܼ 3"Di;�|\�a�w���� ���ˊ�f�*�\,��_��嘐��{�?�=X+0NʊP}�3����A�.T/g4�\�~7�o<GL@��IF'bP!9Ļb"}��� T\:A`U`K.��|yڤ˵P�r���F�[�2���K;gB�<8ݍ`���Q���%��rg�(/Y��o~�>��>mÍ7���o�������g���42v���2�sW�oةy�Ջ�h�����'=;����R�x����Ǿ�׿o��u�]7������}晵oo��y���`�0�ڶ�'�J��e��.��k�y� �ƒ�Zz�]#ÃKY��o+N�):c�t����>40��TQ�
�yl�B\�Y���X�,�&�ts>���b9�$Z
RcT(��L6oR��#櫥=����&V�4�,4(�R��Z�
A��g�l�8�@@Ȑj�^�YBG@@\�.T!�Q޻o��Ϣ��~�P��}��Pr��&���Cv+ �=U�EL��0-t6�������Gq�}LɝB�"�9V��I�2��BĢ�� (<�Ǝ������R>z��r�L&ݗ�dwd2�T&��ؐ����|z�)��:u�S�fM�5k�X{{��A4S�R�K=�k�I��D����SOmʏ�l�޶�o��������bql��BqJ�P�^/w
��b������,��0d\���`�R���kUw��m� ��Y�)]��l���v����b��hh�PK�����.����4�

�[�.�9������ȑ[��V�)�� ӳx)�9�s	aO� �� \pM����t+]L��u�5����ẖ)`i�d����bW���so��[��r>���
���4�\����8+�B���p>�O�^�8m8��7�̑R�Ș�"j���5y���1@} &����b"%�4�u���I�h���M-{n����Ii3.r۪�����X$�N�4���8b6X��o�RKK������xW2�j�R�>�˵Z}���f���-�W�X<�G�7 ~.�g�E���h���>���|��'ox������ˎ��;>��߿?�o��,��h�}��m��Uiv�mi~[Fg[�뮻|���z���ZOA|��s�	����g�9�J2���vjjZ�$S��@؄L�-�_�H��HTZ��۬P6�g#����G� *m�ii�6l�mڲ�@�-���	wL�N����m2O�������z��WA�x�<|�B�:&�ey� K���)F���>&*n͋~��X&��J�H��F��ps1��\��z@Q�-8&W����Bգ�t����Aຆ��a�H�A����6چ"�����d��E&���>�_.��8RC�t�7���hmm���Һ�����ٳg�6kּ���M���~��E��?ڡ�\sM�U�wl�������m��ch``�����RyZ�Z��Je�����es���&L�mEW,���6ݚ\�ք�-Iᄛ���c8�1U !Ǹ���F���i���>bdmKɅkN
G� Y���X�r�(>G�6�gn�l�����3�}�ow K �X3 M��m���4h=���3��}���dSkCu#d��(������TH�*�QǱ~4>a�\�n8�ix�W�A C��l|/&�7�T>�A���<)q��rV�73֌��>����6����|xƎ^f@<MWL����D_w�L��H�v��a�L���T@�X��W�V�r�1�\���c�j5O��\WH��}�|nP1�K���b�x��OPo����m#�l���,����7-[���F~����ӟ��|�I$� /V���=jeӵ'� ��50��G �rт�v���eG�{�i��/�%�L"�y�;/�����C�9S�z�5{FT'>�;�5s�u����iYg�ŚRlԃ��j�J��e�|&+e�L5���}F ORxQ2��vl�(�d�&�./��rMQ&��|`E��ѕ�F��]:��zi���^4����@�.��o�1�����ѩq�1![�yL6���L�p1i2�d)���~��m������G[3yӧϴ &̓>h�@�����B�RY��E�r]��ϟk��W�Aln���ea�~�C�t`��d�0E��,g��	ɳ�L銎<�H�~x�R)?����Lgw��,�y���,����ٳfΜ黺�/y}���e��jyr����Ϭ��v�}������6V�U�]R�T#n@���=�������ɀ�6���u%UOKd.1���bN=��c67��,e�5�XiN�E��b����`�������5�Pň(c`���K����`-uW,�'��-~ 댭���S=����� �7�s���֊�hs�9��:`�ɂ�Mu�ͷ���1?a܉��(��{���'1f@)�l!R�ώ���Ğ�|Js�貨�r�\����1��g���H^JAìk^s�� J��&7c9N�E���>�Q(w�Xx/X�L�\pO�G8�܇ߛ��j������SB�u�n���j�4����v�?�sG��_�����.�`�[n����>��_��g�9X�S�L�uK�ُ��\\��n����v[��o>�M�-[��ww?_�d\r�7�p��W~�*ו�Q>��N9�d�(?2��`-@�����H�<HHU--���0�g)\À�!�[��a崩&�o@�I���&7�r���(8&a.�=���/u[D�.s�=�~2Ӱ3�N&L�`B !H�
�1CNJ���r�pd�S��C0
(�.V�������e
�G�{eh�h1��#�5Ǆ"�����7��vП�B�*W�s�"�"XqJ���c(+� ��W�d�h�_S���Y$��m���=��E
8���`�̃�����N��R6G���������t��w���'���I����[n�%}�}�ι��[�<�����8/Ƨ&�ɶ����Y&޳AV�}�\�+59��_��G�t����p�mpu!3�hP@�,j�� F���H��������L΋o�&D�� ˽��#�&T���5a1�g���5�HK�[(��Q����7g�ʥ2#�A<�[��O����'A{,���Ş�v�q	�D����C��D�K�	�������o�k����aqC��3�2����O@U�R�0�e;k��Lx��I��W`z"��L�dx���#�Z6�c&+�v�T�?9�碧��d܆���f�<;K��>W���;�:��u?|�q˿x��>��Ȱ�����x��~��7��gHM�=�Ǻ�;� ����T� ���W����X���,_~�����l��y�}{}��tS6��5:4%S��oN;=�w�E�@ߎh`p{���ʬ�x�9�P�5�k=�T�:M4�Ы���Q�.�`B]ͱ(��}CQ�R�V?�TtۭwZ�,uR�MNM*-��RҤ�&��M�T�-b���d�1"�f������ �@P*�]���%<�nY�Z$j�~��\ks0�:����p��~���<�Þ���KOOO2��	���,y�Q���_��|��C+�v�p�YgE�w\t�o��P^���Z�7�}�Y�P?#e e�U� V_e�K����ن����rq�_���8�/]������?��S�����佲m=�&K�Z"B�朂Q��1g�xP��֔c������.�cC�T��&�����B*ǩ�d�\(=�^5�a���A��L�X�֘��ɫxz��N� k32Z�����Β�F����du�dM��vjMs,��a��}��C�B���� ��������7��=�Ʌx#6ſPK��(��j���2�$%C���r�LC!f�����<h5����1�����W����@� ��R}��� 1Ib�􊋍s]�n0]���u��u \�gkl�Mڶ456]��W��s�9g�K]�w�yg�7ܰ���o��m۶�n```���g�O�:Â�K��a� -֐{{��ǫ@$L�>c���s?�勾x�Km���j;�����سu�I�B1�F���Ï�]�
�@fk�Fc1�[<�+k�B'���&^�F����AQ���5�a�DƂS�nF�J4>V�֬]���ۣ�1�KQ6绩2�xM���8Km"f��v�S�u�Q\�(�Q� y�Q��I'���kD0p⺟@F��' ���֐"��@�+�{yE�ݢ���5���N����O��~xN6��`!ѿ�U���kOz�?.]z�����3o/�X.yJ�،��������\V֭����מUU�^�Y_��d �(�����#�oؚΤ�^0����={�9Ӝ9s^R �j�ܯs�}���~d��=[fn�ֻ�w��]|��###S�y����2��?K���wg�2�`	G�j<���e<�l#�ʜ�^��+vA˲��C��;����`�0Wp��{#��Y�n�װc�oYe���/�,��� H�f�u)`��P>�n� ���(mUMmC`�-����I    IDAT�<cOG��,e���P�(�I@@2����֍��'��B�C����
b,$�B�!F��_1=<'Ÿx'Ӏ�H����?zl����!;����������� X�9�0����:(س��k~A��ؑP��7i�z���@��B6��J�l-��ʙ:+�%�X���v��\@�k�ǳ�%{�Zݞ�gnZzء_�������e���f�����C��=~*�R��f�cM�-�&/X���]t������;�������K�oܗZu���8�>}�R6�@ƿ_�����~x�����|>��o�>ѫ������c;�667D�t*�[���r�A�+Q���-;�W%�H���T�R��Q�8>6^�F��t*3^���J�D[2J�fҙJ5�4�7WƋ�����j�6�-������r�`�%�Iɉy�Z���Ȃ֢� `r0���w����(l�ǽ>dX%Ә�eⱐ�`L<�����`da��ӀڂM�;FJ@lMh��[�,��А7a���]�淼�m###��{����Լ?�l~oim��]�z经;�5�������ի�qdd,X0%�=u�m���~��WG7�x�)�P������|����n7��gശ�E�Þ�TjcgG���|�:��G�,^�����k�N߶u��uk�Oٸa���m=��f���L-��]Q��EQs�X�%�\.אDp[j]l�n��SÜ����fA��S�y���e>�6ر��,�N��@A6�1�_��������1�Y��]���TI@���Ч�s�>�۲ys-��{*{�{�-�[�M�����­�I ����S?Q��u�7dX�B�"�?�b]
�͵|*�(7�b���Xl��}�u�DX<�e�y�)b'p����6�"C�ku�w�����
6exԋ�	����d%/��1
^ޞ6�\C���\!ra�]�w��z^�]�b:����S��'��<%�u�L@-������s���m�V���	όR �1�)�T1��r�Z[�~�AK�<��C�x)�-i����^�<��_lܸ������d���Դ��BL�v�����Q/�X�iq��B�'����w,[v��{�/\B��#�=٣�?�i��E�b�3�NwL�ڙ�b_�X,��RCKso>�JfңM��r6]HUR�J�\N�S�J&Nr�{g��t��.�J�T���-GKCC�����D�}/���oڴ��5��4Nj'�l�Kh�����(�b��� Ջ��"
z���bU5�$Ne��W����HQd
�b�`��2l�����5��S��ڂ�w=�b'm�5kVu�]����>��/s����Ư?�n�ۚ����:a�s�~��_<�j�?��/}���\:�]��ߟڼ����ם�����}�]t��6�=��/&�+^�8�/�}�Y�gώ���J�]/�%��/:���wo���;��EL�?�C��j��k�����L�G�m޺�U##��+��r�B�CJ� AjB�Y�e� R�a<���	3��ص�6�
�@�B�Z�Ж�ؘS|�pUF��e��jAxR>�����؎8�^A�
B��0#��]�:����f�奲�6��j�x��B���ߜO�����i�)\l�b�d�R�P�1��\�d�n�=�\�J\2��*j�'��\q*rpm���0/b�l�J��-t�%h�:\R����G�F.\�+Q�3j����ދ�W��YXj�W����g�rsɸR�M�Ċ)����b������	�b�Q ��֤��u�9�L�g�y܇�������vc鐋��-@6��
�If�!�ym_����:��TK�|>����n�5k��N8ᘕ/6�������y�mo9��o�ރ����Z��?c�4���fαv��ز����%���e���X�l6���(��6���O|�g��{o��3a:d�IH��ш���w{��'��j��&~r�L���$
���J�ңr}'W��k'ZhJ�
A�=���o��|&���	ʱ0"U՞*(��gYq;8D���;g� �@~���}�kO=�S���[n�e��>�K��!�t:;<<�_�<�����/�H]}�W�ؼy�T�:s��G��'��e�����u�]�,4!a��GM�:��SO>i���C�Z������r�g�,����fM{��-&�>'_J������OO}��{�_��U�7oZX.��D�Č��B��5s�#l:)RiwƽT�4cX%�RhΣ`�o�1P�^�m</8`a��|_���<<���&���x�Hs�6ln�A� �������~�e��\�2Ǫ	W`
�$ӌ�ɐ�������Rq����A�X@g��(�璛��^m�L?B���`:�u �z�.�����	'bp�^�C}��Ԧi��R`y.][�HrDl���|�L,	ó�։��6m�s��!7 �T��)��{��=#�ϕzK_�%�8�ɐ��s��i��u�n�#fKL��_�E�6��a�}�6�� *�J
����$�	p��r�i=i����6�Q2jo��)Y����t_gg׍���{��ﾻ�9}��m��6���s�w�v�W��l}���{���6�<��y�S�L�����]��	K�Pm<���ܚ�\���h�9\��.̝;�K�w�5��j��=��d\�����{W_��R�Ҏ��N���D�d�L鶼d�4�SD��u-M�P�K k��c�JS��h`&��s�d����oϙ	o����ߩ�X=��h�lzs"��T���|n��{�y��?���������;V�^����%��޽�5�y������7.;�G?��7V�\����%�d�+��׷=zlժh�]��>��/l۶�w��y7�[�P���F�~����z��iO<�ȾO>��1���+��̱���t��ؤ	,��$���=Kɭ3Yc��O�b���/$$ �ߜN����8D/s={� L�&��{3�������ܵ�K%��
���u����m�g�̦�D��Xp����!�%լJvb�-`� �g����uw�P&��C앀����T�x�9�"���eK����3��]����5+�����P��UQR�5�\�K Cc-�8tx[<ND�A��j�g(c�vlﯥ�Obt�]X�JrQ�H�ՍWŬiLu���� S�?2}.Opa��s��X�bPOCr9�`M�h2 AQ-��x���J*�� �V�G_	�i�(+�p)Y�;���������,�l�+��y�G�y.�Ɔ�Onx���G�u<�fu��O={����_,�����1P&�� ����n���`�z)�6>4#$v�>8[`����ۯ|呗�z�I��"�e�dP���~�/�J�P=��PB���b� ��|f�1h&<��Κ�4e.�aӽ���-y&vcN<P����lLF&�,1e�(]��B�.H�J0ˀ�8���|�yeG�E���v�V����)�ox*��ܻ|���Κ5m}GG���ŋ��Pn���r�Gn����X�rU���!�;�0k�#���^��W�x�߿~�v�.~E�\sM�-�ܲ��GV���o��j�:7�J5��V� �Z���y!���C�:e�EK���)�% �6ב7����!H�9˜d�]徐�&�LsT>v��o(>e@ 2HW���5�V+e�K� ѶPh��������l\xѾ�#p��w%�6S8�7��J�uY`�(�r��6�j����zp�S޴��g�Q��~��H�L�;��L�1�W�U_�
S2I���!���� ���
�4���m��%�hH���V�ʣS�Oʕvi�2�<%7��ԷRpV�EL��O��c�8��`����Wf��������vH�>	H(����Љ�A^�L�2�>.�}���X1�+��J5D�àU��@�����]@����s���yǢE�������+W�[�q���?��k�ث0R\0^�9>^��dr��u�9XA�D\;�h֬��yƌ���\`�L��T����dkj������@��9� �����y�{���/+�A����o���u>+Z���Z�;{����wFmln����J�pI��U.��ɨ`7<�5�1�	?���X��|�Y&1�)�Kv�v �
dA8�g!S	 b5D;�J'WϚ5���{��{����o�c�<���-?������7�}����Lj����q��Y�t�����/}勯�c���tͫ�����o�����<}pp�J����|�vSUlD���@��j�U(+�9��OR�[�:n=&Is�Kp� q�������V<O>u��Oh��+mYЀ��0m�n��3�����5<8���!0�ʜ<`ů=K��f|+{�o ,l[��#����Sw�{we�F/Y�\ۅo=>��M6J���k�+)3N��û��'�;ƙ��[�j�59�Z�\G��\�N�s.���D׋������<�[��<1)(8� �O��S���ೞ���c�?�m@V1�㽦���b4A���^����eq�N׶�"����{�Ma�n��y�A1\��Tu%m�1�|c�T!��, @#����k�\0�4~���
lU)�����--W��=�y������}�o�W���'ə�Jij��i��p,*%�6�/^޿��/ĊЯn�8X���<��9�;c%�T7���-h-�r�;��s��O9�?}1۴�!���d��s�W\188�|��#��8Bƀ�jJ����ZZ!�v�����/Ƃk˧
 �"�Ž��,@�0����|Q����ǟnjj��ŋ�w���޷t��-���]�X�jՌ���M?~��G��u���f�r��>�+�A���V�����n�m�c��O���k���7_q�M7��\.����k���:&��h�L\R8g��5_4�u?���IP����Y�r/��}��i�Ah�jŷΖ�-?:�k(K^N������(}Yݡ��h�R77Z���d��%�(UU�^s^�E֐���K�������@�*NB ���2Y�&���,��y�^π>�ڊ�7#����%��q�0�o��
�HQP$�K�U����oj������Pyk��-��c���.����묮��m��L�&�82�I$�%)�$Vkt�Y\Q�T��R|<��<&6#̘���8T0�'+�8�w�2#��k��.��'�+����̕��b�l-��Ҽc+
h��	� �^��K
+����������l+
l���(����������LG-M��'ʄR��I�|�s+[���_j=[>o��fWtvu��駿��˗/����'�_v ����?=��G=�P(,L����j��H�=[-&��"�q�)]����N��R)��Ҝohhj{��'jnn�U.�l��jSG�JY��L��z�+��I��W����zJ�rO�8ޞNg����ǆ���##��S�NM�R�͛773y�N�Z����6a�R��$i��[:�~����7]�q�ѯ���O��6�y�I0��իWϺ�'7���SO�w����
OQ�ӧO���:KsfϹ�k�|��/�^/��/��yw�}������ޒHDK��d�-;�e#@P���H�H ��)�!�T)�$R<�NYg��!:���q?��&�?#+_B�/K���>��-�%�f`�z�)hi�@���V^ E�G���.e�gV#��ˊK������#�Xs��r�3�,���(�����|l����c4�.����o z� ��0�H�ϑ�|h%�U��"�A��M� �o�w��F�$���P|��� ����D���V�(�� 	���b�A�\6��v�@�\II��2��А#>��Ɖ��\0\W�bqx&b#�,���yW���܁�a���K=���+^��������(�{��(�����cLQH2|<eWc(@(cV�N��P�\�ˬk�C�B)��Β{|����!����1�Z������Y���ؿ<�G'�|r����}Y��?T�]s�5O<�D+9�ccQ:�'�1]*�ք�d�Z�T�
I��t�Z���|�Zi-�˔�[�h�U�}�{W����y�m�,:�����k���~~�ҥ����֖�կ~��r��>����|�M�)K�FF�R�L*�H%��d�\����\��ᅋ��ᤓ���E���o~=��������ܰq�!�d�]������S�,�9s�l[��ޟ=�o�򕗒����/�v�����r����MMMӕ- �0F9��w�Jm{��&��N0�TuKE,���	��C�8+�pI�Ǩ�%�  �K��
3):��Jo�����h���ӴIU3yצ���fA�x�1ZS�b !�K�JD��N��GR@\m�f��6�B7e�~��"�-k]n%	l=/�Vl��0χ��1�eP��'�W�e`!��b3Ԗ�QИ<��g0�?큯:W��N���Ox)[	C��	Le�C���D~�e���؊��1�'����j�1`r��]7:<6)&��c4��	l�Z
J�H����>њ�+N	.�d�� I�<���Y��Ix�+��¼�i�G~�U��ܛ�7�y���V��\;�˕�6�cY��ݓ�OsH���>q\mpq��N�R+gϙ}�I'�p��4��s��/Y��N�5�����mmmI�{ｷx��'���!����%��p�W/�r͚5�n޼�����M�+��pju֬��{��Շy�%g����m���&)�+V�<覛~�����#��l���OT�����l¹��ݚ8���~S�c�N�z�g�$LD�"��2R����;b ��7;.�MJ ����E�,Bh��� yi�0��7�j�)/ALl�!��^e��5�=9O F0ڬ���s�3�W��=Dx�b��N�,�PًRW��0#���{���>���"�{�)I)C����x��K��P�����=��Je�T]V��%][.#Wz�V���ź��>����X^b<��ʮ�fw�Y��_ @�.ߩO���=��On�mŤ� !�������('�_�B�ɮ1��d�h�	F���b�S��[�b��] ��ȸ�����P�a�%�Z�b7��Ԝ�55O#�qu��1,���.�r���Z�����_�l���O�E�K6�d�Oh���=����o���{�M=��ѳϮ�����-�k����3��Ϗ^u��W|��-Y��e���=��3�;߹��իW�90�@Sc�m��`b�����
��L\�jk-#���Q����R@u6�}�\OԿ	�����d%�(�/+�c���,���:
(�0
]B��ǄD���!��~Af�A���3��*(�������().�+�r�Yzd�(&�����L,��K�-Q)#��!�B����hn�j�,�P�� �t���,�l�,��_ŽB�]L����LH���4�K�0�;{���[��|�(`- Z8Wc,��3�e��/��da�8�NI8{�?��d:�
��D&*ǁ�:��0Ł��Z������vR�S���!vO,����P	k��=�g�$�g�Gc���rM�� Kk�[�o�Vc�bw8�`�T��hNO��=�cc����3�̶���;w]��w^��ew���'��c�^���3�x�=����z�Y�_���l�һ?~�5�%���D��O�P@�Z,�T:������?���w�]/�.��.�˫���c�\�M�H���RE��Jt;�0�T��|�q����J���R\&x"r�Cy�*p��^��(�	�
�w�Q�`��N���و�Z�y*�#几�����JF�E�,'�E�4/Lvv8��D�3��`��\�Km�o���A�BpO�){�:�9����@��f���x��vP�
)�uޱ��� �򐵍[��؍R�v�)���&�Q}�qw(A����#*]��J�J5�{I��}�\�WVȚX")�)�P���Ř�\��B0�i�ޏ�i���ZrE��_}%�!dz�7[�O>��P_�=!���A��5���X	���������K�S`p=�6-r>:(~    IDAT��!8`����]�]���j *ᮏ���>`S5����t:�&��������}�C�^2�� ��0J�Cm�袋����G/d�oܸ���u�j��߈~tk�I;���LE}mm�����k�<��{���7���h�خ������=[�_�~�	���Md��"��O
�Dy�Y�&�1�����^6��[�̪.Ĥ<�!���V����O��h�|��G�n�*A�5�xa����k�J\OB)�P�f!Z���
d�!�p� * @�1態��G`��(C<�`�294b\��=�c�3�����ϻ�_t�2�,Wj���1WPV�����"���ewy*%u���%�!dq�xР�TMQ.|8�g��2(T�k�)�Ul�Ȩ�H��n��~�i!p�~�+*jwp�?/$�)�q��ҕ��� ddtCpU q��'E�F���y�J��.?�w�))]����X�������q�#M1g�c��D�����Y�7W��|4L�NԜ���;�=s���/��S�k���x����20*�Ħ����:::n�u����W��O��|2�� ��z���<�������n��v(�zy��u��(��e�#��#d9�၅����y�C���������e˖=�|���T���������𹮮����B�W.H%�
�g�ٶmB�Y�cq��5���l�iӬ
'BS��1����r��;�	)�*�����Q	WY�
���V�>m�,�D�8n������\���l�1������bY�Y�JUA:����U�|cM�c~������E"&G�

���#C�\�R��ഗ�(i�3
u��`�Y����{�s\C�,:(�����f}e�����#t���_����������UH�y`�c�)V��Ǜ$-�7�%�z�+���hs�ጚ�'
���1	1P��+Y�Y����K��٠���"Y�b2¹���b|�wM�z�YMڊ���h����A�#!|���k�MtҤ���g�4�t���z�i2��T*�����:�o?p��?Y�t��e˖�����ێ?���c�ˎ��o,���{�*�-,4� bbc��,YD��h֣�>�qFF\����D"����{���<��E��]�h�e���5lw�y�n_��W���O�����Ͷr+��`�
���jݺ��z�c��EaKAʢCL��U���bG�(�w��<�K�#{�G�2�5Op���B���F�ڕE'z||l��A���u/Y].���K �
�"ӵ9BIB9��x�+mV	��ŵB�\l�g;N��"�2�or�T㮉\��ܪB6O��˼�ZR^�{�-E�|ߓ�ˁGR1��ꪫ�*�ִ��.F3F�q�	�Yp���	�EE��3/�ɩ��V��i�P��s�;3o��믫{��Wu��ǰI�\�b�y3ϴ�^yR[�bS��lH�+��H�g�ﷴF��^�}Y��qq؞�s"�Q�1�N �*vE�$�3��NV��-���]�2��'\q����1ʅ�0}jw�v���\�sL��(�e�Q0{Z	��"��G�ɑq��d-f�ۑ��1� AQ!]cHܞQ��������!�������JU����2�g���TY^�I�m���W��>�aSq5��T��ot����a�.[����R#����/"	v�`���\�>�jJg���A�2�HĲ��������þ}w��6=�{��z�o���^�m�cO=�v���y`�	��WF�}��k�W	s��w�t�b��Fu�؎?�\!�� 5� c1��O���'o��)`���?�i��J��s�0����FtO�,��4@U��V7hu.���������]���v_�\{�qX�t�v���ُ�%�ǹhɞ��ag�����%�/�H�����b�`0��զK��̑c8UJq=`��j�� :��� ����ϔ����~���s�t �.��y��:�I[�� d�>Fa�.6���؁ª�zU�	� t�LIj��z=5�;��[	y,r*��D펟;�y�(�=�D� ,P���8���y$wG%��!X�1���Q����� ���{�=��6{<�P(\��Wd��Y=zl��>��~����7P�����9�Mi؉'v~�_o�:w].�?$�f@C�΃?�\�s��/?Wa���T��0��2.�����xEEE��:��ԩ��Ν���ҥ��k׮�`0�VRR�ԩ��D���:G�u��}�&�������t���H��j2�Fe�Ca/�3�P#�+L�#�ҧBC����&�v�b�-�� j�G�p:~��l'S�I�J��\�D�z��ag��(�L�N�%�PS�A�1 �]Z!'��	z�h)�J��&�R�W��5U��U��r˨�����2�B�\J�D���+U��%<���Ϡi�sƽI[�Z���%�fʡx]RZ$���h�.R;����� ���TQ�;A��D���5��p�h(��=��)���4L�8p�o����KD#�J�|�W��$=�5G� ��B��=�@�< ��dM�\�q��{���E�E�eœ�%e��L���������c���$��T��f��l.�3sa���A ?_6�����p�d�\n# ���0\���x�\6(DPw,`��^�c@��l�@���b�������aTĒ�_-��q�i{�f���p�Ì�\�v�����V���:�p-��}3:Wu���V[��M�x�N�\/H?�'r�mꀌ�f�M{��+W=��S�L�f�e�t:�/=s�\�h����`�0�?����:Aͷ�q�" 㐅�>�w*��e3���z<�6�����mE�E�E�%�%�+��KꊊB>_�)���K*+3.�;�v�s��Ş%Km1}����ZZ���zK� ȓ�J+ԑƵ�?ܘ'��|����\"Y]� _/������@)Z��d T�i!\�hI����:}�ǪMM$�p���B�'�@�N޾zsY�$��qL��	j k�#��*�*(�R�@��j�t�\������VP�$x�5�6��
�\1�������0B�� ��`5�*LK0��m�W��-`_���y��rK�P�S�\M��~�u$%�
�D<i���Iʈ)3���/R	6��E"UMii�s�8�K����`�LNW܅���?�����KtF�n���ˊ4�s��"��3�����^���x睷_Խ{��_��QБ#��VT�����nw���������N�R�L&㫭m	�r�h4N$"�D"]����d�$��UfR�Rӕ)N�M�˕����t�|��ș�`�f39������!���v�\�va�
���CQЂ�BhA�vgq٠������i�\IK=:�u����*#�v��������^wSiQ1~k�*�[���**��u�V��҆�{��=�2���Ȏ?��k��5{օ�T�#�N�V5PY�I��$�М���T"��B��U�qcU�g���g`�R�XErf�Z��L2�L{<�,d�s�\1�����É��6p&R
z�W�Z,�# �sO�4?Ng ++��_V�ՕUV����#��ґF�+��^�X�*� ���hM$4�D���0lMg��a�}���D+T��\�)I���zW�X&a~�H,��V�|3�M�+��"�S݊L2����:�A΀�V���My���!U0q���~zo�,4�m�l�
���|�����q>J�S0���y#-"m�^������mq轠������(�F �xy���ڂ)��Q��^�%/Þ
��m���qa'��țO��+ �L#�{f�(tuƗ��v��z}�<^��-:w}{�=w�r�UWm�:?�	��O>��V 	7׆�qW�����݉D��v�}��+hIO&�a�͸ݦ;�1ݡp����\2
�r���0��2�:t�e25ي�xfs�@�-�䀌�e��h���{��/'L�9���Ji�O4�A-mdYK��аz�L�e�t@$������ԏ`X��=�?��2�`}�{L��E��![�
���0�y���:X���8�-�z�C@�p��yΊ����ȏ��hl Kh�D��2�x������Gm�
�X�8ނp��C�6�j��2"kKS���ƌ6�f��4�RЦ���V���Oer�N�6s�ۂ 1�ӷi�	\(�U�������b^+�GQ�FH�-�RH3�N���W'H�ypH��V[m!�ù@��>�����`��tJ�R ќ�X�i� ��F$�&!H��Y�xY^L@�Q>V�ฐ���`'��1�/�_97�҈�~'A�4rf��2Vx|���᯻u���N��4ذa�q��l9���,����d�����;n�_xvX{[�l.�)��
�n���c`�LA��j�������N\�/lXTj����
�B+d�{���l�9W}xM��N�ز���̩�	�(@�-�hą�7ҧ �Q��[�.�Z�6"�q��W�((u�$�JD \pR�#	EP�7G��b�``[��X^%��J��"- ����-[b��4���@����0:Z��a+�[lX`�<�#�寸f�LR�2!ω��%��^|����G+$J����ƪ��Ag���bd�y����#!ꔕpg��\p�O=	�+Z%�KEE� ���N���(ȴ����.)�����I�.9SZ�+��%���uW�IH�G-EZB���:�}�q`�� Xʨ���9��41�#@%�����e��I"32iH����B�E$ʣ'�T�=��7�Ls���^����nѥ�;��ܛo�������9dl��m������咽�|ٲL��+�Bt�\8'63R���Ñ�	�81�X=�Y���u���� 0���AKG'�V�EXU�Iӵ����<�������G����^B햰U�\��9��#F��X�&Ǌ��t@�<��`���k��ح�_؀?d��Z)g
Bb�-�U�F�(l���Hy`E��!ڠNUAq!BZu'2��R� ��#�����hX2��b� CW����7��1�V��%����X�1�ư?�y#m�t# x���}t"��Iu�J#*6��C�ϫ.��H��T�	��)��ĳ��[�#�^PM�CWR�Nh��`�q�b**=4�Bm�|�ŭa�$,� yB�5T&\�_0^,�0.�o)�fe|�p8���{�u��Yee���f��_��խ�{��ѣ�:j����`~؜��58 c��r�h̘����N[�d�L��K2�=�Ar�2��6?��Ѥ���-���X���J�L����:i9;��xO���g��j��S|����X����z���\ � ���͒gt�	E�J\伷꺅TM dH����#E��y��c	'y*�E��:$-�N	�@�@D�|>��#Ays
�X����3�T�5�r�1�q�h�pxΙ���p�LIX�\(K��A���J%�
v����	��+���Z]�(9,$�2m�H���Y�~j4cV i�b�<	Fmt��t���#'z,hx��þ8&8;�~`D00VYYY��r���n��|䑇N�������9������-������v�����]�pрl&�c2�,g)���:Bj�$�~|ƒG�L��+#tܚ^A	�F�n!�٭ �^:4���7�Rط����@��[rO́� � �K��ܲ��ݡ� '�h��r� i�C�d�}@_�^������8;*]bL�$���������h�N�ﶶ�6p���`��U�B�<B&T�XU�J�8!�Z�!I�Jc6[���J��9����P�c0"E�R�N��z��
(�n�85)%t��Cz��2�G�*�	׋�����k�ؼ�I	�T9e$�~��� ?)�P����?� I�����a�DB�' ��p8�r��[^Z��Q�\;z���-���G�9ݍ��ب.��3���TL�2a��L9���yߖ�D7�\��r�nii���\����24 2 ���;�`�N���1{*���#܇@���*���ʅ l'"�6�l#s�&�F:�1�x^�Q�}�C�++C����d��N	1p޼y*V�R>����X���0|X۲Á!���;���/5!��¶*��+M��\��p�J�q)iΔ�D5��K�%6+Mp|�U�t	��
���c�q!��b~v%�t��XHT!��I%Mo(i����� ����f�*p*��s�C�M���$²?Ik����v����8,��P�ʟ��M��|Y^Q��!�3��+�n<��L7w8 cs������'[~���͜9�H$�]6��:��i*B��C�.����F���`�$<J#�
2
i��;E8}(o�._T|��6��S$�����X"�US#�}y�r�pY��(�9:�V�H�`,8<�p,Z��jO��@�%�ad�I	<���;_r�Wa*�o�<� ��́\�|?	��@��-G̴�b$�Dy �d��i�V��:��`%�v�+y]��aHKZ�����J+��AR(A�d(#��ԑ��tYk�-S.G;�"T ��~����S*u�/QA�Tk����~���n���K����9�c��jd�Us:���L�����{��N��}ΜY'466��$z%��D*H2ď1���=�R<���K	:29�����_�{��c�
�EaZ�+g����s�88l+Q�2�g:� �=�&i�귺xb<8��b�	����	��kn��[p�(�a٭���R$E���FF>�`��A(/�-+{��<�B8'T� -�T�����*�@�l���A��s�C���~���h���l'�b7*NP*�`K�C��O�)|�����F�=Am���>�S2L�ډ�7^̇m�4D��q�pP[y��	�-T`p�P(8}��}.+.�{����q�628 c#�`��t�/_~��}�o̜=k7�۽e(��ek��OW�*����!X�"N��e����ډ+q�B�I����P�#6��p?V����?:q,uVi	���5/]P��$��hkѕu<�-��%M %J+=����'���p�t��\�~8��ᡄ\%˒#���t��?V��Ƹx�^�/���Has6샨�inn�W�Ў�r0������=�u!QV�K�?SN�%t\0����8>;Sd6�]0rsi��)�UT����\G3�<ޗ���G!e�H^���#;�����`S��;��Y���5� ��4M��X1oޤ�3fo�t�҃��N%S]À�h�ae,�#(���C�v�z�����h\�H�x���>�,����h87lk����k�� �����Y�,:pp�.�3�N�V,$�)K��_��]n�8G���t���ܨz����!��(H� ��Ab�@�N[���y���xɳ%/`A	u%D*�a�#C��lsn�� ��N�Gm%z
MӨ��k �S��4z��^3�1�A#jx&0 9��v�0+g�"O�C(ΓcC᠑ˀ7�hQ���$}��t:��m��t�^{�նA~a�I9XC8 c�l�~,��g��,\��l��ť+V�w��]ѻ��a�h{[�D"U�m�4LO�i�E�X����np�J��*�B�T#JB�'	^3�/�H�3�ʔ��/O�K>��������	�J�rW�T�\S*Y�h gJ'��t�T'�=Tg d�A�%���;	�8U�T",�5����%�P�����@�$�.�l	ިH�T��j�D , xpn�mH7Apet�:P$ �g�s��+AH:�)����Yi��i(���da��2`�����v�A�7��!nC��Ϩ��F�("q������ �	���nݺ�����Q27    IDATL���vg=��#�Ϸ�9�c��gd�=[:#�c̜9�d��Eյ�WTΞ��s]݊]&M�|f[[�V�ب?�\��@�� �
?���S������N�az8
{?F2x|��I-DW�F4�&N�z�W>��.���m��%�9BO,n5�bڂ�{��p$,r��zt�.��Kp'��LjTPQS�3�&@�=�C�(^ϝ;7/���)���i2i�Z&jWeZ��Jl�ϰ��!�:��#Q!���/\�������I��J\Kr3�F!(`��>"���Έa�h|[2M���wd���PWoTUW(I�-))6rfv���g9p��e��+�α�Z��2ֺI�ק.�誋>���rE�B�UD�2Sѧ��ހ�cƊ��T8Tu�=�������p�"n%}GT��\;I�ɹ�d4��Ϊ�p(i��<N%����Ph�ș��@��(�%3M����RMF M '����A�q؈�yv��-s1R"�&�ϧl(;1:dx4�Λ�S!LM0����u��ؙ���oo�J���nH��QW�2���5��h�>-m�j��Y��IL���{1b��p� h8gF9p� z���}p ~ .�Њ��E��<"Z=z���ε��۝���<�>�Gα�-8 cmY�g�Z����2kּ����G�,X0�0���� ��@��j��>��
 � ��b8&���<H�#F�
��Y�b���:${����	�rHc+8�}$�5"��pt�������Ao�+!p��+�M�yju�*zbŌ�<,��`�ȅ�lX=g�B�q�Z ��4$�2� �{`�z1�|�.�W�4�衪£�,�d*��ؼ��K>
{�P1��Ɣ;Ғ��% �jJ	8y�ca�x�G���O�Y`,���P�#���l `������^�E�4<0�J$�-��BlU^QjF"����!�~x�z�B9w,��,����dHg�uk�4=��2v�o����W_}hsc�����[4k����dgB2 K�� ���������a��p�U)��p\��  U�z���J�#�<���j(M�����	*���,^4��Pc���D4�v�c�#�Y��!��m ���E��$�M�>�`SH�����h�-�a���W���~�H�,
���N���"=��HBe��$\���+G��ɳ���5��jj�eNHQ`*��j*E#&��y�v #�4��<y,J��T�1h+V�`|��p| ��,ZYU.s��B�U�����~��c��w�z��T2�UuuE���m�j���4��ч�oݺ�69Gs,��Y���m�����[}&N�f���g�q��%{��E�y=����5v�e��o�ͯ�:�m
�_B�p 
pp�Ŗ�%�6S#  pV� ��r��+!SW܌^��8���e�
I�   ~��IE ����ŵ`u��_T��>V��L0��Xi pI�-�+����$��ŒE�%�Fc3��_A��{P����U��QB'���+V,�s*� �)!����\�`5	�% ���4b�@�U$*I�)_��qN8�F��{/Q�!6S�֩��Р�M�EF <�&�30�猔ᾁ��/S$�d<]���T�Պ���ٮ�ŏ?��~5�z뭊��:oqqq|������+��X`�Z�����������O;;q���;j�E���mg$\���@�O�>"���5>�#@� ��Q����RMt��#a�$�'@2�	��g(��SL�أʯ(H���@'��!B��tJ:ע���X�"��N�L:H��׶���8i���-�SX���`�58a�K	����9Q�~����2R`W�$���D�T��H��d�q��F/p��l��HDcy�C`A`�r_�����0JU^^)�����e��c�Z��e��p�\�B�K+DymXu�m1_�ၹ�02E]���ƈ� �)0t�]�_�~�ݯ��޻>��{��ܱ��ddlJWs9��'�z͘1{�ys�Y��Ч���G4�,PUp�pp(��e���;"�5�� X��.����ꎐ�F��*�߳���Np���J?�`�� �%��$����4]WTm����.����֡A�;%����.iPJ:���߽����s�Z�}����d��y+�����BL��M�Ok$��j�vz(<�$��H���_���
��hv�_ǅ> Ѿbhg�Kܑ��f��9c��oeXi�2wè��߁��U�I*v	ث�IHJ�>���<MM�$qB!��v�9��	��^�����Z���A ���V~"Ll��a?ӯG_��u��`�4�w���،�����YRw(�x�8L4��G�����r?�>F�m�Ǳ�e_>�Ԧ��NAv��j�����Ji�?fg�~�M���y&Q~)�T�I.B0�D�l�"20�2a| �g��B�D��%�H}���h3f��.�G�ط$�h�F�?���o֥ vZ6/t��l,'c]F�փX<HTCvJ|ku�t �#@N��E7
�CBS��An��KG_Äl8V�^�E�" ����a��ҵ�^�t1
r��oog����-��b۝v��$����ԓa�){������;l���9q����'��1�݊�f�: J@��eiV=�P�r�-^O�������o6_E�t�?��B�$��V.ձ�to2�D)uL�:1��f�߭+�3��������ieo���sM�x��{��!��5�g�����<*�sGE�G��1�/,+l���}��-z���"P슊[Qr�,>F\,��^Gk)G�F��?	
{�gM� ����F��=�$�.�R��pp<��xC������pƏ<�4%�?��1�ɂq�λaC �!�0���إ@sB{ՇjE��a����iu�滒���N�?����Z���혬\��x�h�Ē����pbdd.5�-}{��ȅ���yn�f}�|2��������
�8 h'aQ�=ZZ� �eJKX+Nwx���(W�!��l2a�L�:�}�,s���\|�Ҧ(��퐷��jc�5�{eF�<ݟl������e1y�WI���}nrm���m��l��,z =J.��Q�7#��H-�X%�n��,�d��Vrp+c0r�veq+R�Sg��i�����IKڵ���l�A���.��H�bpb~��n)���A�F������늹9/��GC���
��$�<��,�����,T���6~m,i2��Ȝ������N7-2:�L����O�����_��Zk~+K���uD�R������ء�I�0OL�
���ξ��$��|d����`#Èp6Y�t�Kׅ�A��H?«�������*C�h7�'�u6�w��V�z�B���	��4�O���`F��-������Q
��ۻ=�}s؆�C�ODmP)�K��55N3?~�(�h؅���	����l���K�c��D�i`�Շ*Ƽ�[��ڒ�"l�R�zt�ްD��!��)�0p�o	ɚ]#���H�Й��^��h^��*{�ª�&"��&!b��ᇧ����Z4��q�(~�z�}���
pAU�05��5+�h�<&�f������e��J�֟��p� �(���Q�M��� �����[�[ヘb���0�W����-r	D���Ƶu�:^�'0p���?�*+C�,alw�9����f�Gp]>_�n�a���NA}���P�p�����0�!r�����l���6��H�3$����M���*�7
�'u���H����������UQQ�\�f��#��N+n8�7���,�>�A���G�
*:ݸ4,�u_2���3��)�������e�Y�[B�&ϬRۧ�U��lH��[��d��8���b��o7cM�zkYE�3=obd��韞&�׻
{q1�O"���C�\�@J8�`
�tp*�tb���dm�_$M��@����0ovDQy{g����?�>u_����_�L����-?�.�TJJ��~�2�$�.�Z��˂'3P^�`N�����%wSKx�>x��F?I��x�Y�,����U����܃E��D	��e"Λ���}�3���b}�]�sO�ES ѕ���/#�^Y,��z�y"�~�hC�46����䗼����}5r}x!�ֻ�B�:c+����8C*���t��n��/^�5�:wK}�ꁶ�d�����6m��-P�F�J
ЎE}�i�[r�Ɨ���NƑ���]G�B��=��bM�m̄w����pmM��1���8�
��;S�C9�8�~�hg1�½����,�G���?*ƍ�۩�:���tvz=�m���y�u���s����V�A=�}Kb�Y.�N����P���t�����g��ˇ}
��s�qD��;N55{�;���fl	>Q.�p
 �B��	u���$$J���v,,U^��Mj��`�x���,pp]�/˙Y��� 4���^���q��3B �1Fx'Gǉ6,D�+2 ;��"j��&��م`,1%*��^�͕���te;DYe,q������	�Z��b0���ղ�D�/��T�g�&�A h!�Ѻ,�o6�j2.��'�	`c�s6Z$B��q`�5G&ӷ��ZQ��)�����&�5���0�,|Pp�s����%Ҵ����\����n Fߟ�MϾ���F��������ꌱ�@v0Zl� n��/�� cF��)�nI�µ��f�>b�>	���F���=�WT�I�٤ �����58A�o��ܬ�+��T�?9E�n�8��Tݷ��=l_cv�W�z���O{������}#�C��/�?�z��(eh�4Az�s��ٔ�H p8�r�\<H
"q�}bt�"�ѥEq�#�>7�!!��Xr�U�r�r�c�k~�
����-���hR�� ��`�ña�BƧ�͐�3p��E�mº��[�����Z?F�2SR�8����K�)��9���X�� ��P7�@�|�}���R��9;���q,=v�-靓�~�e���jE��X��}�V��]�δ%:P��ض��x��<��.]N9k�u�@�Y��ٹ�H�{�t����T=�[�w_ϴ��w���~sb�-y?O���^S������;l�h*�/�Q���a_����_J�D�ѷ��� ��rH ��V�|������4$�����A�\]N�	���Cr�0��֌��I.��p�Y3� �kO�5�D?���Q��Ir�2����DR��(�W��g��I9T��	����6&O�0��\*tX>���G��S��F�[�H����&Y�W�d��HX_	�Ƶ
�8�߱��(Qk�L�J^�\��@���x�9�!z�Gٕ� �_�f5�����H��lgd���V�I{�Z0g|xg%1_}"��d�k������0�*�Y/��Ql�VS�'� �CZ��{G����H����K��<�_��r��.�>��O�7@V��i�9���@��x����y����A����Ʃ��Hg��1���6o�AU c�}A@��{�o
6Zl������5]���ka�����0s"&EͮX���OV0|�{��D�F���$���~.��F e�g(X˷W�خ�v$B�q/fUbAָ@Ke4�)��Z���]kKs��b:VS8��;��R3 !���&����{��%B�k y���}��{�i^*ϭ�ϻ�G���Aa��ҷڷ�`�.�s��L��޹���(�B `��������c�M�w?{�I�b��?Q��'L��F688(��%h�r�W:�D��m(�i�7=�3�o��	�6�����y>�
�Y/v���ո��$�uA�~7[� >z�I���+s��]�H
��L����$�55��hC��B�e\D"�̺�f��~q�/w\��}��tP��R]�����Q�z�(V��7m��*Y�zQ�1��B��Sڸ\�^ק8TZ3-1��:�S�,���+�R�-�:����?Z+�M��0A��_�!�]Ƚ�=x�m�����}�G'|T�u�y�}���#4$A��[�/��|�)��JfCmz24�4V+g��m��Cb��mz%����5�맦K�ڎ�a[�N=�$�a��uS�Ex���D}�� �Ū�O5��Cj�d�:��۽�rE��Hn�#ݯ��1���i����W���oE	#�wW�������AnQ�x�X�����l�@�1��]D D�����rh���E@�_謽��W3�$^�S��u���"�����6�) �>���3�+�L&˼���=��@�V�L�@�`�&6+ �����k�r	� �K��F��������ŖsG�b"���3X�åU�+M�F�k�|=}�8�^��9�/��<8�)DV�ǤL^���r��;y&��J�
A���q�V�LA9N�q�:�~g��s��?~��r��WWs{�.�u�ɿ�!Y�R�eN���W�o����"�R��aHwgPo��n��;�ZUU�5ɢx��t���n<_0���b��P���Y�5W�O^,I�'�qb�w���%@�"*��cda����q+���=�o<S�K��$Q�0s�G㲴�3�ODZ��\���\�#� ޱ�b���7�a؈Xb�V��pZƎ�;��x�2癐���\?�����&�H br٢�`*3|���ȴR��ؕ���ٕ&���Zi����{�<>E��6ӥAP��윣n�����]
F���������i��XAz�����GM�]�5�x�������h�Z)��Ib� �o�2"���7I�ѱh �����#�K����+u�i�?��U��ɽ	N�b#0�7��j��|Y�HF��
�7�4���c"ʀ;��1u�hS�Z��{t
ߑ�ח'���k0+T��!��Mj�_m��	�@17w.9� �ܜoc��e�@VD�,ez�}�x||�&�U����-O׶�R�l92jt��M���C�(�B��t�q9����F���,��'��T��A���T|�p�8m��(@((������DX�f{��@���y�ϋ����hɇ��
LA8�x���̑�E���\>mK�#�-�J���$�e<��
m#�ܫ�]Ɖ�#GV<N�/o�T��R��-!���S����<�fꪵ��uL�n�)����C��|��@  8c$cW�����;�%1�B�/��|��??uվ�w��3���iU谗4V\���5�j�h�ՉH��,V؟���qrp��JQ���]��9����Z���,���S{����T�^[**.��Y[��SQB��S��ӕ�]:���l�ce>��wtX+x�=��z����xT���PL{�X���^��m����E��4�a�6��0��>p�Hۦj���!3\�**<f���V��}�	u�X��*�/L	-��pKѦ���������  a��d��P��ߒ�?��Ճ�C��9����i�h��������Yuߕ��N�u�ߏ�#c2�����a;Ʀn��m�:"���8e����l/�=��\C�"	�D%(ZJ6�=�;5_pڑ�����P�Z�&�(-EB��T����鹮�-z��ބ7�;j���X����P���۲j46G7�����EI�S%�;ܡ1q|t+���Vm*,�����cz��&�����qG� �����]Qc)D:]�+���Z���쭗�Q����8;�L̉������Z�t�#�<%�0��L&5�F�����8��N��+�s���Z���US`���@V<dm�e n�'�tj7�p���C2�,��AL�Zccq(���0W`�% ��H�k�A�'�c���w,���ay�	d����Te!���
�
���>�$�]�q��y���)�R;�r���{3��k/:uԫg�f�(���޺��=�W)�#�`�0G��~���6���S���u��PG�1��������1������s�̀ �KAIuպ�AE�.��B�/!X	�F�۫��r��UN�_^�d�t���;�Zo�������"���� ���z�.����%=J�צ˟l��-�>�k��)d��V���*?�<u䯁���:x2��"���2?������%9����迪���)�F��� 7)/2��S�����x���{�椀��N�lB{H���:䲼8�[!Q����?RB���QVWkbo�	zb������Wg]约;l��{t	�M��%���G��لt�\����U�c��&����>��Ѷj�~��zE,G7e1S�0������
���;�nܴ�ʔI�1�Ê8i�40BT�\���-W�53?�����S�=�+͈��;8�_���k?�s�AOOEΔ�9">� ����U8Utq��: �� �0��Z��2aT�ѠAS�`�@�Z+h�Ƨ
QL]�PM�.�V���YR	�6-X�`N<�d	���bґ^����!*�Z�D4��?8�e���%l�J�Ά������*�����ٍd���u��ܞx���/�:ꉉ�n�B_EA) ��Բakaɾ���t��5�]���  e�N�Z�k�(��ͫO�JVZ���S�T��9o���qL�֯&Ȑ�f�*e[Z��)(�">�s��T�p�ﲸ�ʹ�0��e�㉯���+����'�f��6���@3?��ѧ�>ם��^l՞���B���AwkU}����;6��N��G��,q@�(ݼy�H�#ȉ�@IveoqD�A�[�`-wBT��MA�XFȥ�B�G�ЁۗdGذq������0l'=*^��C�=օ���u]�n�5A͑{4���\�\����[8ׂzIv��]yI��]W^wx��������_���$�\>���k�/O��U����������>�p�@�@�z�4�n�zs�邂E���Xb���ǎ��^ݕ�$��ߣ�G_�lr��������xx�x������vj}@�O�8�}B3�Ǆ�I�ӆ�����Q,4��H
s��T�lj�% y$\���tD��v�:^,$0	�O��Mo�
�v����Z�Kr3T*Dgs��LT$!�\@�X?��s3�r��ίy������:s!��j%=.��W`��X.�/t��9#�3��ד�7��~����Y�ܸ�W7[�ab�ؖ�c�����N�8̘�F���qU�ɍa�է,JjUx�o�,�v�c���������φ���w�^�(s*nI�~m�[=�L�T��(1��	����^\�.S�y-CM#�T��Á�t����B{L��f������ �����Q����QNP̅�����	z�Й���v���t'u
�`6�ӘEQ�`���f(�ˆ�d}�����I֨Xd�5G�Zۜqc4䈠k�Н�CM�D����0@�D��a
*��&PܡTu�{)���۔������`����cf���7�0�/����|��x>��q}?9��)��I�瓔N�]�X'LK���QU\r�6�`v0���.x.;������D�?�l�y�<m�P��N��(r�6`Qs�̸:�F Q���8�'-[�4��]��_�p��0�x{���S�R^o� |�WޘeLg@��(�A��CkYYFm��p,Z��㱠�d��.Z͠a�Q�OV�Lٴ��x���Y��ލ�+�'�������3$j�C���/~���xĎR�Q�4�Χ�U��a4s03����+�����EO8�z2M�����"����
	���}"��nç��Bo��=s�q�\�H���R�X�`[}<�u�C<7�8��(:�8��໱���y�Og9�{;�t��}�8�<;x��ϳ�!�x����8Hs�(|K�1�1Ē	E9�EB���i�\����uڊ��s��. �9� ���������7\(U��z�n�z����f�ev��?3�T�I�0Q���O�96�S�N�E�©�\�w}򨇤 �x������<�(;�+���ŏ�"�x���'�ę�ۇU���S]%�(*F_1�áIi����ʿ�z[�; �9k����_fz�C�7�B��\��pa+�����4�Ku�J	<������wm�S��GQ5~TV����~O� �g�w�ש,ܐ�ݘ����Y�r ��d���������[�)��O�	�扚�戫@��x+�&����Yj�!
I��]�+��*�Dk�>7y�upX3���@Ts��C�E�:8��@}������0�~r����!����RC�`�8����YB���N�i��쓓��mahlK��+m=�=���Q�X @$܁��:�W��LS��5�{'�b��FTU�qq���, ܚ{e3�� �[޵����i,ݴOѳ�"�)���(��)boNɊ+}�����^�{�'��F���G���"�"4I��@W
^�^�0���v041�'E��z����4�R,^��}L t����J,�z�}ί���E!��d�G�_YhHC?F�_�7�����}����*�׀0:7��]��&�m�Zp�& �`#�
�4I��̕)y�L�����p�T���M�_�yP\�c�����/z����E����~�Ӎr���i�dW⟳:۹Cͷ�d��Z�u���}�m4�����4�&׻�w��ޞ��]���c�sj(�8TTh*J����"uIg{f9�hl�AP9��R�go��jb�j��-*x�zN½{�������Cp'��׷i�7�(�NE@͞�����jK:��l�졖.��~�`9�i�	�f�B"x���ZY����&t[��*T�w�:�p��A|M�z��Ӻ�W�m�_T���;P� ��D�c���x��_���xW����sy4��q
�?t�1��H�qՅ����j���W��NX��Pd����V� K�&�p| "9����5�{m�����9N���񞶵����N����zv`Z���E�"���+p��5<���P��χ�U0z6褲ҞIA���E@vBt^�ZLP
�L�!�mR��X[]{wҽ3M���y��X�p۽=1y#c�$G�D㘀��";����Bۏ��G/Л^%��?����M_K���eJ�Ё2�}~f���_��r}�v*3��l|��q6����[����D��6�}՘S�[��_�����u�+q��Ң$�/��oF~[k҅��	O��l>kR�5��c#hK�V09kM?�O�"c

�"�&�Ò��#s!�큓\^�Fo����O�6de�6��9y#��)��ٛ	k88��v���t~�����,O�����b4�~���UHI�v6�1����B�)��V�44���{^]5�AJ�뽺z��
��$���=�ƒڍk�%���͟
��B��w?$ڢ��9b�.�}�Pۢb^h����l���ݭԞ͈����7eX�f��w�0zO�u�����sL�1����)��r5똕+� ���k@���s���
Y�X�,�dg��W��v`3���BH�OAΥf��׼��_/oEF��f"�j�F4韄*���E�Y9|�ڵ��8��B�M �<i�=�����F�7)ۮ�Ο�f\������rv=�H�qg$"|��
��WD����Ƅf{�$%� M��-��!�rD[5+�hi�_E_y���nR�|9�𦟋�eH�	��"`3v���X�8��h��bQl6��!ec���O���EZ��׋{1LqQ���y}E7�{����F��]|-9M9����>쵺�#��^<�
\?ã칞�O5��#�-S�ݷ��!�R�#bQ�4�Uk����cQ�e�3�`���uS�4Ѭ��Ȁ=F1�>�
ha�� ����e�Gɸc~TM��BO3��FK���f>u��/֪��9��96J����D���a���?`������z��S��Yl�:}�!��	̦���B�'��|W�W!K ��J��̕�O��p�#������uw�U{^۬�:�k�λ��e�*�z!po����!�][�������q �G/p�@��~y�&�5��$O��آ D�J�ٷd�Λ�iec63WgW��1�ٿςO>o���J����N'^
Kw"�g��a�`Y����qXЂ%�my���MX��1�X�*�U+|	uK����#�Sy�h����JyW^���w��#;�v��[�4�����u>wg�^�(/�:r�z��)���,ά��;�����>�Xo*i�v�e���� f^TV(�̄��g&�U��6��c͞�T�,�̰.�S��H���kSȭ:~�'Y����|y9OW=��;gN%G_��æ��yv/tW���k&!|��U,�d|Oϸ���@�1���qi����`��P�<���R�J)��������\b���-��q�u��ey��~c������隍�:�~TD��=�����w���o�wT���k��籾�[Ϛ�e2+hw`W��wT���V��@q����
9��/�?��ݕS�>���at���O�\P�ټ=�7{�#D�7h����W��\�M��lo�Q��M�Ty:��O�XIȁ���gH����(X-0�8������� ���2�#E����
í^"%�����Ϗ"L1�_��˪^��%e��2�%%+�/&�t�L�D*��Q{';\p�s����f�fi�
L@fc#��$G_sf�c)Ph;[�ƌsA��u�@���GֽS��.�Q`V�?�e������_��V-၎"�6t^  �?`�����Te���,�X��)��u�m��&̗$s~�������bs�J%\W��*l���� ��Ӿ��C}�e��g�꨷J�'�����ܰӧ�!-H�ֹVtZ�c?����ʶ�G� A��8N����EВ�삀�����YN�=̼Ūj.}��90��\�(�
�UUCi��x�͓N�B�3���QhЌ�ۜ��^��H<��� �^n�������[I"7,5-k+�x����]�G^���U���d�������Ό@�|�F6�����S��G�ú��ܒʖ^�@D�Կ��˵�y7��^����D��q�ndSa��^�*��@`�Ї�D���
ݥĔp ���elսd�*&�>�@b7�U�t���% �t輸��@��<�h'a}��,��W 8�VZ^`�:�Д==�֫�t�������N~V����B���HB5��`�
�r&J*`Ë��@��B�Ɲ���l����v���b�n���i���Ӿ����ݓ��W�*�a�o\v�B��?T2����C���㰙��>tq�eS�����I�I8��q���]�+q�D�ƫ�l�������#�|m��y�0��g�Og	�FF����+��:��Tn���ӈ��Ϗ�F��4�nx���H��UWQ����{�d�U2Hx }�P��0^��oHa!U�bD5���,^T�A����/��ꌩ9�!��J����A���R�LZ�pʙ�s��p��j��Y�+E���^}�ՠ�x���U���Ն��)L��˭�����߂��қ����Fb�8>;:#V�&�
k�������0
���֞Η(����oh��J��~  	??��	�U���i��'�31����&�������W���JC�?�*������F�私��]���U���ve�%\�CP@&)m�!#�VO�~�z���XF�i&�S�m�h�O��J\'$��V��SYd�иˎd�0$�$y�#�^� �9�h~TC�-3��JY�}$%y�xL�F1���Ԭ�+���z�0է*��A�|�u�]��{{+�2���Xi�Xi��Ӽ��l-.��I1�"dȿ�f_�~b���@���E���N`leeeٌ�Au,x�3</�)�:�u�?5�=~��r[�[(YX^6ʥ+X����t�ktiF� ��$�ea�G^	P�_�1�\M`�럘u��7�PH4��Q]��1����!܆d,I��bٔ�樝8��e=�tD~��_��K�S�'�i����h�z�����*�����6�
��Q��?���ZE|��_zA`(�R{�L�ˍ�`Ħ����d�J���k��>'B�g	�����T��f�\���J&]�qT~'}�Fc�b.�Zqe�qF��o,�I��A:��c�r>[�y0WM��f >��L_C���m�z0͗lG���.�3�Õ����>����{i��7��Y�sEfmv ��R�qw,��ܱ��"��1A�>&V�3��Q��o��JF��}��;-~�J�EL<�-�Y�>�lhM.U�G�3j�<M�b/����x����a��R� ��U��H���V*!�y�'n_'/�9J�|��s	��h���)]���gN�Q�x�?~=Lh6v@�$��k8�ý}Y.�	FZ��u�;朧2��q�$��MG����a|� |0��������i�����QW�l��ѥ��/�uK.]0Ckeo0v)\}#��tV�X!ln�׭�4E�ii 	�_��c�=;Q�l��nG?O.96G��CT��r��)��&%ꚑ<��d��$���s�Q0ɋ��D���I�n]�=H�����|��E}��|١L���>~�p�$V�s'$E�d�?.)j��P�O�^.)< ���� G���S�_QD\ϡ�399a��<|@�<�-�U�"�|.=�7i��r8����KO���N���˩;T���?��\���4h�+[������T*�Gv���8��Z.����c*}�^��V��Չ�Y���J@�:=pz�ҌυAWm��d�y��v0v�׌��U�ʣ n���V(���^N��ѥm���7�2����_u���%>{�n��Mn��v'����S�����o���t8�4I�Y#�i�b�E��Ƴ��%��a�'�N&�V����h#��l�y��E������D~?Vlr}5��@�$�6?ٿM���ie�&H2�R���H�tv~Nl5x����Br����$>תCA��(��=+���p����t�A�^s<�*�ޛ�U]�?Y���`�RI'#���d�l��� ��şY��.~t�w׫�Z{��9��LɸG�Z|�h	��̒���:0>d�PR����[f���k�kY�]�g�M?OG����pR�������:��(�v�,'J1>-1U=澹�x�[4���D��j�e Bk�=� ?U�6uɰh������@Lx��IC��	F��{��A<<������\�Yyz��:��ߔ�����x}�#U|A�_B�ra�
"6~T��.3��V��#�'皧f���A�������]JN�A�}����C��TY�n�g`6VZ�}�]��7#-9:gα��.,���e���9�,�a>Sd�S";� y���b7��wC_�8a4?=��ѯ��嗻e�<�?��}*[Nm�zv�z��dbҲo��&���C�Qx�I�w#H�����4c�v�w�s�)�R>pV�G�c�%rf��8j�P��p����31UJ^�ąF?�⿑8����e���P�!j,��C�e^|�`���IF�8��ޮخ�_��	����g 7�y��a�4�^��:��]%�>��)p�G4*�&]�����}3�����隷V��i�;�1�d'ǩ��=T=���7	P�/6��Ƞ�9�p3G���2v^%��Z��T(I�S~ǳ��x=�8qpR��w��:��D�����I���'��ù�g�[�y�~��F�}3��Vg�#��T� r��� �ƎW�d���]s著K����<+I~�W+b�)���[�"0��޶�������I՞㞾yο�����4L�w����ῢ�+�!�x��5�����V������Sé�\ixv��`��)��{��a����VCT�A�~���E]5�N8ha�z/r�,�J��h��T#�_�Rb��8/iF��_�#�WO���Xt�k�Q� x Q�O-�u6����"U��g���G�Y6[�w���C��u�����]������6�u��n��qwlQ9��WԊ�'�>1"qE8�G ����.@��4r$&,�@hK���1�6u��~8J���`on��~|I;��E��O��[s?M]{ˑ5�I]=����4@��y������\߫q���/�<����f���솆.x*?/���"ofM�K�`��lK9�Uu�֤�����B^v蒓 ���}�����A�QۧI�x"�_���7*e�i�Nd��������q�3�%�a!��y�s+�um"YSUx��Y�D)��ʉN�c����а=q�f�閭�������$����U����ʙ����`"��V���!�a���mS��G�ElB�%�k��%y���+��2RK1��p����e旯r�]�=p�ߠM~��w�U����)��Uџ{O�\��%�V����n��� ��{�������@����FJ �a���Dv|_3�ƙB�R�(4`T�E�n�DR@���`l��\V��&O�dk|Ǣ���Cei�e�T�)�	l��	��j��v�{�_|�����%2Cױ�(S;qD�Q��R�@�G�O��wA�g���:
Q�O�����.��?����G�<yZu�{q>^���P�1�"�U� A���z	<��w�w"��LĺU��_Ơ�`rj��Z *!�eDd4�!��g-���S�nu�����!`U�sg��qp�x�o����z�rh��?�>�(�>��*�G?�����K(�S���0�eBN�X�!#����8��c�߱_���5v ���w�~�+�>��I+�"��j!�Ћf�'��,CCA���>��b�t��jq�Yr��S�C��+͚C���o����0`��9y�ձ��Kϧ_�Wc���cr]>���	of�G6'��w'/�QC�Gn_N�Y����8�QrQu�%��2*|F��e�'g���̸�
$��h턀/�Q�h�=�1wՖi��(�둕��˦ך�y�᧛t�U��l����4�wt6.S����Y�qW�2��ȟh�,j[`�!�7T��*����^О�yj�d�̲ �J�W��5�k�ś�����Œ=B��;6���<Ϟ`ء��
���A�v.*!�$_rڄ����Y�Ɵ���u]���/����f5%�\��-HU�]:ǥ};~Ĺ/^�m��Sވ9�}F�����ӷM$��%�x����J�Up?�?�w�8�g�+p�ȯ%��9m���);P{Z�	�JG��AL��E)4�!��K���Ο%��ث��C�c�9�| hNe�x`�h�Yu���7ܟ&>��be$��΃��i�;����¤��l�J++|gji��i<�����M�i5��q�k��S�7�XRm �`��l��';���"��65��]��p���N��=���	D.���'hrc����K(���`,hp�-�5��I��'�ضQ�
U:\��O�e^h��Nɟu����aV�%b�&�����ӕ�}d?v!u2mk�hoo/h촐�����Q��xp��P�Ԭ���VҖ��k�e5̝�(X³ǡ��ѥ��~R?Q�"���L�O�"��⤿���\��<�GW�l������5Uw�UiG��R���8���՝�](�37��u3���$ǿw���w���]��+IWTr�;������jj�v�|�)X��7����1�֤�\
������ӊ����d�&9E�]�{>�\��I m#M�?C�<gz�;Er!�X�����:��i&Z@]܆�A舞�����?&�����D�d�:"�`5���3�AQ ҵo`�f����s{��	�R��v�����k�tOb%Ӎ0��3�el�h�¨��l6��>��*�(�PS�����&�QP&U>DVA�nd��Q9��@��e�q��P�j�v�U[3��?cէ�D�Zm���ǗG&p�"C��[R�2p	�t��\@v$@���$�O��m���� ���xx����%z1"�ٷ��d1S�z>-f������	�Q�(�$q���cc��`m��{��� ѻL׃ܯ�9��uUN�7��oȚ�L�Yf4��]d �F�dm�������(]g�(vb����<D�I
Ll��h�����,��A=��U�b�Ra�He��?����L�<�QT�.GY���W@�{9�]�Y=��e�oF�~{���i�鿲m��*�����h0}Fh��2�-P6�-��|y��%I=f�ă��QR�ui�%&߾�c@������/����1���2����=�AO�����qWI�Ȧm�%6^9�O��r~&&���}�]z��0���j��}S<$�/�h�(�� & >�ƅ�����bW�7+PMb@]^�WΖ��>�۔�d�V�;8�X*�ӡȘ+v��:�5�#<�o�x�����6��H�j'r���U�Et���;������APr)�nX)Ab)	A�ei$�qD�%�Ni���}}������fΜ�9�9gf�y\Ek�9�(�j	j��:�������Qf�}��|W�6�"6nΗ<�.�E���9�W54��ƭ����U	FK)KN���Bo���`�8h����d�Vl^)�8w���o���'p%�ؚY �M"���i�׭߷LjM�;������+�Ob����nc��H;�/.�$���GC?7츞�L,�m��}��S�W fK�5�&�Vw&�'��bK��`��"�� �'���2��XoJ5��h��q#q(�����Z�C��﷾X�k�Ct�o����\㼘_=_���0Ȝ�N�l�z6B^�l��{x�O�ठt���W��"rq�ĎϷ�*�!]UU;-gx�݆�`)�@��(�D(�U��$^|�*��͙����}K��B�վ���K w��βg��6HL��3��j��fn��r�|8���K��/G�HD�Q��x�VM���Іh�=���(o����p�>��H$#`,�r�H�Z2��8��2���hD*�q��Mbzln�Y
z���C��f���A���g�ò+�rin��,��)�`�n���_�T-r�<���V�Ŭ�;����+�͜�4��xll�D炂�S3�F
4��5�l��BB�ܛ��#|<C��������\7�P��y��#������� �l�y!\���`�����:�d^qs�y?��|�����R��a>FJ�pϫ�_���L�W��RG��bM0 �e�6��άĥ01>�`3�PرP{~ �]2�^W&Vp������8�r-G#����tO:��ؗ˛[9$)��].K��ż�v�P���PkZ�0�,�6(�Vy���6b0�=Ъ�Q��3clj]�p9U{�
����e/3��|���#u�����A7����:5�_���*�ڛ>S�3[~Z��?i�-}�P4mN�+�ͭ��%�V�ZT���������� �^�T�,c���7F���*��z��ej����M�����o�����f���	�G�/b�k���p
B�fK���DNX�V��2�����mf������d��(�I�H���2:�`�)�S���g��.7`�_v��;e��!�߲��>V	���\�v�ש*�I|�znR�B��g�;�4�,�1o��&�T���pU���������Dd~���r=��$�z�}d!��|Fw��R�W��k?8��os�� *��3�{���-O�A���u<M�r,-?���)����Y���-����;�`B���^Y�l�R��M�B�9���l��l�&h�k��x'������Ň�Z)�:h�{7?��_}]Q��R�����G$�]>�XǸ�ňˀ
� 17�1�|���P"�"��cji$��0ꂬ�cd��%	��zqa6�l�}�@���ZM�����؁P[xa0����-���Y��* �ƣ��h��6����Հ�܈�����ɶ����2]�zn�����JQ�TJ
	y$J��N[�OEa��֤��U��*H��;S*5W�����QT�Q��w��vj.tqڣϊ
�$��# t�;��$�(t�����e^�	S?_g��)u��6ܶ3h�.�j�~�ձ(@�G�W���M��~��r��`	1��X����AZOb��7r�>��)�w��]�N�,�iT��`�E+�fT�V��1�p�������|c���חǨR��;k�-�4w	:��� �[e���F=�����f�y�]�a*�Y��u�T]���FgN�笚E��h�&dҟ�.�;���h���~d<s�|!�� T�S�5�u�Ib�	�Ó�l�^� ���g�3��i1=%�;]�w�B2y��0�m��h�y1����_��*|��@F�o�rɭ~R�K&E�n�LZ�=�m�6����v@l��}��ZS���4���~wP��wN.泷w=�=��f o�����`��H����k4*	Fb>& O�o6
y���O��w5�
42��K5����͉���� Q/:llETE�PK�ţ� ��Ӹ���అ�iSu9Cu�q8p��wwֲ%;�S�t��杍�+�Ώ��ҙ�:`z�X����N�ԇQ�j�֪�� �]Nn�QxP��}���ܰqR�}N��/�>��k���b���i���������Yk�	�g�����w��ᕕy८��f�!���ϟ}t9)Zg�v���5���O��
�%;$ؽug���9����x�	f�𮱰�k+�pH���w�J ��ܞ��zհz�b��֦������o�t�=�mU���*���fs7j�Zm�0?��!��)Sʹ�f�V�57�E��-u���375U�B19�>��!56iM�x��8�*D���T<2x�A���O�	���Ȋtn��T� �#���S獍J�H��ܫH�;��4���c�a5x���$©�[_	�+	��0Z [��d��St�~_�59@�ȫ_r�Uv��'M�8>f�ȿ�H�J6ڟE�".0iY��&�"V�J���nR���	I?:H	<�B��v�hnNU��ii*ɡ�e<��?1;���pQ� *����fi:}��9���GWW������و��}��K��w�g�&?�_˸�w��5&�</U}�6�C'��Ic#������\��ε����l�
�|��!����b���F�W�e MƼ�/!((�0Q�ϱ��o�]:�k����:�3KϯJ|����dl���3��n��N ����9�_�T)P_c�p�IN5�ˣmZ$�o��M�l`��N�;��.���B���62��w��nt����b����Rhq>&  �C@e�c:��utt6�3WD��k10�\�'���
C������??j`�)"�ޛ����r)隃W!���|<>�љߣ��u#�_{Za�q@,��V�#�'�&�~�[��ϓ!1�q�9��$�P��Ҩ3@��3S��^���45�aI䡠�&MZ�Y������[&CB���:<�^ݯK��U�Nvu-�+̝��a���qQ?��􇖚�\v�x�m�i�"�w�8�Ƿ�ʾkeڏ��j��W�{�*��idK�P
�T�)8��[07R�t�=b�Lޛ��n?ƕ�N����WYTd��/�|sT�NӁ�	p���y�z��"�Wt�cPֱ�<=�����*
+�$��_r��e��;a$bz��)��P�f^+I�]��[��
�����խ��ߡ!�[�iesS9H�a'�*��m�c'dK��P!�S�3�4��O;ǌ����.b`$�����!lV�X����[C
�	�iC�Ʋ`�6s�1��S|����G(!!�!�9�¬$O0�B�-�������5�M�z�;e�����6���IH���Wv^�Y�w\�[Ӫ�*-<c�F|&Er\`u�:\��=|�VW\lwH��������nJ^�Ӆ��\���w�S2P����+k�l�@�Xvc��H�I��{�d����'ϰ�oHt�G�S��~�l���U;�Mq��uq�3#�3�?�lmzJ�Q$v�ִ���X�l��?�H `�����h~�s�+C3�uȟ�kS���?x�?Im��Ō|߮�����;����!��Ti>Is_92>�ό�E��1��4%���k1�rB��%��ԙT&c�D��uǖDKk����~��pm�[�k�\f`N'@�o(�#8���8|�x�BlHq�^�Zn�eT��dڸ�G7�XS=b�{r�?��T��ӈur4��}2�
��[���?��uB�!��)���|�r�-Q���:]���͈��0m!ܖbx!a����� �?���	j}i���p�E�wR����~!NqKj
��'�M)3��*ϫ����AวJʐw�R�p/q��c�A?]́�����.�0�w��]4Ќ���dE�En�J��O���]8%y]]�'-8�4u_ma��~t�����5p��~f� m��s��!@jS�h-�o��z�����߫���ǴL]w�ԴOp�z�܂h_�/����G�����tz�;��٪�_3���d��Ɉ�i
-��N��P�3F \���9���t.▖�0}pZxv�.-Q��j^նw�������R���t *����s�C�]xD"�qI�[(����l��"�aM���F�,h�>U��4�BG��q�Zt��T�Ӵ7�����>���UGi�;DV�j�,Y�#�:�ҝ����FFFA��_k"x� tw��n���;�������x�9$��\Û�������ƨ� ������#��ŽNv�����׵��^��W������*�h�hrFD�E�ǅS�ק{kAF���At��rH��,:������F�N@�2�{�[ȳ��ၚ���Zw�&7���b���϶��Ob: �{D�� ��4~���L�O�5:�;L<����,�h<����?�Zh�b=9`�?�9�X>�m����  {���?�C@h���l��O���$�K���=�kR�?]P��m��PK   ��W������ �� /   images/8db8bc11-a89c-44df-83ef-15ccf3dbf879.png\�sp%L�-�9�1��<�mN�	&�1�3��;��m۶Nl�}�V�w��ѫ�Vu���]{��U;BEI�	UVFB����� ��"�����&-Q3E|A!+!��ip��M�����Y��oQ��ǏTSX�U��C�!8[#��t�Qh�;s8|V�`6�>h8�������h��K����/����9T�t{u�c?�����=��'Ιwc8_����=ӫ(t�HY��_��#�<�zfLo(�L'�R�u��2���P�Y�n��T�\P�`��.�_�0RFH3_0�{�bz� �'��F�����"_�-�i��� ��?��Q6�)��PޡQ���-��9J��w��<}q�ǩVÄ� .��oS܃�
�����N�1�]�5^tgLb�M2��ፔ�����y�T%�I<�Õ!CW5xt���r��"B�:�$�,2�qs���6-�E񱉇�D!&,!3|"�7��P� YV]���� DJ��?�5�u;�!D�*�uA��Ct]�7χ�#�M�L�,��R6R��g�*�|.��~�ݟJ�^S�i����Q�~3�v�y��ص�<";���uW2PU	+ R���`����#A�#�x4U5a"��a4D,1KD4aCj�#���*"U��"�kf!P昷_"�b0�Ex$�0A*��Pe5�H<9�c)����Z?B97��a��3�8��jr�nƺ�˚ �xt2�p�� :(�px� W�Z���#b����5a:�����e��tlܜhÇ��1�֬>#�I�Y�����XS��"����0�d�1�"Q�[e��I�س�<��a���I	�1�Ԝ����"�"�o���E�;J����b�R��Lx�j�
�u�5$?��%Q@%�qp��ќ�� ػ5�I̈|�Nrz�|�'$�!{F�"co)ub�ɷ�b�֫ %�?L�,��D(����}��}l���~x�`�E>��������_$��(�8$���Y�ú��<�ƳؠN9J��w�55I�
)yO�gQ�Z0��b~7�5�Z@Um����;��<'�O�Z����ۡ�@U;��镉��m�J�8y��1�2~	��_�V����Z$�YTu���>�r�T�P�e���NIth��8�T3ݘj�׮����08���*6��!v+R]�O��� 
�px��p���[u��8�[�~�
�t�����I!a�h��s���w �� �D�\�~	�EH�\1+� ���#�*4�z�@�pgf� ��	}b+W�A�م}Z��3��&�VK)!YF�D���.�,�_fM����@�=��2�O	 VF�_��Ǧ��t�(�C�Z#��;#�",���1�-	$����#��T0�a��!YG�1<��<b�i8C�|K�u]`@	|$��&�������fLo\�&&��oJ���j��!��(~E �e���8�'�|-BAC�Uy4��B�gB�:���)(�m�N�D��J�D�Z���d�G���Y8��Zh$���J�l�Tu#���!t���2�d�nN�0�Ua�V�����>BP���I)�g�ZBl���h�IR�L~��ò��A���T��q%���;�n�A^��
�3��|��	�q�@�!�7��|*v��x�A���
z���&�,_��9H�,�L��*Բ�����<��8 S�ȵ�5�qݍ���*���Ο�O E���'4�Z���?<qs�g��A(z�ۧ��m=����Qf}�O�Rl3�Q%�ƧHW�ؾVg�%���E%�t0C����{�~�e�w"I}A���#�P:���'tz�%Eb�ݳYi�n���,�,cDק�N��\D���������q��ښ����6:Ե%�����=�ɹV�������Up@6q�ܷ�z �9�!���������}��+`(~�`�
�Ƶ,"�8׈��t儢��Pӣ_�	�N�)m��u.�KaQ_,��ؔ�*����@HQ��A)�2���9b�ϠŃ,� Zcր��g@�Ԍ����e	H�,�mw)Λ�*��MG[�m	9,\�?�lm�S�de7��W-V�4��L��2%D��5Wh���߽�z)S�24�&L�5�6�E0�\d�o��L�8�9$�9�����q9��:ؖ�l<�ps&7D��7/1H��y���� �"/�"��
�O���u�a�t
+��@#�L�H?�D�V��PBXB�U�PSBׇ,����H.��u-�SAh�vtV�����ht�Sj���JNjTp8�;T�g��� ���-+
⦍��Y(F*��Swa�l~d^��qqU�1�����ҋ�� �-3��֣�#�P��� �����ah�
����Tpz�̊B�*�s*��M�� .E�u�6(uTΕ��q璽�BIz��*"8u�
���!��>�����ݓ��LU3G�7]Lz��	���xI+�Y���ID�}� F
�g�$	r1�D�<�4�AZ�*?���`�Z���q�7Av�/�a{
�>��q2ӹ�d�.�����w#�O�'�ϳ�'����&fq߃��FhP��E=f\@5��������*["�08e�F�?��|�E��Y~� �����&��]M�{�6J
VZ�.�)����+;�`i%�SL���n��<��	5�:��
+Q@�i�R8;�+$"�I0K����]nv�'��
�o����£�(N�h@����x��J�qs�-VjVWö꣙Pz��9.�V��X�:~n^]���;݄���1�v@�/:�H�^4��H��ՙ�Md�a{l��OgE�2@�'�ik�f9]��95\�W��o���b��!­�#���O�u�@�uo:�G"�*�U������H��>>ѷم���|[�霏b�C�kS����8���tu#s����i��\�<�u��S�^������cr/sCo|�z��h�_���6�z[X0�1�� z��t�-�L���P��ƠL��"��)'£�٠�E� ��WK��&�n9��,���� ��`��ʀ����d	�t)�2%���&^��UD�Y�u�9+'/��imk���&a���ϱ��Lp�����-O'��ߘP�Uc��;�84�*��0�%[����(��"�f��[���Ts� ver�3��I2�٠̻�'f(?$$��9ZQ��
�*E�/so�2��V]fz��|R|$�~4�u�?z��R!��.s�h��b��b}ъ�'�}~8��4�0���T�u�%l�wn!]fmV	����ܻ�L���#����=;����BrD���Y W�T�퐍bĂ,�����Qb�! �K�m�7PG��V���U|��u{A!/��.� i�����S�z:V����+�H�j�?`Ap�RPk�̬�ͦ\Y�k	��n�"���
����"-����,�)!�1�.��M#�0Zi\��^�~�f�߲���Ň��(����_+#O&�?h�k�2g`�l�5�54Q���Q\ſ���������ҧ2�2a�j�
�B@.j��N�_Lk$� ��$��B�.�!�|�>(�p�����T���č[r-~\�}�^����5ӽ�iFK)��Z(!|�kj���KSu�y>X�H��!ܨS���B�+�����Z�2-���p���e7-�*�дŒ������f���v9"�@�T
�H �b3��L�H*���-["�o�,���*��k�p��y�f�M���9o��_Q�ӕ�`���s9�����|��;I��2��p�7��1?�G�,�N��a�?�8(L%W�YO�N�x�s8��|���w��K&f
��C/T�p^X�K�n�W�����A���D�4s�t��n�/��][C�y��&]�z��/����xM�2�2���mA�B ��(�iߓ!�"�)1v��-���a} T}s\]�ٲ�^��R��^�Ua�o��Z(l2��M�z�2�ׄrC��-
��\b�ݕ���]s2��K�(�$�cK��Ɔ���2O0��Xhewb9Dl6��3�<��|�3Q��Z+�"6�w�TUu"��[�y�0��BIXr�!2�Ȏ�֗���T"��]����π�	I�u-�[�܊?(G�l�E\HE�ƌ�H�mx�<��]����t.%.Ne�}�e2@�gp?�
g��gHAZ��&+q{�)h��o��p[�	����^y|e��w���F�ˤP?-�|�Tm"�z[�/���>����w=&�R�q�ZD�r�ƭ��
�����\H���Qs2����)��=����[�>Zm��ՖG�1c���n{(�����Z�������z{E;Uj`��dǹ8A����9o�pu���}鷆Tۨ�갰pT��aU�-��ö�Jw��$�o�$��ppp?��a��4�Æ��9���/�K��B�dkۺ�M����{0̰q"��s�I@�OaQ>Rm:��n��B#�TΘo��||s���:/���sT�w!�T���x�?(֝��0�{�s��1%Z'X�R�gk_< )BJ����ҳ���a�Sp!,9�#���"�]�SԆ�%��|iu�������W�����Db�ŧ�}:k,��P9�.��H�xⷷ�:꜄�H Ӷ���/~tr@ج��#��ؖP�F�%�tʣ6�TǾ����Z�O��k�or)D���*cQSF�w!�D^�A֦�#&��%X�]󓿓��1"O�jn涛<��RΘ��w�!��}�r@w����7;�~$!�Ai�-k��d��S0��q8uu[)@d����K=<:m�Ua��"u�:moAף?<M/���G�Z���U��T�̋JG%F�;���A<��S�N�c�C��7`��T!I_hf��[x���g��D�f��
a����0[�n��Z .�XTY�Ѿ��<��ԶJ�ʾ5@ϡ�㘹/�����`z�+���U�c��t��^:[=|�Wi!�r@���As"�ݽO�&ɸ�P�a����׍�Ӆx�;����+
/'�8�wض���l����Tl+^�><�Zj��k�V�7QvJ�062����J`�(�<�(M@�Dʹ"�ׇ��i����0�C��Wԟ�y��0,�C ��2��}�SCz�)uM��ϘAJP�܍6G��++-�F%ڐ�Z�,(��o�{5�&w7�E�ǰ?�p�hS�?�e�c���Į���FO���2�+$#-�\E�A|�/����'�b���>���ӯ�~������G I�ԥ�� ٴ�1��3��� �E^�<s��e�C��/j;�L��t���+��ʝT~��Z����fȤ>F�]ϡ,;����ϖ����<��N��Q�~��-7��C�.����,���do���%��:��(Ý��������Z�r�$(��~v�C��N;��<>q��u���V"V�<Y��F�+�~�V�w��;O[�f�i�X�.moDB��JN=������[M�����U�TP^��T�����y���0<V<�4�������V�b2쎂�nr�ָ�pB���H�T�G�����x�Q�ϵ�i���!�Eo�a+�~�7jY�DY�_�a�O8�o�[i��.�Ψ��2�w�6F�~BN�CɜWT��'[�LXu*0��n�h�x�R)�7&��Վ�<�@�N#��УDq��#wYk�i�*�$�#�7P�
����aq
o>���%|���(�ʒD��g��W�M�	�������v��������~���8L>��K�2�^�'���Ĭ�(5)-
_(m�>���6YM��_�+Q <�H�V ����B�:��.�AlQ%Ĝ�θ��O�=�Zl��K9x3G1��E���GE�>߁�����ȯi�zG�L~��N\��x�hQ��
R�����yM�E�^��鹧�҄U��OE�Vr�b-�!���G��f���z͵~;	Q�C5�Ѷ.�_`|"|��?�D�銯�^	ΊD<h�l� h�T�o:L��!�E�V[�N�u�R�����y�\8Ub)=�����'�gf���G���
�/xR�I��7�t�';%Y����3k<��_\4U�����vR�6�G��)�^��5+Cn�,�|�8
�xC�+ɲ�[�~�.ٰڻ\kD�j�,��M�7���.JZx�����k�h+l�-����BW���3��(K6��zTqx�B@.ɗ������_z�ܜ}����r�t���R��e��"k��i_y��
��#���HH1L
9���ͮ�[;�su���2�y�J��5v'���k��>�Q��$�"K_/pGL�ꨁ)З}�u��r?��^�]l��?}�<�	[�.��D�;k(���(8%�C�`�B|%��ՈWx�eik���/�췾�f����s�}�cBɰ����{����H9/&aW���/J�J���q��i'���L��y?�������N�S)t��􎹇QϠ?W��Ҧv��߃�9��`.�z��OQ1�,-D��Ұ��HPo�/��]�r�iyb;���L�>i�p��Fd胖�y_��rx3Bg e��#�Mˠ����^��$�n��~g������a�w��y�7�ꆾ��&h�� ��Zsf�!��'��L�R���-׊k�1��]v���9��z��4��Vv�M�}�Ods![d�b��|�=_K����_�*�:cJ���98��\�=���ͅ�+�z�|�N��2g�ׅy_xtU&���?���a������e�La�K%�Ji k�	�G���/�%�+�i���C��oI7@P������H5M���|�����6Jgv*�ҫ�����a��V�$�� �cI�}Sަ36��9��F�[�r�̩�th s��˝�a���Yq�W����R޴�v����*2��[���/A!�y|�2H&��ɓH�_f`A��]k�o\Ư�+Œr.��"7C��������>y��/�����BU|����q-�R�,Q��:tN����&|O^�cݥ�ǒ%��4�b!��[q��� j��Zz#�v|�l��i��9�U�U�vE�P�d_�F��B�ˣWm�g+\-A�MBWs�H��I�a�&�� �*��	Vr���\gBFs�!�B�pX���=e��l>�̜��o���@���8.V�K}��+��.�&�eaՠVSܟ99�^`:�y�Ubid�e�h	��a��?wS��ïu.O��NC��C���;p��w��cE�tPmz�޵�p�Q��T��^�zMv"薳�j�*w����N��=q���B��?{�ךv�q4�~�W%�(�Jϒ/w$�e�4�=���t��:��f;)�?��3#��������>s��m���,)�#i��ɑC�9p�%�Y�ոH4��Ήv���wC�Y����};t(�xDq^��5N��h�v&v_����|LemҦ���m�p�C1�ͨ�;,��Y��u�οsN������Z/Z��F$Ï���Fit�������Kd�����w��{5&g�萘72ݸI���8�s �T��O�����Q�b��.�ph����X��ڟ�D��� �~���f­�O�ٹ����u���Z��Bj�4{�+7������i_x�%���TB�	�{�%�������z�fi�a��5�9�&��$�W���Ʊ��+k���Ni��ɺ/��K����S��چ1�oO���P<�`�����?���ǹ�!SG�_�6��C�u���6r�L�N�5ݻp�
g}����y�0x�^�Z�BD�ݟ�8�:�z�A��ޓ�v������W����WW"2=���0��齔�	"|�
��t�Q�&7���*TP,^�;Ed���_�F v�6��rB��-e��̩��am�1^������Ab�c*E�s�?�͕�Y�ҽ�z]7a1��t���d�q�6{dƒe��H$Fh�o�]�_4FaH��+ڬ�6E���3��2O -!I]X��[���R�I�=���uoT��� ���S	�]�˻�Fk��7}�`�`Ps���EH�n��������B���j���73r�8���
w?�䡧�s~�[�,��H�x�(|,���
>5��xU��W����I�??���>�!,�O/��ݗjc��BK=!{���7ơ�I���t�X;%�����wa��D?chi����T�YL0=Nn�wx11ɤ�GKZ����P���q'^�?&T�����0��@�1�x+ˁ���U[h�M�V�c[>�2���\�[���p�r����k��U�*�L�%��>����xq�� k҈"X�y�M�}�/�{��yG�Ĳ�s��fe�̷03�*V�H�yYl�Q�/<6NΞ���^W]��� ���r!8�Uѕ�"F�~�2�'���U�i�L�۫�9fRaoT[,\t!�q�D��F�.�3�*���ft�Õ�AYW�N���A�*ّ�{Y����rO�-�-�w	0�{AM����'��@f�҈-KbA�$�cn��P[`�ɇo:�	������U��b��#��������q��+B,)o���f�;�.2OHɯ��{���8㳥�����=��_C�`K�^�/��;�^�������h����ӊʿF�>��^7�>��y�'ߟ=�BL|?,�m���5䇣����a_J���X����?M���&�w~ �>�&r��rҺ@���M�j���l��Ky����L�Y��O	��'t
����,Kb��|��=�y�^�Wn�*u<�7-��+��I��^�/W�)��¤:�o�u<�?<�5�����v�?'���E�8�ק��{��l�>��U@�5~�t������f�(�WPi3����Bd�9,$P�`��G�*�Qy��X�Z�*$ٍ���;�\�W�H�N6~w���	�.��)��SÇ 2�l�C&R���3I(J�>���|�s6EҨ��(cfv3��k���?���Lm4��΂	`E�+Y�#k��[D�� ��ٺ.u�1��S��c=�-��م�:>iL��X�a�E�~`�[��݂��z ;�1z��M�5&*A���2��̣O��*At����K�a�4�z�3F��ۭ���L���+k#XeIJ֑����,���LduJ���ҭ�R.�Q� ?�/I�;)�ŏ��i��Jdeö�I4��n��>�<��,�������$e��k-u*A����D���wjI1�Ļ�����(��-��DC�&L��hTP+�0�%��q`>�on��C�R�E��SVE;]���������ǒ�,"�rk����ggV��
�� �B�t���
��Uk4��w��Pm�ۼ�l{w,I��HDF�f�]����0`�0���v�zZ�,V�X�M�L ^�EWG]��hU��g%�9��K#c�9�	���a������f�@�����+A�a��ܤ��ߨ�":���N��e�b�Q��w�,���q�vd=�b����啈�S0��UȐ�/��q�u��KGe�s��r��������e8.�q��PX�3�����g�����%��N�Pe�@��g�BukQ��<�p�Ѓɪ�u�������ml�����[��m�)~����(����h���?\�́�G������B�h6�c�5�y^fm�;��Vn�u���ɸvϒ]�뜇o���rX��n�o��|T���l��5ƕN�Ŭ�ר���~��ʎ�i�-r�)ҕ�7����_��B�����@�5U�n(X�#^��$�03��	�A~�]_o0|��el���֨B��
�����\��B�cb#�v�H9�R��z�4�VϹ���s������l����E��D���:Ը��z���zp��5��/���f8���Z��
+�Mоl>�p�AbgZ�B��m�+�����r��u�@}�� �_9~�Wּ{�Wg>3E�^��Nŉ���u�PŻ,*KJ̖��2gُ�ơ|_�7���<Q����h|N�y��!��l��fDBz}��/�R��~ѧ`��sթ�%�Ii�>4�j�i%q��uf�xg+�[Cݼ
��&z>�4L�ʪ����e��EXB���&�5��m��w&����" ]�Eu���f�����9�w��
�q�Soq�KD}���F���޶���a��6��q�6�E� �v������Љ�1L�Lj�{^��6������O�ku�vs��P���u"G���.On��*���ߪ�"A���d�eai>��'�\SW�ǿ�L4G���y?q�r	�� hI����|
�^mvO�W��*�
H�EJ���%K��@��H�����Bǫ�s�b'�z�f&l����Ɓ#�H��Ō��V��ԇ�U�)W���~a"�ݳ�N�J��k���6U��ɮx_gˁ�Y��ILưw�@Ī�`s�LbJ��h�M�U�5�+\&lR�/
�	��BrOv&ި/��!L�PW�ΖK�2`7o�(�+	���׸V�c�g��g�!�x�h1) �2ɥ8O���(��M�9�O�9��ޒ �a`�R�{�{�T��A)�X��g�.Xu�L:��a���W1�wy�t�x�O��"�?����m����VT1�ʛ�&������5T�TjN������V��DJ]�uF7�pe%M^B{w�*�~�.�M*W�� ���2Z�UGl��������<��$5�dio�'c!,���Uj��-OƑ!EW�hFK� �k��|r"���F��+
��,����[��x�%t�#^�GPTTi�����-�l������Ff�=��v����ީ�b!�A�CM��m=�3�̾�Z5Fθ�1g�ܣ��n'��-U�`��ZN��Ӊ����#ȴ��D�S�L���2Y�4}3���UX�iZ
I4E��6�ʛ�F2Vل�SN�'��Lk�:��@����C����u�C �����Z6Vl/(e��)N��oUh�WS�+�����$�+e���?l�}��u��|I��k�TNA�\FZ��W��_�H�w����qqE0R���Vb�U�8<h�:&��DLo5��Z����R}k�kܿ��#oe�l�W�
����	�\J3+�Qd�PA;��as�ƭ��s��PP����d���q-��I5������7�Cލ�����!2ߔ$��i���,a�e�:N	��>�ģY/�D�_%�kil�t���¤&���!�׭��'/��8���i�u�,���=�v}z�K�U�����He��YL �S�g@L���R�����9����Ðj���vh���;όƦ��-�U�>Ӎ�L��uMA�&���X@A<4q� �k�?[v��H�%߷��"�^|��H�����!�gI�q�4qĪ5R��B���
���b�c錶[��]��D�՘Y�4��mJ����!Nn���j��S��?T�%G������+o�ћ��qT<_o$�gQ=*W8m�}k��0c��N;��� ���FN��O�a6���\�&:�	9e���!\��Cs�|j���![�$��<�(Y�2O̾B,@
����߿�)=��74�T�7�0)S�c���!Fn`�N���)�ٔ���8E��稉�2�R��5B¥.0�D��E��,&��O�E�:L����W5��2%��j*b%ؼ����jDD�~�8۞!ZRH<;逭�%�
��q��ƨBK+�X����R�]"3rG_t�m��L.�x�Sm����$ͫ�0ю�g �& �x̵���������ٹl�<�Ǳ�4����+�>Ӱeio�;�$���[y�a�;e0�����@�J�s��Й`"�{P,2g%8!�W)��O4��k�&����k���J����t�_��X�0�%d�P���aRc�B�9�Z�GGC��I����:����������H�%�2BJ2���jcɫ����K�����O�M�����$���!�D�Fk�F��Q	Nx_���en)�*�쎗��8݄&0 �edJ�'��v��U���K@�.|г�>�/,�!1�R�XIb�iF��ʅ!2�6�^�|�l��n���Z�]��[�K���0z��ko{�gGȫߕî��6�N۸SZ���:\Z۱��`Z����r�Օ<�t5���J�vo��̑�;�鸴���F诽���z��'Y�~�xx���%d��}����淣{2�\�K$�V���j;�5|V�k�_D�06�0��~��w���K�
2v��.8�L{I��%�)��w募{K0(��b�&���1������^�d��m+�U�؂)�섚�#Ku}}��#��UKN��h@J�ï���P0H���V@�_�̧�ʗت�.�p�)E�����8��̯�Ǔ~c�E�~�Z����"�~���#-�4e��|��@r[L	��OC.����ngr�{����Fw4���qg�c�s6�)Dbl ����TV�-���%���9�Q)�m
>�H���h��Zv!{ pA�p=G a��*�H�(��%�t-7�Q�ȫ:��jc�l
��Ue*�<�B����B�2<�E�����*�19�T5X�%�Y����'�r�T��*,��Oϥ�sP��Nd|����!�PA�1��_������v}C�d_��Т�BQB����\��{�Q����8�ܜFǏ$+�,�BCH�],��r��¨���b5D�wpp6K	�]���D�ʞ�D�9�q�$�-��CsG��;k�r�T��.���I�_&}ǩ֍pPy}L�MD8ioӲ���
�4���ꈪ����ˡ��DJ��s�пF��GG(Ζ{���W!p���-�VG�Ӎ��}��{Ц�cB�or^�|d_��������/�ˮ?�C���x�ڌ�h@�rαPʸѴ��q�T����m6l1#!}&�i�~�^�Q�M��rB���h�����%�mȜ�y|Ś��������E�c���� ��җ�0��+���� !{3�c*!��:qe�4���O;۹�����2��W�M�^	�`/�2�Wx�a����{�"aJ�Z �%����;�DB�����`s�ן~l��n�7�2�wkL�����?�x~�G�<��[M�տ���m���o3��d_�]�T�Ch��tsٲ�����4X����V_��U�	�~*����k��>{��Ƈ*��Ȕ�PRux%ɫ4��;3�ކ$�S�}+i��}��]���^�bw���'��P8�5j��$RP�M���Ď�%�߲ �&0��#��9c�b��E��#Ҕt����?�{ޘq6#ƜZ)���	2J���n�Zr�|�^�'�?敠�E���N:7[��Y���K�V���(��g�YC���q�c�g�ύΦ�[N��g���>O���3,�_`ߟ��O�$�k�ͤ�2���8�$ߢ��?ڤ��� }���mf����p,�!�l�M�����wBOH
8��\��}!�'^x���$i������x�n�=fM�8L����t��ʃD��n>j!̇n�A�H���.��K�tn�"�

�m��?C&�)�]I��'G�n�<wP�}�Bg>b�/Z�wF�D�w����V��ꨪ~�R��JƫA��_��]�"O�K8y"1`����l
��#��%�L5NS�g�6�vA���e���xSC�%ԑ9(ڢ�h}�?��?�KjT�9g�p Z��u�nh�r>�fy�L���}H[5�3%�]/�����ْ�4�5��*Ɣ �2Q�L��}�\c>�ԡ�\��3�LdJ[v/�{�C�d�Y��f���T��V�`<U��/5�"�Y[���W����qu}0$���6J�k#%>��-?S�xL�֙T�b�}�8�8��qgW���ׯ��3z;m���T^�׸��3Ͼ%7fK�E�5�#s"X�b����+�GK y�R(`�p��h��Q{m��u�-�f�R'�fK�� �<���*Nk�+X?�p�e7����+~Y>3!>1���-��l0a��8|z�Ydk�	��~�S�6���
p�O���/;\NRs�[���N���{1��\8j4����,��B�Ci5��o��;�IP�е�?_ϼ��w��J�p}�O!J�btC��UB�3�~�;2d�~�a̆v��=e�}���~1�e��
� ����h���<B�(�<�1�|�!ei%I�;PvjA�!�Z���ƨ�R�2����I� ��Og�y�`|��DV���-�L0yy�|�ڛw
ɾ �n�O��D��B�E�8��j� ������	�9a�$�\����P�ow`����C��~K0xТ�Y�4�zn���z�C`��?��(���j��nO�5����
O~�ʂRn%�$+(	*�E��Rr�&�^�ו�fH�qr�������]���cQ��+�ֆ:_��[)1��p�%v���Sl��@Q�����Od E{�;v�W2&?�y��O�wA~8U����<���u*��]�F�(��_�4�Ƈ�2�	��Wq1.��-Ȏa���>�<y-
� �i2Ae'��c�@Ͼ8;T묈�V_"����j5b�s������n8��]m���Ƥ8�6YQ\��F`=
��윟�8�f��
��ϖ.��)��Y(^@����p��*EH�4�b-��pEw��Ֆ��f��$$����HD�H�繥PP�^�З�s�@_1R�'���	]���r$�y���Ge-�1�FOtKm*��ΛW���-�� ����'��P2�,8�J*`��9;�=(��B��l�:ɦ:	�!���]�-N- ,o�Wa�@�ŉ���d_F�#���{f�摞����T�@����M�� �~x�}f�-q�/��F�%�UD�A<:�������J9�T�m�H���
CiΪ����\�����V�h�g���p%�:��ψ�����Y���¯�V�5�Zk F����ԉ\k��}��SF�w�H����7u=k(�����Q���H�Kh���]��9���R-���Z�g��.Mָf���e ��G|ӥ�m�.�Z�+r����L	
�}����M7s�]��ф�qQ��WT;��m�����yEvј&z�~)M6;`8�Gx�q4׸��؇�����	]������]�r��39S��J�N0C�NK�z�v)
�Ɩ/�O"U~Aٔ �s�:��E�G����b�)2_X���`��9��<&;�yPU"�����_s���S?��N�?�}tw�ԝ�M�&,�`��m�c*;��O"�d��R����I�5B:��4~���V��ؙ�����	�Ej]b���f�3U�Lt�Ȱ����߄�q�,q\�|���6�P� �hR�F�"�n���L�F'P���F�x���d�x8�G���(�BY��r�F��"�/wcz�<�7Tҕ�GA�⟹νW���#�:�rHRHI꽄C/S��ԇ��wD�}3+��A��qJ��eh{��M/h-ae%��y��^&���y
w�I$��L�U�הﯶa\c�DWFɊ��-2{8�2�vGV��6FӒv�K?]�DBl���Q�_�B�ըb��j��	�x�-J-%|B
�Vށ؁�y")��H�`]�'H���V1���I��E��huiɢ𕶳��I�2<�IK>�9w��R�>�U��vIȆ ���Ȫ�E��k�Az��H��"EI.� �f�f'Xɳ{����\��
�C�
�m2���L*D�}̘�e&�p��ߵ3T�EJ����)�L�Au�U�4G��P�r&_u�k@��W7��
��c(����d�L|���4���#�r���N�I}�-C�0U�ldA�]��}`�~BɄš��E��Oѽ�Q��y@;Q}�䚒;>�4p�;N~��M7��;�eq-v&���[~OZ�]e:�!���􈥵ա菀�.�0��Z�NJ��2&#�PS�$�sS�/����d�Hγl��Ysb$���y�G����U;x"ǟ��TЋ���8˖���z{,Jޯ"=�5zYoc=V���K�ʖ�c�������/��0-�7��Oǳ~�����EXe�$��ZOV:�]�����c��i��{;tk�H���m����&�+��gC>]w�4ٍ�P�Z�
�h��[8�c�����l�:�bа�6��ZzR��X�2��*~U�n$Sb�����rF��Az��E?�0����1d�͌?�G���^ �Q!����Pv,bj����:_� �W�͕�M�� D���$b����ї�f�8�!����T�>z�W���k�_�Ë�4^�è�T�}��Q;�!���<���u�)��=	�L��h+��� #@ܿ�����"���`Oud����"<j��8�e�hoieC�H��'��(�A=����/n�@��Ts�j\#��(P4X�pZ�qn�7���$��G�t���MTF@N�7�`U}�o��H)r�\�V���`�q������'D5��ͭ��%��o�V�@�ݸ����w*�H@��q��̈ 5D9�`��
��fK�;/>�ߋ��v��!�ё���hG{k�Ũ��=�dY��S"�њ�CX��T�������Ei/l~�����֤!��Z�e�hjlAo�L/]�{�n�9��Ir�:
��s��Cs[;^:�{�6��<��� >t?XuNNEb�鍌9	��pI$(���===�?!oC��;9.�ER�W��E�6�ߨYL*��ᾣ8r�
�"�,Y��"tn�����Ʀ����a.�۳�#�������840_K@Od�/D@jp��r�ip��)��%�P�(u9��_���!.�:��#������ڨ���{2����A�)������wQCZ��BR�4i�e�TH�J�BiN��&�JQ�j�iFm�����""l����}VI�06�=3���sx��qpxN��s�4�Q(��b�J$��7�R�o�����)�:ĤpZ¦�,(����m�z�Y���{7�v�k����@qah丂J!���#�a�>4oh~{�w.Z��+O9e���d�'_���O~�bf�/�Z��$ǡ��2_zeh^�XgC���X����x��o՘�x�C�6<��?��5y�eKy���k�Xcϑ)V���F�j�#O+z�X}$t��Й�"}Mh��b,֦|���E�:@y��*Ι���A�҇�p��2HX)n�⑑�ST[��E2��W�.ִly�Y�v�@�E�߾�{�1�L,_<����1L�,px��}}Eܷ�9���##тj�`�TB���
hmk�'-춎��1sO;�ݷU#��L�܋��w���X۠g�(+��	�����$RIzb����6��i����A��~ z�j�A�*�G����Lu��5#�ej{Է��!為h��O�
$cG���y|��ƹ��9n:���8i?��#mOe[��X��_&��&{�'���[Y|��X���qǆ./��e#~�U�L�Ο��T�T�j�r�jlzl����Qƒ%��I�~��1��Yjj(�H� �J��]xU�
V._�MR�I(G� 0%a�tQ[Sc����	��]��+���Ӽ����x����	e#"JX�tf͙�߿��K�ԅ��Fz�G�4���9j���e0&P%p&������ʿ�H�#4~�p�.� 3f���nܸ������6�9`E99�ǠN�fϞ*Sz���ػw?����N�L��Ck*3Y�F/^�\.��{�ؓO`��[�k��l@��yVGF
�S9�*�A�&�n��֤����9�A��'��D]�Na���2�7�ho�1HE�&;�R.����_��zD�ڿR4mp�"e5!Rv��?r��)eB���������	�5֞B;�〮��ͭ ,�1t�7H"���#���F��G�y�s�65qʐ�*#�27�JJ���`L�(ĕ 4�̂�҆ʀ�����}�E��sO^V�f��gw?����_��H�]%�s	v�J|�İzȩ�Ђ���/[��e3g�!O���G^���'�����]S�t�(��2�.8���K�-��s�ek.���3f�C�ǿ�g�C7b���'��5�$T�[�G���ᧀљ� �t�R--=;�vE�K�9��Ƶ��(�&̐�=�QH��7&nP$@�7(r���By fy���W�?bd;gV`��T�.t#��ᥗ���g&��F�L�ރ��V(*E�U�9�����<k.\���C�1��B�`��!<���xu��B��l��##jBK�����6w�k�,9�<�|�è�)�Q36t�G��~0������hU�N#�I!�6 B����б2�r�vM�m(U}��BՈZXRbʝ�O=#�t�Gs\�����u��@�Z(xŭ�a1w���	�uڇ���/���\��&���=�x�'�\�W��N�o�L����d�;��ֿ�<�8quȺaI�r*��W�Lc\���&G��ꝝ\��%��s���E��SıC{���{�74d��э͛7��u��<�-�i�dr��H�l���^��s}Æصs'S�<�Hi,|�ZH�[��,>�w�Z��M��~	d����7&"Z��+��ܹs9:��j;w�`j�0M��)�������oꚮ㡇¡�Q*��;��CR4�ѓ��3��N=u!��w��l~�>:rS�uj�I����~��r
7����b;��4p���J�̐ք���	��x��ʶ]�9T��p�$�n�FE�p�i5LV�Ǭ��2|��%�4ş'�5�ߎ�ZDu��Ԛ\"�ǘE�� ��ȕ;����Or��v���-�6PM7� ���8ym$�e{˔<�S�`Z��^Փ�G�őAM�&���U+Q����WCp
p���E�Bs������X������E����ݬ��f]d#��B~��dC�*.��PO�0���ՐU�Ց�����>t�]o���DI�{��]�����J�>_M4C���(U`����T�N�n����gްlf��O�2���n�����`���WEF�T�dƴЁ�
�ͿޚM<��3�r����=z�샛7wo~n��g^���TcǅU%5�h��I�I*��ЙN�k.��s��\ u�^�M�R���0�M�'�q@��i�;"Q�-�;|O�4	QD��X=.�DCH�2�P��Qs�>46d���SO?���!�j@�⠩�	����d�8��� ��65�36�Lu|�'�n�QM�90�}��p�Oa��AJNH}��T'ݒ�6��v*�!���Ђi�`���ֻףzp�������%0��Ǝ�JI2��h�d:%.k�:NG3�A����F��r�{r�"~�@�f��L�����T�\8	C�ι��H�S�����K<�9�>�.����D�~�H)���o��>���Ll0���le�A�>��;�輞o�6�����O��zLH���t9�ki��s�=�|B/j��#�*0I�[�#�o_s���0�������ɏ_�ŧ-��}�{��m�܊l*�S��Ē�hz��5�\����~��,�c���oKjq;�ı�xA�Ӗ.�(���Gƍ7ވl:�F�Ɩj�i�P7��?�O0�=28�{�۷o��<.E�t�l�5��O�S\�V�T��oȇOɧڒ�MX8x`3����s�=�������x�)ޞ�BjΔ`��?4�w��J��W��Y���^Ǐ�f�mC6qʤ�|n�r�袋���hj����]���}���W��5s�jCU��IP��惜���1(����l�9P�'�Mf#G����`�娫�f�H$<Q�.����ǁ:���FmR̔�?����e�5�v{w�g�~Nz�=!���`@��XGqt@G��SA�( ��K�J	!B!��v�����yߓ�s}����I9g�w?�]ֺֽ���b�A#��C��ƀщ���6P~F�nS�l�#aW�j�1\RcQe�W��g���rUP�"L�Lբ4+�^I�$V��Ŷ����T�j^ �@@}V�VU&�-]���{![���/��>]��<�*�<��\��m~�o\�M��u����q�`���[뾴c��OM��p+R�*�N���Z53�*<�\d\{��K�ϸ�s%��7l�f�ֻJv��D����D�*����Ys>S)��V�f�Y�w����p�)��=��>OGw�Ю���b�<�j��,�V_��R��LMU���ć�� �!��	"��UJ�5)������:�>g%�R�(�`��.Mf
��ߋk�ɂR�.78	EV
0�"pU����^İ�z�C~$z;�r�?\׈-�nA,�5 ����VS^����YC6�����#{JU���@o��ǟ_�O�u��
�W�(�(te@�a3��fG�ȑ6a�����zx�m(q�ͥ2�-�ēȤ��Ȳmli��_�|.�ة�8�v�j����<��4IT���@g�.�C�3݄�M%n�<�$>�j�U�Q*��ֆf\6e "0Ϗ͝�%&���ӷ�L���I�3�]�O_� r�?�w���4Զ>�F��`EA��J�L �9+aY�q:�~�����Rlp�yN���Y��0��XRՉN&c�"�@���s�c/� ����%ȑ�ΥV��T��f��R�7����݀}�~�j)#	��b��EȦ�x���g�>1����R'��c�].Y��o��$�w��(�UXHz��
�_#��h,%�������#��[����ϯ���&��Sn�{Ȥ�{���X`Qv��*�B�7��떳"L{�M6�y���зlۊ[o�U��.8����(۳k���=���}7��ήn�����v�鲰�g�B ���g��_\~)b�^X���w����O7sΟ��C�x�&w�ꫯ�wo�A�h�yi��~�\Q��hrbؘ)8�ы����C	V��*D@G�:u����IH佥����(1y� ����UW�ӹ����@&����W�1.���sˤZ)���"Lm<�iP%/��ht缋r�e����(�[��iE�My�눒�����wB���I���	�J�b.!�ՠ�u�����Ջx���A���Ī�u�) �#�������j�l�xR�'*�MM�kl@4�P���A�3v�7�ȡ��D�\@�L��8��)�bЌZ�$+�]�*̅$|�¦�̾��sgm������a��!O���?wF2��y�L-N��j�Fhu�`3U�[�o��ٳ��������ؽ����	�^VI�%�ZM9n++	C�R.ej�B�V)'-�J�f�^��K�8v��osy�e�f�̜[ɬ�Me��O�
j�S�J�: #�I��egV=�ɮ�V�ޮC�<���e��n���J����i� �F�P_X���� �?x-5��:�X�	�{�<,�?{v~�\��x!�-S�"ErX��WC0`�C+a��x<f��8�L����V�7r�
�8��]�y�}Df4��EIXд�U�	�6;lf2�lZ�4�;g)���o`v�e~^*�c���%����E��Z��&a.P#�����C���O�dε�j;���m^����ga6���p��E����y�8}5:ڙ-���ҥ���7)oh��	���w���w#��멺L���BW��5���R����nd�W^7F��1���y�ube7�u�D-��g�pGy�3D(q�ɟ:��b�b�S0�*X-����9繭�[�[	��AƢ�r.k��f�?��-x��pp�'4�B!�ŢE�ce`{�����#���d\^/ �r��x�_|���N޲�=���*��8��.;������R!�1c������&?r\V wuu���A%fX�2fa��_����-[���n{W~� ̪
".����믗��P��?.?����fA�\�n���f���۴�����5�::����P�}|$��2&�"�O�?�8l\���ඟ�!K\�9��$a�]%"�bA^׿��X�x
���.ٶ�pP�Y�(j��_@Go��eT�pd%�r���T!��(8�%G^t�SšZLdl)7,W�Z�DY&WnV��˦��8�<&�<��, t���̳���n%��0�
���Ha�s�eX���׫�i�'[\v��Ț��JaB���7>۪��bL��2���X��E��ل����.ŀ�,��v�4Y`)��Kb�);Xd��fOO��w��x�~��^7�����X���L(*b��b*�M�b'q����ŮJ�b�!���ۥ��U5�J��kh�����_���F��o��������ښ��ع�6�;4�fv�3�<�~���2C�f��T�_3�o����|����Ǿ���?V���|�.	]g\	� �>r�Y�H��,ʥ�$5�X���|�<d���ӡQ ��?TZfHx��� �r	~��<H��g�)c��*eU�.�e�ftS���UT�pH0�Pz�9�BL�2�<49&t3�ݧ��t�>�F]Ѝ��F���]�������`�J�D&��x4h�"*�B!<N3�.ZZ�{��)6�5��Ďw�![0�Tg����$�
J$�Y���jlmhliF�b�ɮ^�����;X��]0	NND����֢�ܨ����J���Q���s���a��L\�T�_���_��g	���F�9����lIvq�$�\��m�]�G���C��Gf���f��ϑ)�C��*��u���"���5� �稾�}�����M�G��\dm�°�BQߵ~�\�`�*��tM�oͤkS3A&�t)Y���1H�sc!���)�|�P�HХm��}ɐ������I�?nl�hL�"̕~tӍX��oس{'�[����$qs{����j�� i6	k��=
K��,��h� 7l؀��m(��fU�YaA����6�����|�3����.���@Y���s���j|�k_����e?�я�l��&&p&�;��~��2ƺ��{�w�����StЄ�E�W�e�.��~�3����܅�n�I�r��'y�����e�]x��7�)�ا{v��w�'O�B6S�R*�.�NJD�z䑇��y���W�q6n��ۏX:�	Sg�/]�?��0z"I��22cq�W�uʎ���?�-����;��Y>#oS�����Yq#�F��������܈��ȕ�����5тBQ�\;��pHB7�]&t,��#3�J���}�a�A:o�5���T
��_8����
t?��M?c���#3�3�5e�����Q@"k�a!Z�\D9m��l*�T,�\&�7��_�B�tJL�8Za1�0�5��bD<�����9�s0Y�:PFcj��"	*c,΄m���l&Ѣ#/⽟�jox���s^8��������h���+o�۲�ӛ��.p�B��)�3�Iv�%��b �췙z�6~鼉~.R���?��[��[v��N�Z>W�"GT3j-?�Mt�)Kg��ĊV�Yd��)��Q�Yf �n�
�Շp��č�Ř	YM��T��{ơ�"�aJ0V���dg�J�U<u�.�2��w�!�3$��X��Gy��d�D�L�tJ��nE&��fF��G�@H�,�Xq��{,Ҽ�q��r��U�\�1e�,�JKB.�.����&�\���p�T������C*XJ�ʵ��dY)�IJ�xnTs8��q��.�k�m�6�2\:|e�{�x����M���f�#jX.��IL�f���L<�
=��K�����Kȃ`�RGZ��ݦ���yJ�x�dn�u᠘xpcW����$cј��^բ���/.Vgdi?K4:vvO� 'T�3�a�2�DV��	�)����D.�߾+I�tszqȳ*��jU \�<�݆�r�B$ɰ�Uݠ�-�j�ىH��3(-4K�O2�b1���Z�ږݕU_2��O�XE����� E�P�����-E}((c���9��B�\F�\&��7�:&N��)��o&j���U'Lș�1��$A9v	���]jI����I����S��TƉ#��L�?7K�Ё��띝�%���QI����H�|�˘>e�<�+VH���$EcI���qhVY\t�2\��q�*��R!BwEnD�M�ϛn���G������x{�fٳ���d"�ӡ�=+䲂^��]�ɓ'q���[�iHfX|�2�;w��7��CR\��b����Ĉˇ8�ҡu�{ԹP����ι:��3�eR�G�Z[���xEr�Ac�y�	K!ANzɗ赡��N� vf/������{WE,�`��a�e�L9���y����7#�ϻ�s��0[��	���̐�d��    IDAT�x��� ��
�~��~�%����%a⹦
��ɢ�J!��+p��aÄ��'d\C����	&��:Y�"z)���D�|�"��XS���/�7�f�@�2��QJG��X���pp�̩S^?{���1��	�II�H�;��Б�ol�<gߑ��k&�<���.���hA]}X�'�&G)��L��Q�u��x���>WB|ö	���zE��M��B�� wY��Z��fق%ZJ��1d� @0a�uCJ7�|E
��(�>h9�e�}�g:�3qY��_�d�)�τnF�T�K�)-$7Nћ�Ŧ>S�$��$5�M�%8� w8�y�8rɘt�C>$S144���X�c'�!�IʥK�2�q�J�����*�;t������U9����0j(��Y-�a��E"&��V&"}���!U��r5XnT�6�=�%3�o��%�ŦCC4���7X��v�O�;5���"�Ǣ�AG-E�ʶ2xcV̟�����`s��Fp��!4}hE2���l3��f�t.+sA��9CeWa��F H�D��	��:iX�nq:�g�V�8[	gbO�ad������&�?�uTB��g~�U��s�unB�3�����X�?#V�vMf��t	�T���r:B�Bd1��|�j������[*á9�ֺ�r�{T*�ē�3�°�Kd��ul�$ౄ6:c�_j�����ט�Y3��g��-f$q��u��?�91g�R��25�:�����e.��玝���|N^�����fΜ�P�N�-4i���a�r֬�kNA�),Z�]p>NMwkּ�����+�&W��I�˯�Z6����?��G��Ȇ�,=9��MoE�0w�Y�1q��Ilٹv_ �@@lomN�<�w�ۢ�+�U�%�b���J��-z�� �y��,g&z2S!�L�7��:K�|}}���3�P�A��K9��͢��Ӣ�gm�4y��נ g�/ce+��3\��N�Ю�f�r��97SIc����X�D��P��jD�:����ſ��B-�NL���Z��<�)�?Sr�(fԽ�ze��5UP���qi�B�\�L�]��=��0��d,�l� �ǃ@C�8br	����e�d�U>�Fq��6eG����\
~�͌B2V�Lծt,��kw���nm�q����h����wj"�U�k�f[[�ls�����$�B3'.A�.5�0����ϲ��\:��~��I�׿���杓(���BY1$t�$���K��ʩ�3	���dT��|Ht���/��3^�ҙ譗���>Y�E��I9���̐��lvs�$�
�6<��)�%e<!d~��yP)��t_W��H�b��:і�fD�}ȕr���2�#���.�����U�,�T�ve	$&�SU�������B��219�ֶj���)��
��;�3i��NI�@b�i�!���/�X�瑔ڰK����H|��N�3��G��FY7��� MB�~�)A�g$���Y,�q�)~�^��;��4	�'�E���e�bPK��v0��Gck��}����A4}v'Y�J��?v�dE_w)�� D�T���;%{�;��>�-k,��b��u~�u����_ê`A"0���a��ՙ�s�4��I	P"��D��l�o���j8����G�8ggd�.J�&�E��Й�y�U��\Mf�u�4�TḤ��_�Kuk(S�[)A��D��\6A�d�M.'��gK$=V�M�r�[NΓ$Ji�B�+���A)�����q���	��*�fH�&�!ÆJ���?�^�b�֦>Y�&�����=�w��޽[�/��Y��rv�W�������������w7�	���y���|��a�����
X��߰e���S kei�d'q�Ϸ�[n��\��_?��lx��v�v�K�/�uܣ�n�h��Ĺ��4J!݄1Ѥ���2$&|�����;��u�2�9�T�9j��Λ-�(�����=>�B~T�V�(i�Vp�^E��i_%��P�kr2��z'Ji�~��pb�"Y�g�ZA�p��,Ks�B��+!�v6q*�(�6=]HB��eY
U��z�%w�\�b�Q�[�7��L�ׯH�e+[I�[%h�*��<(���U"�w����f8\N�:qZ΢��9!��9�>+�Qb�3�|!D����sv>��,�����$耝�B��J�R�f�\�R��,����VO�w�V�j� jf�7��ɳRrV2u;r�L9��V������7�?�a�W���`U�΢}ᙄ���L�4=� Cw.����nїAJej@��y���I.���Vۤo�Rd�~R����c�7�y�%�' #��j�S+�U��iG��V��Z�\�u����Rଌ�Ó8q���\� aq��@P��wv9p���B.�G>}�1=Pӻ�(.k���E'�j���rM$LESl�x@�Yv�&�57\�R6��Y9*KT�y=v��)(CM�'DGw�\NXPj}�"f�[��sxܢk�K[����W	WUK4ڈ!˽�t��%M���v�t�<�DX��9e(e��4��������h�����iX��:X�-�JY�n����H�g6�c!E��Й�H`Qi�݃	�*�]�W�,.�lXPI؎�Am��
	)��=�3�9��0sp�&p3��|eZ�֐�E���>!\q�#�
 Pr}��<����&����xP$��ͣV�&	0\���ɕ@��A�M��%i���'G*n��e�8� ��^�E� u���U��x蕏 ��R���K�2pZN��B6'�_D��j�+y���e�A_n���%�p{\�=�й>U�4at������A�7)�m�y��L�A�򃧩�fs�I�f�pqK�*c�aÆbܸq���p;��ߣF�<�B�9y��s������on��W�`Ǯ]rƅ��,�kTL��+���ӧ��[��+�蓃�ٹ<j��$�]
��Y��ֿ������������.��$B>{�j̒:'^:z��T��ds!���Y$����!Ţ&���T��X @�~��Ȧ%�a1Ɵg� TB�S�$f����k���~U܉�S�(����0gB=��;hr���C,�����ϒ[ 	7�����߫VaR�ĭ�)��)>�U _���ml�:v{�hnn��Bn	@�T��6���66Ib;�3�ŕR��
���4G)�*j"e$S^T)�S`%T�#�JY�$��2��D�v��ETLuj���"�l���&�\	�s%����7~P�w|��c�?�����ЧL�G�N?�ȗ�|�U��*x�$��{�J������8ah�uM�?�6X�,��^�_���.[��7����L4|� \v�E��8��Ja'�Rʡ\ʠ�),��z.�����r�K�<2)���A�����������Sx�����a�	�٪�,yI���kr�2c'��$�F��pp�R@��u^]w� ��ԬҌ�CA_.��	ϓXR�f(�
�#���E��Q��uQ8�a�@�29#�$��m�}���h�aE[}A��ZYUȜ��E�gȺ?x����-3����=h0<N���L�$����f2����m!�5����
0��k��Y.�n,�KZ��
B!8O(r����"n�@�z��Ku�g<���kLq��ᕠ)rȚ@�żZ�nS�i*�Z����	;?S��20�ǒȈ$�2���P���N�lH�r>Xx���g/�������<R�_���g�˔[��[��Ƣ��B![�s�y4���S��Ύ���~>�EM��t��ZD!i,��H�T�o�U�`H�b7&�F�[lfaƓHĢ�����fe��7�	t^����\&-�Q �;)|4Ս˯�l�"ɗE� d��:�	�v�ۣ6R���HIm��f�f�IƢ��"�L���AF
v֚u��Y�:�=x }���rޫU�	�$_�U��ѣe��r9���a����)w�w�c)���
��e<�k�U����)��qH�pM:]AE<n�OL�F�9`��طi(ռ��|B�s�\��ht��@$ǐ�av�9��y�n��[Aĉ%㜑����ExV|N}�CH�6��l4$.�8D.�9wb�ϸz��O����V����VM��.>9ƨ¸�|J�ο��E�8U6�%1>�7;�#�X�[ ���N�u;z�,��ݲ�(U,C�ln�3'c�$Jz0�._� �9�KY���X���K"�D�J��'UF6�Q�X��0�.�����Τx]�n�HBh������.�7��5C`��9�o�����Ȅ��r	F�Yd0=S,�C�OH�Y��E|s<��/�3I��BI�/V�R��ŉ�=�����%ܳ�ѓ;SV���S�b�A��A��.Y�L�矍9���?��tg�5�H/���Xr�8}N�R��Ί�x*G1K	VǏ�@<���^�
L�1;����y����_C_<���nؘ�X��,B�ʑ|�9_Ռ�?�L4.2�	t�*2���8�"|G�/��a"�tLLX�ȳ���
[ɢ�X*��9;Y&}aiqH�H&(dR雄EM��B|��т	�x?��z4��9~�BA��XR=/U]}9���BfW$�]p��56���Y�I*ET��â�w��xm�6<�j�>�t$�SE�i	��L������N`\s�B�����]>��|��8U��Q:mr8���0�T�dīذe>oz��T��"+�\����>f�	ٙE#Dm�v.�P��64���1�q��_�"�h��L��A���l8t��z�i>r��0.��rL�6MX��`ԇC����t`�:����x��pz}�?M�o�m��0Lv
r���#�\<	����du�٬<��T��>�4,D�u���KQY��-������+tH/������i;��)=�d7�!�hj[�Uى�5l(|^�3@�����"���h2�e7�v���]�]nA|xn)�c�a�j��BO4�H,����2Y����M�T�L��7n���b�lA6������Z-�
ʈKPO.�tJ,8���u�r��5)%�,,��ۦ\�ؙ���&�!�����C��N�S_l����B��n��H.M�p��1��45�RAe�*r\@� �-g�gẗQ��=:z�q��q���ğ��n�^��z/SJV�͏D�{/�Ro.�DZ5I��Ig��1��Uf)_L���M�u�l
8��<es�^�X,��v��vt�(� F�D�8Ƒ&�dd}Lf1#_)��r�D�x.�B&)�+��<;.%��XE������bp�<�0f4�ɘ,y9��-J��+H'!�T����L�!QWx�>$Rqx<>�eNoTy�[`pX�
A�����ώ��<'Z�q�B�[M��J�|��ED����;���/Ο�����cz���/�,����Vo��Ʀ��38>U��P�}i$��[3�ˆ���W�	v-�L� �$)K�f��l�Q��C��\�ǹ	��7�؀r����7���ӫ'U��%�Z��8o�,�;���(g���_�)�wc̤Q�ԊB�	�� D��eQ+���#���m�.܄��'�oj�������ĳ�#�*!���QM:��٬�t���p����v�\ұ��<^�d˄Ҕ�3	V�,.V;�cvM��urNX��߯*B�a��Y�N���)2���+�I�'T/�'��m.ň�3�"L�n��_�y�y�>\�t)&�/�t�� B�cw����;ҋI�'`��H��=s��$|�a:q
=1� vѸ'<����r���"�� �d�ĶZ��E�1�j���. ��<�
))���s�p��C�,	V�P�\����e��Tũ17���	��j�:G�+5��Y`�\��|\�`!�x���{Ɣ��<yB�=-R?ݻ���դ�gφ��A�P��˛�A�*w]=��<���o@o,�L�nh.)r���.����hN��D1��qnB��4a_. !��c�"ύh�p�0��z��tC�e���aa+E��9K�5�#� �J���Y)9��(�n:���2��46��� ��.�c��9G "Ƣ�2K2�w��X�iٱ_�lfL�)��4mvyM��ڇ�^׌O����Y��sHg����H���IQ͎�]e�zwJ�"\2�s�[�8�{��s�z@D��xvK�'�JI
&n��n�=t�8l��M�K6@TFE�������Qݟ���fCS,�oÌ�1u���u�tw�O�>�M�f,�šc�xg�Θ0j�,<�,�.db1�9��{�9@��[]>=v[��/T'a�)���^��P t��d�8Z��,#$���3 �X�B�����(�B9r*�R�} W�svv�2�q��$7B���sq��I��4�됻�w��-�\>��R^��H9I4�x]r�x�Ydi�|n:�z0dP�C^)\��b�z�	X���N�SY4���Gd�c	!�
	���EQ;�QU��ץƝe9s���r��>9v�Ѕ�"�O���˦$r�&2s��R@�a��k����������w��eǟjZ`lZO�$[I/�w�g&��)���~�6u�u��rټ�Ej����ʋƤ/��@�,�3�e��YEQuFR�9�Б,��`��],,Y�-L��e�-��/��Ϫ֯~�
\p�98x`7B>��K�F���d�B���T]��N?�\��gP�s/�BW,��g�Ť����u芦q�y����,{k_X����]�D\��:,E���-�êu���8q��`+zx�Aa.g+"i0k$�@�d����h�tN�	�9^6�x��(HW��<Ov���4��#��xAY J5IȪVF>����SD�O�����ŗ��cǎAO_��<�A?��9/��O�xW�L���p��)%�z|:������(��F�[���=x���g
R{�N�`�J��^ݼ���X���'~D�)DxY�^�T` ���p%����Y��������G�J"2:�alt�Z���C�*�I�u��3�̐�>,��|Ś5�ſ}�L9�]sfN�����'�2�S�`6#]����Ǟx\f��&���T<��">�TU�3^T ��9�	��f�z�(T ���^~�L�y�RI؜j��ʿ��C��H�qs,$��I�����1et,�xC��p��L*��.�)ϛd-v�t�}	] Q}�P!����'��)Oub�E0~�G�����뾎{��=N�:�I�#����C����g����$9���{�C��ȯ͜9��@o�W �'�}At�5�&,�x,!�\�z�p���Q��UHp�hٌ$y�㒐ƄM���Sݮ�w��B��lm+�Ld'(V6�+2���i�-���<g<�D2���_��[�.�V���<���~�ƺ �����������X#[.��/
4}��p�up�lVP\�H&�T���c&�mD;:����q�n�(�Ш�fA2��g�ED�q��yOD�r\�C�V>/}�)�\�E�����UB'
������-���<���,�{i�ZQ��E�k�����VW	'�>�n!W�k��	�Cpᢅ0�rp�-�KDP�)�"Q��˂\���%Y����p���a��	�Fz��[�Ԍd6���(��24w ����壝�
��I3D.Hw/ϵ�qǨ,�(�%�'&ABX�!{���yH���8R��n��������46"�C�JA�����9oф{綷G�?w���ڸd��([=�9��>t!��	�/T�����"Ro�JF�פ����&�i3��͠�N����8$�Z�E�	B&1*i�U(�QZ׌@����3�A�(�V��u��X,;�E�����?ߏֆ0���/b������h���tWO�Vu<�$K�N�l۲C����_^�T�]�1o1���3��7�߼Ͽ��!/F�N	��k�����`��)����.���2�\��}	d*NtF���Qbǉ
�ȣ\��j#�B1_-%
��ټJ����(�A9/�<W���0�P�}毫��ϋ��BJU�>1�`B��t�J��7݀�SG��啘<~�u����    IDAT
>r��dr92YY
�"+	��3c�Ǐ1��a�ۛ�k�a7	��6l�s /���'�/]v%�Nl�:N��ϖA��nǚ7�tM�D
k����5�yX�Xm�d��Zb����YV� B@���	�RI�R)x=.A{XȈ��1�	���J(WA���jq��Ht�w�����){$��0H��z�^�e��W�ݎ�׋�\{-&�+���i5+��:���+]:����sjmG��O:.��%�~':�p���BZ0�o�|3�ǨQc��sϧ����9kچ��vb��I�]2�tZ�t
�־�L2!�
����@K'A���jQ�"���(c�LtG솫,�u�_��Dֳ�J�BW*��toz�� *c�2�N�2!�<e�8��7��o�M��K.��l֯��i3�������U�O�p�	��ύ��9mj���r����`Ҝ�x��j�f�p{��=�Q�I��p+5��G�!�o���p�"��� �e�DV
w"��}GԲ��9Wc"���Y�e��#���֭Z���FF*$s�`���BĄ_��mx�Ux������eҘPU��un����Å�_]�=�`����oA��B�c�`�Rn<�l	p�p"����lƩ�(<��
}�u�DK��y��A�R�A����+	�F��CM4R���H+�J�:�010�*2Z#�S���[�y�At���`�k�d|!E�[
�|����pɒs1c�X���c"ښ+�H%d�.��X�����=�4����?��G��j�1㧢}�(D�EĲ%��nb9*{4D�1Aq������b����= 1���"������9:��n��Z-�:�az[̄�j$􀽖�Vw�9'�;��@�w��e��ﻯhqcBϋFI�&�fR����rU�
�Tw9�B���|V�J�m3#��"텕�K��'s3Vw4*��<[�]]�{��,e��`L���ofq�I�Eu���"0i1���sb��I�����r��?�Y$�>ف�ӧ	C��	��x�*�F"xػ{?Z��P�b���/����ƌy���o���#���/��"�s�����Ǽy��bs�ǻ0b�(Y+y��~|���+�_FGoUG��.�γ����8�~�}]�(繀Q��	A�O*vv�	&f^�j'�U1�1��B"�	�<;K7�e�'��K�*)��\>��Q���?�����O��]y*�N9,�!&���z�g �����S�p�E'W������f�z�q�08���ឃx��8{�9��W.����nxf�=�؃\�w�l�sv�����ӋW^[��~��z}�m|�@ E&���d����L���V.���"�I�L4�Iy�G䉆�[��(J�ґ�_4��9�p�������$+�ϙ��#Z>�k�^��c����ݍ�p�_�O�܌M�6�� 
Lǹ�Xyrv�3�	�Ǣ}9l��c�ۺ�p#���"C�ß¡��p�����6w��7���Yg�����{	�<T��D6���ttvJ���cCYBB%?3�b!�j)�݂X<�B����fs��9)U�W�%���(����J=-��g$��,�3��\Ȧ���1���wq�o�C�c������.�A4ƥ/�"�E��.1B���9f�����6qj�)ȓO>���CP��_ ?�$��̓1m�m�!xi��8k�L��4����>��׋��m*�Hc�{�!�� ?�&��:e�#GE���S�6�݄��J�iH����gI�kH3V=+3�~-���l����Z8t�l��;nÖM���a�Q���!n�X���ijh@WO���a�<����V�����j2/�y�P�,N?���ƣ/�BӐa6dh�
����8q�$��S�2�da4l�h�lv�ڻ�ty��.���,Xg�\$��\�Jj�;���=�����Jm��i��]�j0��/AǄ�eH��/i%��O*��p#Fj�o��Xj|���0hp�t��{$��vݛoa�;����ꫯFKCX^g�D:�ģ';e�%��5�k6��d��$ѫZ�u4<*���S��,.E[�ʸ�����t�S�A%q�(B(7��j��6I���I��W�UJ�)s�x�T
�ˉ���ߟ�`�}�+��~�_x����`�/�����O���WJ���E�(�-���r1.���j���@k��7M��:C�J���8��+m�Z	I�lS���c�!�/�U����W�KX�t	�������an��71i��ݽ[�h��J�2��ۍ�A����%pc]X$:=�=8�ܥ�5ࡿ>��X�ˍ�/Y�??��&32�8.XzZ����Jq���1|�2T�'N���[?���.���l��c'`r�![&��!� �<�4��j��t�E ɢ��i,��Hw
��@Ʊ�Թ[��
	�)���^�K$5����%0��p�"����
��V�ӵ�|G���s�Lŵ_�
ɾ^?tƍG��Ȃz1�'L%���&���aР!�<n$���S ���1l�d|z�V��&ڇ�ƹ�'��:��T���̖]E�jlnA:W�K������ol|��nG�lE��D�Û	v�K <5T+�%��h��t�u!�)v7Y��.jΩs��@�J�a���Ը�:	P����Kl��5�p�e��\�����}6���3i|��#44�j����P*��3��H�(7ߥ�2e��>ݍ�6	��
n}�)q��K�/b]����v�e3Y|�w7��1\�������_���H��t�"ƳM����^
�%�֊X�����r��)�G�6)ȥ����Lr�ܫ��ĳ�|T�^�n��sK_�����<a,�Ϟ��V>�l2-H���«��$>��&��N�0)��6��6��`'N�B8� ��_|��B�--X��{غ�S�w�rL�1?�0Ξs̵
ϟ�'�+�ٗcѹ�����J�n��V��$�w�S�-	��k�Fwzh�T'�,��9Sg,�dR��j�e�*��
�`<�B��K����D�A�Id�#�˩Y�\�-7߈�ﾍ�V���Q#q��bX[�p4���8�lFg$"z�t.��jn�TL�1[�}�X<�RMCc�Hl�� ^z����Cڰh�<|��^��/�7k׮ż�s�c���8Y�SA���GX�y��6kt1,pi��֐(A/(7�0�*bÚ�'�yR�ϸ�$�����/�@�`��r�Vv�F�>�1O%��,$�'���_CKc��d}����aڤ�Ȥ�B�en�<.<��38t���r���rL�8�&��V�7֭�O��E�/��Y �&NĐ!C��[o"�v���E�K���N�>]Ү�n��x'�u��q�@"�&���U]vK4Q��'�R7�z��|&���.	ݯ���Bw/]8��u�q�%��:��l�6�HM���MUUi��%��9��*��Y�J�&Vlze���P�gQ�3���1C�`����e����N�q�K6�/�z�8	�Q���4�9��^Ew_�`�kW�"=`�Wҗ����k0���ӽ"����Kq��ix�7O��"�����o��Dv	߼�:�>ў^twtc���?i*�����L�����y\���E��p�VD�z0o�:B
�>؆��VL�2E���+_@��C�ǒϭb�F0ٮ��PɊ�&	p�Y�4�����<.L�"e_���E!8Qv&�d������nZ�ڤ�K�\΅K���d�pˏ�/	i�ߞ��Y�p�����i��"�O�O�M&��z}�v�څ@(�Qc��?�P��1o�9ر{?V�ۀ@C#��xх�G:1��;w�����Yg�þ����z�:\����������6��f���R\��C�r!�l�;�U�Q��o*�#b<�Y��*,$R�*�e��+ZT(m��`��.lzs߹�mk���+L;W_�^M~�f����A�g8�fP��bhkn�s;N�<)��̙��s�.��u;&̘��\�j�<�4lN���5�0j��z�}�)y/������o{�	�>���"����P�XK�����i��]��+x]v$c=���p{Of:t2Y��(.����Z'��W�.f[��%�2�f�袈�b<D�����sf��'��b	7|�ZL܆��	ǣ�����H4*񠳻Ç�����1t�Hqv[�j�8��D�4c�~�/�x��8�/�G���ݏQCa�ԉ�Էmۊ=�����>���vL��O>�����f\l�H�bC"F<��k���[F4-tYq��)%��G֬v%Y*S�������=`_��r�;�R:DVē�e��o_'	��gެX�h
���'�֖����{}ș+�{4�qDz�d)c�I��{�A�������{��{�I�q���.��=�&N���`��^-���,�U�+_}M$��jٲJ���W�c)��I���.!�1����K̢~]P
�6I2ӓ�@͆�,	���E(9���	�;�ǫp��!��o�=�R"����'�5y">޶E�qBM�eS�W�+�7_u] �b<����9|�m'���X��f<��3��9{�B����c,;w	���D���?Q��X-��˯H��1����V9"�*����,\ҍjd#��j'��{g��8Ǳ_B�������\���=������c�fkgB�p٬C��ɺ��f�B��C܅�?�Sg !D��� �V�cD{.��|��x��#W��6^_�=}Q�]�J��������h�!��-{���'n�W�����$���6c� ��c���0c���ǻ����U�����X��Z����0f�Y����
������];v�QG<�����KfM&�C���\<���K���{P�f�L��6K�m]�,� ��Lg`w���{�=�ٿN�C�Ƽ��笝�#���s	$�O�.�E>��ٳ�aƌYؽk76n�(]v}c�����l��a�Zu泱���g:�r�$�2�Gm�&�Joz�����+��ډ'�xK�����c��M�0ffϞ��Gذ��S}1��6_�����"�[���(�,���_�����k7�4�/]�ǃ���{W +�(p������K��R͌|��gW��#�N�ʹ�ݎ<�e6MԨ�(��t��&R���t94��wP
���"�[ ?�e8�6�,5AUH6�f�[�2:�&�R��P�p�V¿��6�7�;7|(����ɣ�@����^��g���O*�>ݵm-�b��c�n��T���fã�=�D:��}��0u�4���;�=�����{���!Trd����*$�Q&������2*$�U�r��ݟ�ZA�a+�B:�xO�b�Ө�_��/�I�d�	�tݺA�U!��8�<I=j��C�G�ѥ�4�L�r�'O��?�����s�����¥0��b�B��:�HȎ�#G�J�N����Oa��i�y��=V��Ł�on��ݘ4c�9o)�y���4˼9���I,_�\>g�/�UkV���`޹����t	�AKF9'�Z�&�M�[�,(\,��K+Y�7��K"��J�J�8�B���.Y��s|�g1J��/�"�I40��r�p��n��7_ú�����c�Eh	����w���tL\�a��/�D"��p�T@wg�$��[?��ՃRɆp�Plٹ/mx_��5�	O��_�(�C�eRGt�����i��_���Z��ǟF��1���rM)=.�l�7s+�\�X6�I`|�=H8�]$��j�J��KNuR��i�vI�(5>���%	��9*��`.��xs�*8MU|��+0�!�]nC0��7��u�/2iCs��Y�M�0y��!̜<�D	۶~��c'�+��)P��>ľ�1d�p<[6o�5W])�`��'������/��ACcԸ�X�z���noBg�N	�2fS�� C�Y䶈�J躯
Y�ʷ�
S�֯�ؘ���^��yv��?�����ے���slueե���}�jS��V�B|�RjA-�����y�f��s��)��'(	�б�x�GE[Jf��4�?n�)Z=ؿ��P�ǃx"���V�X�:y�Y��ۇX2�"�4�]�+H&"���%�4z���u����c�	y��D�=�%c���������KJ隒�Z�a�Y�0t�H�9N��Y�9�/+�Qm�ϯNe�
�7���TJz%x�V${:Q���m"۵�]�x���a��ihk��/��}���Q4�4P�>e���o���X�����{c�����TN6@Q*'���k��(�CT��7^���n�3O>�Esgc��!ؼ�,9g��0�i��T�v딤�������n�z�5�[�Dj����,�1�2��}�x��\AT(��RU�:� �P䜩Qٴ�%��|�8?/����*L�BV�탳ZĈ�F\�����>Սӝ}x���8��O}�DC�F1����^���}*5с��D`�����w�Ɔ���6X�!I�d�"3Wdr�IU��k�AC �������[n�>�򁼯�.Z���6���@�1��S�fYD'(��<����l�;k���@w1�i�z�iTM\����,F��gN��t*��7c�С���䮞��8$ω��j��L.��KY�����լ�O�������'��
2@�C�N]4�DnZ̉.<��J���7C4������"���(��M1ʅfO����������4���X<w&^��JI��F(;Ȯ�Zc"�����}}Q|��GX�d� d&���؂G�z�{B�����F}��G<t��t�#���ގ�׏P�{�ĊU�Q1k�g�B�������r(�"��s(��phK��u��JH�i(����ϗv�ԭ�������eM�1ӹ�KU
\�I�?��l�
�M�5����݅��=�WW��9�f���.���F��hi�G=G�4V1���q��#�:BAU��ڦV��w^Gժ�axq�z���1�u�wpذg�ǘ1c�4
�'O�ɓ�1g�ttt���w�n��	�ї�`Ś��s�ьՎ-�mV��f�TW�Z&�tO7}=R�q�������Dgb鴠�|�%�Dp����`�W��˃��\� �ق��ȝ����N�v��Ez���݈���8��w���L����n�i��Y4�����*n��ر.@>��%<Κ�=;�a�ڷ1j�4��nT�uxu�&��b��I�7gV���H,iX6i�h�q�ÿ��&�ٝ0e*6��re��\c���"��%a&M�a��Z��oP���D��:b�[��$�'߸�����P�z�rBQ
;οK�"KS���b/�L�x���{�0�6��ʋ�`��1H�v`��6kV�?r%hxsӻx���R����~7n��Ԍ��Kgn�0�]��a�u8v�?=�5y�U��@��Y�0o����,����J1�hm
�,���4�g��y�fY��k��i"�����m.!i?ZچH�5��'_@��Y�v��,9�1�7�Ȥ���D�t��%"��
=����YS������	����_�
��|=���eYJ� $��t>��}�HC����:@��lλi�N;	^�C䖋��Jh	���-_y����6JV��$g�vu��I�"���D9�C��G���@��,J�;�5|��?�VB���K�7�gm1�H�"<v��L��\�g��"��'�7Y���oq��7�,��ʥ0�!����]���;n�<x�ٕxn����5����=���|��(���	�DM�Zp׽��o��E�u04�W����U���R��˯��3���/��2f4���BP��&�����L֩��$��m��4�p6b&̙�7����?��l�3 �&�m�蓌ȥ;�x^�_�^"r)������T\�54n����(�=y��b���m;y
�G�Łcǰe���%�	�EgK��%g/�yK �d��$�]$s~�k�����Y5����    IDATQ�iH�*����$�r\��Ĭ���}w��'8v� ���K|�N�Ĳe�D��{�╆����	&�����߂!C#���HW7�L��G�^�O������u�����=h<�C��=;y�Ĩ��&�|�F�8z��9R1l�bh���J�b=G�ÉNΚ3C�>�Ou��n�lH�bB���.fL����&h�<��aVwo:���O�b�J1Rer4S��
)4����/n��WV�����_�Eb�'��߳t�b�<y���Qh.'ʵ� A�ڶ�#ԅ
�a�:`2�P�z���x���=y2Ϟ-�������O��/|C��Ώ��㏶	j���&gu��oa߱�����&/�+���J��L����*�=z�L^�͍���b��݃".��W�@�V���i���mg���XCB�9M�R\��GY'�*�
�)3!�D�_��j�:���/� �]r1��:O⢋.�3z�̈Z{wOw���G����f�9xc��@�jF��+om@_2��'`ᜳ�sǇ��`�;�u0�>]@�Cj6�����;�3AA��KQ�i]�[Y뫚���U� (����s%����R��K�O���������?������6������Іz�� ��]c�$�h�$����]D�"����;�0��9����~ϐ|w���r��q�]&J��{��o����=U�j\m��,��G�o���&�E����1�h^!7p�I�H[c��M�l�����.�ˬ��j���jl�y �����dd
�4n4&��|�M��ٕwAYyo��λX��f�ʠ�����P,�$`"Cy�2�6�.�M��b<B�7�}&��ܹ{���8�_v�xt/�*�5;9ž�]x\�J�w��;��@8k�yQC���g?�lA��:���@��=f�:R1���i�ǌ��1j`�ܱݺwAC+�]е[/�}Q|��W"���0v�p\~�8q�
���2T��}!��ڛh�`�͇JoF����m�d�m�n'n�{-�d�7�"�� ��Pd}F��7��onmǆM� <�p���#Kd$�h~b�Z�TCKE_"��K�b׉�0�r�N���'@8��!�A���s�)�2 �-t6B!��DC�#�T��:�Y�Ŝ��㆙8u���y�;�p��9�t�{�-��+�.���"����uwa���Ҭ��#	�nl�wo�)̹�08s�R���D=Nb0�I��kf�o��ذv⡀8�雯ʠ��U"Cوt���Fr"�0��`1K�u,�1�ƨQc0��)hGq��_,_�xR�XB�"�]�؄�L���?qOdЅ�>�iI�cQ��X�7�"�h� �:�����;~[6mDNA��d��ǅ�::vF��(iT�'_�9W���ӧp�M��(�1��!����CR����A�k�Tٓ��d������&��7_��{�y�����8cF���\R��_D�H&�������$DZ6��>� j:��s�0���'����hECS�Lk�XX�.Th��51�0�4E�\�:�f�Aj��F�b	�Q�]m�c2C5ʋs`R�r�y匫p���x���ص������t��?pvn���*�O�Y��V?���x湗����ww��_L*��4v4���c��K�`�����<��(��C8�cv�^_ȇ@2��)C."~�1��=6h��dJ�XJ�u;�`��Ș�0�4r��aÜL���)F@� h��i6&��&y$�g=�&	�A3R�3nmF�SгC�ü��dMu���^������N�%��6Xq���;f2�� �F�A��Lvv�;���vɿ�ds9�������p��:p��sУ�o���<M���k��P�Ê�sg��w���RK_�����6hZ|�n�N���^��JkQ�g0��J�r�Fx�J��Е#�	����In=}�4�K�P�C������{�0�*-�.l�A��0*5@1��������lXTgA���T���/��>^u���5/���p2-V��C$?�;�4ŧل+�������D>��$��܀P[z�`Ҙ��{�X	#G��8����V,��+�4�	<�I�i5�y�`��i�<0�ho����[PU[����Bg�A�/��n�d�E%l�0�|Z��p��P��?�!qLϩS�����h����O<���8��);O1�/=�3*ax&��D�Mt���v���E��E_w�0�qN'��V4�d����K��{`��0~h�0{:����h?� �CO�ؑ�hljE����]Y,��֛пw�"�p�dJ٩��/�����WQyNj��J1�`�`*	C(�qbh�>p�5�^�A��E��jj�Q�� _�'{�!��k�'6�d�s2 �KK�Wb
�<�&�$�g�vY�i+�-�j�U(�-,)F�I�S���]��$Ȥby�	y�Ť����/ȷp��i�B�8���+~ܳ�-�:�A�����w�?���.t�5H��՛��QԵ'^]��\����`t���
�L�*�N�4I�6nƍ���$b�XYh�I�X�V�n8| �V�چZ���r�Mp;Dä��ͩ6IS��եшo�nÚ��j��8�jP�Gm��PIr#Y2�(�,�L�l�f1��N���dV�ޚs��C�i�<t�h�����������D��'N������R���g���\�o��*�&���p��9�6�x
���@]�e����g����}$�!��᱇�����Pu�4B^�H��H��`�H$�s���ԩ3��wzii�4Q����~`�%�@m�"��-鋯�_,	��*��?dI��zr�j��� ^��4�6;ڼ~!ّ�C�Q��1�D��	o3�wC[�a�s�;p� \:i
�[<����;��6		:��k����^����?�������7��ѓg`�)��Y ��Ɍb���J��5ǆG��vmۈ���˻A~��l�R*Gq�Ymi�Fi�	I3_^\}�;E#	<����lvCmv`��m�v�$2��b��$��8X���b#D����0*��͕�h"��'s+�>�iP'�ȳ���u���r�<t�/0����hʽȦ�	�w �7�6ֺD����6u1��+�d:$v�Q�m{���{����]�`��.:�R@AD�:�?ƌ��yA�s����Bi�"�Y�TaI1Z�aSPd�
��OǱs�4��#������1f�D4z���bɚ�P�R�l[�IǂR���\A��:7ND��#�xb-�F�(��\���'��Y��l����sB'_�z�!�,����hBg �����й�����:qA��:EO��*��);�s:��p6iU�5#���E�>���C��F<DN^�^�.�Z��*�Q)0���x�'��vH�ݾ};���_e78u�5��X�~������Pv��\$�Ń��#�m�*E:�����bV#�LC$%�lq�+��銭lF)J,آ���%��2�Ƶjٛp���i��iG{j�ly.j0��l(���:F��Nھ&C1�n�y.J��d� |�n}�%��(�J��A'�z�������T'��;v������F��<?����J�{�� :3�D#���cԜ9%�#��H�W
�d5����dp/��.�@�'�@o}3T)J�J��x�y��b�� ���[�2jx"ʥk69��ԦD-!�k֎H$��-�_V5Qr�@t:��c��Zn��>�kz�eEb�H�����{Ǘ�V���#�-���w~�ԯе�)zl2���*���%��ї��K�VX
�3푘�	1P�A3Jӗ�%WJn��x.�$Ց	�KG�/�y9B�E��nq���O�\��1�I��o����F�v����Jm@R|��j��z�N�F�A���(��Ҫ��$���HY&!d���'�M��G�M���'����1#Q޳�up��a�}���]EBf�JA�1m*.3F���y.�|~�,μb<��`���p��̑8фZ'�)��"��;���=�K��$Q��|�(Lv#�	%܈H���@m�[[1u�TA4X���0s]���=1X�Ź�&�\�#q��}a�4-5��H�DI"�[Y�ͮ�ƉU�Z#a�w�i�{�	)�Z��fs���݋�3'0q¥��� y�k�m8q�.\(�r[K3zW�㓏>y��fQ2�ټB_("�v�Ћ��"��G��0C߃���G�B7�͘��]
�z����SZ/3 A�#~�>wk�}�`<*Ĭ�'N�����@����
5�uF��ٗ�ph?ܥe��LN��V�����DZ>�͊��-B�j�I�>�˴qh�����7�#�Z��o�����OŨU���ըUhhj�?��(z~N~{�W�c¥cp����i+]�؄�����P��Eq�^��s��hE6����>������5r��^�'z��� w��bA�6:��E0��QX\ ���A:�@��*�3WN�i�~��|��QBŁ��a�y*�Y�M��`�&f'l��������E+C1m���AAW%C�5B
��	C��:�L&����+�9p��o*��b�n\!}��a��	=[�;w�T��;��<lu<�������'���>�`Щ��<d����<#V�Q�9��n�7_/�3���<�����lw��[9�۽�Gg^�F"��HMvA$N�0�O��1|�P�4F��`�%e8z�8֮]+p����`Ҥ��`1�/���j��H@Fk[��;���U���0��+��
�붓��Tu)��@E��)q��"QɒIH���H=��_������ ��ҥ˰i#3��B���]0�~}+�ȃ���ɮ�˯����ѵW%�^=_-_%лŝ'�yFeB���P�ݤ�2�x=�����x��:	ʪ����G8ER�N4�т|W��"���XK8��No��dC0��U+��A��d|�z�0�����otg�V����=��R�_�D]L�o��F�:k����:�̙W��Ջ���x��uDoT���Ч��=cz�nٵz}4�I���>D(��v�\�]�w�6w�Dg�5��i�ωM��-r���sA�݂��f؝N�:���~��1�p.��@����dz0�ܨjjFaE���Q���O�&��S7M{�ν�V-�?5��%~�lJS1hRh��h�����~�������r��������
�������Y�P�~�v���_>,aA$�1q�o�x�ǌǲ5ߡ��'������	aZ̦�b�C�y�ɌL4,�&�5�q��I"�����φ�onA���:ӷ������.�N�F�8$uVDx�4���"_�9�iH�$�Z�ϡ��H,ͦ��Y9��F"_*����ńa�����'�����	E�d�۰}�N������}��ӫ7\7O��Wϔ���V8s�p��)���{�ihA�憺�;f�i�����7j20#��z��n�ʆ&/d}�a�[b\Y�$2	�>_�3�Я� �(��F'�)2�4
r�X�wNZa�x�0�&ڂ!8MN�i$?�x��+��{==.��PT:�0��W�D+l���L�H g����BE�B�8�W����V�덦��a1s~����o���o��*���p��<��J|��d�����g_�|�FwL�<q��l"Aɹ� ��޽z�Hn�*#$a6��` 	"�Z-��;�l�2���	�g��(+/G8�\�1��5z�֥��{�4��? �6��'�|O�u��O,"q��.ө����%1[�f�+�b�b�X�и�� �wN��Oq�?.�0������d�_~����'��Yo�qrB�!��o.;�O�.P������lXu&!��Lȏ����-hS���q�Q�Ђ�B���P�f�$����3L&����ZS2���݋��R!z��N1�syH�x
*T�D4���g
Yi��%�XӫG<mmB 
eR���g�~1G�.���+*{��S�L��U���V��*� �7��Uk'������$��������x��[mɩB��A/|��g�!��!�z������ʇ�l�Ȝ�<���Ņyb�����*D��4�z� �1Hܤ��@���v'�A���C	�ၸ���Q���`�#�n"��LQN3��\��b!�G�n�9�Jt)-E$���gZUuN�K�Pܫ~�|%�5�J�c:��}4MIĎV�I����C�-�8ҡ� *�EY�pJ��V �m���<��Q�!�e�_��AM�+���ߒ�93��Tuj$CA�����|��(*(Dk�3����̑����.��D�J�/����,���RW�uǐ��`e�9�N�|�v� ���:=��ޅ��o���qc� ?'Wdoj/pT1F��`��Ù�&�m��5�?G.>+��x噐_ �v� 2�� �s\!�e��ᄬQN�
�5g�|U�k��5j��Kn]��idE��
�.��y��	�a��!�p�{��8�)3�ƒ��*���Px�:�QFJ�.%U1����6F��5�����
�D���F����Nx�$&>7%N	��N�"�GlJ�)-2z+�5
$���]���^��$�J3�ВLR��������f3�p5H�� �ބ�ݺ���I
�}�݃9��!
�S���#���#�0�@�̊��ޕ��?</iy9�������p��E�8y���bh�{"��JAg���=�c~E�������Z-�eR�D�����r��po�&H��u�,ǝ8et��Rȴ*��������-H��v!����Ԗ|N�4"8�UjiY�.���Fiq�H������7U᯿{�T���8]>��Ө��^?�����w�r��%ԨϘ>M��zW��u�]'R2Wn��`?�l1�o݃PF[Q��$m�y��JFż� �����'-tل�S.��!�8�H� )��()t�q�#ʖ�UU$/�@.4�c��$e]�����N4$��̀"���\��Y��q�,�Y����Y�WbpE�&G������� w���s^�v���c/��L���+��q�ԟ��|�-��ςީ$M)K�Q\n��T��S=I��P$B0�S��:���f1GY�ݝ��V�d%��Nm5:������;2�����y�BJ�M(������`�I�0}�����K�j�d���)�c'�����i���Sg�u�:/�>�}1j�p���a޴䝨�X�|%zUVb�eS���o�U�/B�Y��Ĵw�f�e4v��� �!䥓�I����`kr��Ch�Q����̸>:��R�@�7�O\�D�2����"���h��Ce� �Vˤis�#�Rd4<��I�������#�^�)Ν>���P��������-((��f���{Q[[//m~n�U��M�Q/����݁�f���7X��l;r~�h�Tĸ�lt)e*�����L��M��:��A�!!����æ�C�BKL<$���Ey2h��l?��lݾK�\iOK�+Y�=zb���rAщ��Ⱥ�z4�u��e\������@$Ik�h�9�)�#\w�5� v��#,-�&�h�9��ɨ>q�4�|�L$�̛w-
s���D0���6M/�Z*F�ā�xi��0s�c0F$&�r�hG�%�	Y� 2�%�ia�ݨ�S���J�L$C&}2$�OS�i���������{i��;�_6�Zq����{e�[�A���)��)gr�O��`A�dA��)�E�� ���{w̙~����G�e�����iGL(���o���߿r�U�f�La�S�*�3ɀ�2(چ�UuX�v#23R�b�$q�*)�B��̛����g���.�m���?�&�]���0�C���dv�Q��>}*1d��n)y]��b�u�^V&:\�P{߿_1�♥<���as���c8W� �� w1�Ԓ�t�z���X�.��E���i�5��ӏ���x d �x�f�ja��Qѽ,&�<'��f�Q�e�g��ђ��x{3�n��1�+�D�#��7`s*q�i��řQ���Co�US�ń����cx�rTt-��SG�P{���Il%�T    IDAT���_bm��x�װu�v�wp՘ Ң���0�����p�n�V|��*�k���WwY�I��E>C4,k/~/1�I�/l��Z2���h�Q�*���r����@|��YlVYK�aR�J!������@�;wWR$kg�0e�2��tI�%�Q+�`kS�bC�uq�Tj�� 7@ȿ��`	�e�����N'��NR����^�1����N7�=��N���'tE��y�p���C����e�H��BR�g��;s���LzI�����#F�U��!mF�%��
ÃEe�>p�0\}�,��߸ޡ5ʡ���� ���;oE��X�ŧ��y�$�b��թ0e�d������A���E/4�w~�!9x-M-Lr����EIi7o}�0Zd��HT�Ӊm۶!�a�ȑ�C8{�,���;v���L.���*i<`0�!�FE��E+�!/j����������yO�����d+�^�'���'��X�HXTi`�ؤ�k�V�� [^�9*|�2�?�L�R�T
yN^~�o����z�p���7s��	حc��u8s��H���'�Q�9
�.�H*!ų�KWT�/Œ����o���a��a/(��"���/�P(���B)��xH,ᮞ^�
Y���1Ҳ�Q�2PŃ@�6U��r&#��d�O@G?�
I2��L�Ŧ�]�UZ&����H{����� �����K�ms#A"�I��{�Ba����Ia6�,�55�)�p�998]u�v��a�I�WEO�?��y��d��D�PiMX�i�]=��"����ֳr���b�����VTv�)p4'z���1�����L|�D��y�
�j��5]@I�1_�ڴh[�L(���wK��@���H�[\��XK�Ѥ���21l�P��֠�DBc@�<��f������B��i�|���bD���.dK^�p([۶m+|>?�A?����F K���Y!��B�=��°�#�n�KN!���4��]}#�;�;�4��Q/���?�j�d6�;�`B�@B\�TEv+Zj�ĸ��8N�]�ѐp,,�E*�8,q�!jς�T��Y��	F�߶ �!iP��h�H��Q����a�B��!ߦ�m7�B��\4�UjHc�\��W�=���v���-?� �f��;�IR�
&3LN���K�G�����?x�/@g�AMюϵ��U8M�ԹZ��/Cv:�~Y�"W(�R8-���d���%ׁ��'�o��ݐA��$�ߕ���˕X"w�M͂(�}p����۫�\�^S2��O�CG43Ss��i4����s�c���ӣ��������� �rA��'�a��o���k@yEoL�1C�Z:V�;+�${�K�p�i�� ����%��ѵH:��S!�1n��b����N�픬u�ْ��ЕLy��*xgA�+)'t��w`.m�WY�~��I��UZڞ�f]����^U�1����O7{�N�6)��*�8��VKHN)���AR
�Ԑ�N3��8��C��!]8,�Y�b����/��I��j4HGC�	���iM[K�c�t)����q��Y>yZ"h�"d2.�˥��{�s'�a��~�(ַw��\N��_1�����}�^.���'��c�d���"�kh�__x��\��n�0���(���&\&�^�p��	�ܾ=�Ν���ݻ%���c�B��`��p��J�
�I'��1v`��O��	���a��%d��9՟�7�Ah�I�RzS�&�66������f��� я~��4���f�@!\�|w--�#=���/��jF������P}�͝'���=�u�.&,|�H<b�JC�ᗌ�y�����G���ر� ~���b͖��~�N��艑c�"/� ��Tɤ_֥�|���_���F�}�lv�x�9iq�N�LE&��o���g�a�R	��2N1�/�b�͗Z	? JV5�:��l��*q"��B�#�V'>ϱd�o�I$M_|�m����M����&³O=�h؋o>��ó�յ��v8�c.��+V��M$�f$�b�(*z��-7܈`{݋���kbi-����1a��hAo/�3��v2��@���hA��R���
J�7j����ZJŰ�2<�N����܊.X��ّ
�p��^8�Zh�1���LYnG�ci��<�<ߢH ����b��_)��hy�]p�\���V�<s�/��~}��ɸi�,��?`Đ!�v��b����+����Çb���8p�X�h�UW]%g���믿�Z���>�����o�|*�{���p;lR��T�$Ұ8sq���K;�
O���l1�i�y�&$�c���">�&>[e�P�hH����E�=4�pq���g��,T:�}q-��`R�G����RD���5�ކ�.�x��g���e����q�]�p�Ο���ic�T2�����A �Å��A �����d9EE�|=y���E|�z9��=%}Z�\G�|e>�Z�L"yd�K�������%�_�Cj�����v��iD��0�jN#��:��|o8��9���8���%�>IR����M+R�m�Ml�܈9 ��b*���}b#=v�plZ�~O+�\N!�c��B��.��6l��*-��ӥk�&�\���͕�h�D�]�Q����C�'"l����V:?2�:��i�(�g��BT�TB�u�E��.wV`U�����G)��$��b��V�C�DD0�.��]�����G���zmm����/;��}:�5�8�KA%�$��nR�^Y�E��s�⁧�<�Ci�=[Џ#h����l�j�%Vx�E4�W���P�"9�i2�R� �N1�a*T<��~�K�<{����͕'<�y�P�>o�����R�Y�\y'��ѽ+z������e��Q�S��	���N���|B��|N�>���H�KŐ�X��pv)���S����1t����%�����f��ѣ����~�U�f׻c�N>zD�mZ�r/����Tf���p�$���QdFzIQi$eBW|���0_�aGyI�sM���h�"q�H�������[޷�L��/_(����$�%~�Kq!n��z������El(�ΟW����¾}������9sѳ��?���^���
L�:Y�#j���_��7��k�}?��/�џ	<7�y�@�AQI)���q�-�J�VAq	��Z�?m�-'G�,�٥����#F�f2��������5˰s�zX����jB.^�z^����L��&,��s*��@�����E�6O �K/��n��\�����V��x���Ɏ��w�u2�c`ʤ	��Z���g���zSbSo��N|�h��.��2�۳O>�k��i���_~�����qխ�"j���_.��������z�j�7�Ϟ��s�"q������
!�>ٜ��b�G��V���&�R	���9=�/�mZ�߯�!wN�C���w&c�<PzDf:����ِQ��7������o�s�a�v$�9iu�#Ϧ���
7̙��|�)�]�>y
�a��U�4i2������A��}��iP�}B
i<�i�&>���^yUt�F_�,�	�%e=1z�h�2�[����W_����]!�8�a��"
:#*"���w��JνU�B{S-�m�"F�x��� ���=$+{U���I+�-~ʊ��8��&;����a�*��Cw=i�h����$/����v%�ڏ{�@�;��/�?�������U��@*o�ʰ82�+a�[��1t��9]�W�~�������uX��&����9cC��Ϩ�%DC��T��Η��4���q�Lۋ&��g?��"~��-HE|h8
Eyv�?hq��f�n}��I��r��<!\"�4�1U녴��񋳥���	-�0�r B���w�0p�ܹ��^����QÇ
1��qt��X�1b��f���p���Ί�dа���,�P[-���S`��7mEA�J�s	�~�є6��F��ɉ�������q����(���Jq��.����l�E�޹BS�M�b�ϱ�1���������_�m��-:w�,�ʄΝ��KB�]m��$ĹlA�`��".K�gO �?Z~q�i2��-Ck:���&\d�w��t��K�)ߴ�L&q��a�}8r�<�J䰐DĨSa��Q�Z�x�Z>ù�'$q��w�EII��t��NO����޻�����MH�����^��ӯ����,E��A�:y*��&F!�o-S9����2iX.���xZ�۰m�vq2� 7#ł��ઉP{�oߊ�]���)-[eQY$f���K�b��ժ����#C	�^�D�Kz|A�8y
>��3	 ۝���h� '7̛�M�	����

�
��"����k���K.��z��P؏cGa��s1��?v�4��qd�Q47�����º�[�n�v<��#rY�ܴi�$h0T�ݻ�����}�Q�֢a*�6W�6�d�M�Ìۮ��>�g@�ˎD�f5I�gAWg-d�Ϧ�r-���$��1�!��K�]6'�@,	�Ŋ�~\<�����$���q7m��q��W�"�c�a��hm�C��EA^��'�)�:�pX���k%��o�N=&0���Aر� ���{̹�N�F����%�Mx�w���8w�,Z�pݬ���0:l�n�v|�z9�
r��F.����4ױa�}~�-&�v�l�Z��÷ˑ�P�"�뀚je�u��Ia��@$��������<r��,p��׎4�",�3f�Ûޕ�2���[��Ť��}1l@�ݵ}+*�TS��}�"�������]�����^xA���GK�	/��gQQV��k֯GY���0�����g�(̹�&�[���yH�{��x��8{E]���ߐU@��i�;6XDM�3}8ճ��0z&��=?m���Eq_��S�����}6�</��9l��vª�E�Ϗk�W9��2qƓ@ EnaZAdt���4��$���w�H��g�哦H�ơ�q�k�į���vZ�=��������~��*��.t��O�`٪o��3������A\6�J��66�]�C5���ޣ>Y�9�N�!V�[w쁚{sr!xn�F,��S�H��sc�Q��5:yx/~�~��p�]�O+����f�/4�)��DL��gW��Y��9���VFt��C�(!��&�"�����ǀ�}�ڋ/`Đ��6�r!ű�x�伽����k�]��݋Ғ"�2q\9}�L�DF
��I����c�E�q�d�J����@� �+;�DG$�� �#��
����H�U�TH�!���%�1��/���N��UM��� ���/tm�׻8��F�ygxeq���lm���p���|����2�Gɐ��]�])��c�2����� �$2!�h9;z"������� %E�~����b�y0�@Hז��^�#5�`4����cO������G`�e$MS��qL&�sg��e���_� ׉��j8�6T���#/_/[.E�fw�����R��c���|�eX�`�@�cǎEQq)^~�5L�b�{t���_J��̫f�������#G�o�^\;{�|f�OS#ZS[+{�#'�� �;b�H¢7#"಑��p�4��܆��dD��5�NT��=�$�lƃ&�ov�Z���9��TQK������F���2\2a>��S��T�<O�tޜh�%�f�r١����k���?^~A�O?�;�{����%�}Рؿw�ͯѽ�?�p�1�FT����C'�ؓ����k���}������;��kQ��-����ܳ�c��زu'J�wGms�t�g��ђ�CO�K���z6�[��;w"I>���TYB����t��C�4�X�S	x�!�q�&$P�,2O��r㖻����;�e�n�k��h9��`&�Ɠ�����iƏ%�gNJ���w݉����%����Q�-���5(.,�#�=��{�#�WIΜ�Ŗ�1��������>G�~����w+C{K ߭^�I�N��o��K&^u���Yc6dC�eAo����	q�s�o����!��Q���;x�{5v.e	��,��#�N�9�Q����v�¨1"�Ⱥlب��ٻ?-�F���������b��1#ѭK!���	�����&��5�M��k�q�f�X�R�'�E��TWW����� u���1n���(,-Ä����G�����?�uuuX��+a�O�0��}�6X�x��̇�Q̩��	ӱ42�4҉�L��V�K}찡1�>������T�I�jf"�Qtj86��{���=��k&�vlB�,��u�@�H,��6/z��@*)�K�5CCw�H\!	_�s�Mصe#��E&G��0ѭ����Ÿ��g���I���z��z�Q��zx�~��Z|�h1���q�]�cզM8T_�֎ �=sgL��u[�uۏ���C[�V�_}���7=6�OdMJ&]���3t��07Ν���e��oj�I[�ՄL�C��+%��4��'�cygek�Nn	�,�\��N.�m9�����ɡ�i3��Í��_���ޕ����SЫ��^�9.�������>u��A� �墶�<��z9�͸J@:.���ŧ_.����W��}�� (�&\�qCFaŒ��i���@S(���l߱oXH�\u�;����V(��DN2��_�*����R���9��̈́�?*��<ǫ��mu����tٳe���	�1�� �����=��p��0���6�+]~a}+�$t�=v3�C����]j!�5�/ #^�x!{��6?~���q��I�>x=���rI��B!�q�M(�s����$I&{����n�{	���0{:�v2���(+�ƅ�޽S.6`\1�J,��	h7�
���h�P޵;

D�u��)ģQ	H!k�ě^����b�r��Q��苯��]Tv2�4zZ.����ېk��~��,�L],���!�����#�A
��V���9���c6b4&�#�4'�_�Ae������B�J���'�~�J�?���.x{�d��1��Z8~��}�'�� +���e=1}�Ԟ�ǡ��1�۰��u����ї�y�k�"���y7���j�K�,EU]����%_j�%ğ K\jע<q<�a�
�8�_t�Z�J
:��|7Md�f���CZ!�*�hLvpD/�GM��藥�<���e�v��X�v6��] w�悐q����w�=��ׇ�V-GYa��GD��
�q�/����Бð8��ۭ�ި����O?��˾�0f�(上�q�})B?��}�l�����.\:v����Ũ�7��
���ش�E�x�%zؙK�XB�Mi�jḬ(\�46��AGk��_���NߒH��ٕ��
�2�[O���\	ˈI1��q���貺����9v��/��^��(�����b4�\����1w������У{��v=v��x�׿�IvժU�ޭ�4ݻ��i��R�����r�*��_A�w6�CF��+�}GQ\w�8t� N<$��G��/�m^̾�|�d	��;fx
$5��`�J��,��׃q#��[�}�L<"�Y$�G��ʘh�$�%L��!w�8�u$�Є�����RRZ&�Vm}��޷E#&I��)��)���A��o�	�V/G*CNA����A2�ğ��{حV)�����ڰn�4[�{���NZ��ft+����;q�l�\w3��;���E�C1y�$l\��6��[o�}�V�Zc���ذe+6m�	��"�/���t�����xs$#�f���q�w8�w/�F���B>
r\B6d��0��x�˜�E�`l��5�P�լ5�$ћvט���#��!�!�2�A'��UӦ
9u��(�q��0_TTCm��˰h�"i��h0�io͢CC1i�d�|gO�Fmc�4�e}�T\���7���CqAz�������CAY	I^8t�4֬]�3>D�-�����pSv❶Y$�fW�����y����qB�ܡ�?+�::�~��V�/�:��sB�=[�%	F�T4k��LARl3I�X�#��d+    IDAT~���N�=���t��mST�𔢮�?����2��E{�T� ��E�Ŏ8��鎻���1?S%��$4pw�/����cG�kQ.>��p[�Ъ�h�P�݂P2"����/���.Y�d^r�baf�DYVn^��܁[o�ye����BX]ntx<���!�U,�%���������bwH�M)\9y�����($�T4��fNCs�Yٱn�U��Ւ��V��IA���tHa�)����n1��:w�),V.�7a���b�t�_�O�����N�P����|<�����`4iPVZ�M��#��I�1��=�����K���lt����V�U������t��ȅ)cFuUz���웥�q��yn!��cΤ�l�3y�h�k�T1��h�&tp� ԮS#��\��ԯv-�����²/>��8���yj��Cf񕵎��ҍ�x
A��Ԡ��:��I�c��='so��n�[~y$9|7;w�=p�����\w�l�7�a��-pڬ�^���uسw/�y9��|�B:h F���{�"�����1f�x,[�F]6M��m�$�>=�	���J�-5�C�D,���o�Es{��OcJ �LJ�Έ��M��P��z#.�=�M�WC��àM�sbJ��h�����e�*�>!oE��)��;aS��� Ğ3�Ha��1�/(�'��h�|�$dQ�M_�9�f�4������#�H���C���p��7J��7QZZ&�n4�����'�}��Bt�Zl���V���Ëo-���ygϜAqN�pfR��\2U���'������Jť)�CA[(7�J�J2�'����+��G��aA'��j�J�6��p��g��F"��3sa/�j��ђ��{E�7�����<4��s2O� R���i1����Wއ}������"AknkG(��)���{��S��r�y8{�J� ����O
���G���[LDQ�w ~ڼǣ�=��[~§+W���?á}�g�8@�x�|����ġc����=0��d�u.�g �zMB�N!��lT�7܀��6�ľ�H���Hţ�$(�h�̹6S��O�#�"b��:B��tBV,�Lu����H�5�4��ٰ����V	c�e��˥��#!|��Z�E�S�N`��m��Y�]�va��W� �rŷ�w�u4t���DͅYM�tP>hT��X��Fx�!8c��0z��ػz�]z�c������["פ��j&B�⢚u�FId����RI�w�[A��=��p���S��V��2g�� r?����{��j:���3"������HqRG��&�.{�0m���	��a�X�I��<D�rqgR�F�`6�t0R)�֒{b�vP
�R:=��.����p�wc���8z���P�N���hģ�z�T���˾��P��]�JD���т8';���-B��ٔ\o��3q:ep/J���y�=�cxu�8sr䂧	��r\.�+/A��;�dJI#�4�C^���f!/Gt���q�<Ԝ<�û�#��]��&���_܍R4���򼲄�{*�-_$�vJP�І���c��1��%˛)�)'t���~/��g�7Ԉ�_,VL3t:�G�_s�nx�~��i)�<��T��\�`�!�"䉠��+���KX�чX�a��_� bZ�2,#�$��i�w8rd�$���!���N���L��EYV�����7oām�䢵�I0�"��K��v�"*�B��qd��u&�x���2c�ß��f�I����a#���#͘3��|5"��<�D<��] ����:��V�YOQi1|� Z�[�;�G�rxJ�7�䥘AeIOh�:�5�c��7�=���>��j�)�����z�qL6���tÊ'��XJ-�;�)H�3�ho��w�
U<���V!��5X�cH�v�/NּF�����D���y�|>���R��+���>L�2.w>�b1�᤼_�3��GC�:�Qx��Wq��Qٳ���9+|��5���z}��	[ݝ+��������3((*��iW����DC�]�E�V	a��l�^�|�9w.�}���f���CuK3�>�MZ!t��c�aW��_MԦ��]2ZdvK�Xtѣ��<=�u�4
�s����Kh�V/M$Q+�{�09�p�@Rw��0�rQ_� ���^?�*5�q6@&R���*�w_�>�@$��G������*9�ӯ��ŋ�����\Ķ6����9s��o��ފ�}��av�BMn��v�Z�G��Pѯƍ�`�Ok��܉��'���bǪ5���Q������0X̅�GWPn�UI\9y26~�-��j���M4�Ly#V����N'7�j �y�w�f��Vև�xD�3�-х��&�7z|H�Y���L8�T4�_�|��c��o�[q�~?�vXMF�t��8r��0�{���8�Ft��KrA��L�0^d�z�^xH��6�=+��O?�ݑ�C�bܰ�ؽu+F������]\��F�e���hq�� Jn�~(7���]%�!��^�0��JBsv��d~'�nd,a:�΂>m����*j��v�/x]���o����d"T+���2�b'�+I2�����(	P�0tZ�A����~Vw���?҉��م1�N��(޼2�g셹-�8,�m�\\��xɛMV$Tj���}�1l۵���D~YW�H�(V�߇�S���K�"�ᕎ��Wa_ 9ynx�Y6�$�o�������+���/���K��6�3�<>���V�Y��p�/놌\z����ģ1�FE���[�0a�H\���C2�T$��ӯ���?nX��M#�d(�PP
�++D<j'$���BBP*��$�V#��gr��Ջ��N�%�.���'PZ8�c������w�u;�j��ܙ3H'��R��:�э,(�w�B]c��

$��p,���|"ᄰ�[�Z���q�ͷ�O?�4ى����3
7���\��@��G�(!Q������W��i�RR��'~�vo݆�[B���V��)UZ�]�]O�,����g���NΆD�*{4-I$30Y��`��ҵ�uQ�m��!����=%;��^yU��B�ɾ�,D�MͲw������(��zi���-��]�W���Dm�����j/��W^�-�%��@�'�ӳg^��V���8�)�I�^B��x&��,	����P#���|���5b颏`R'��B�Q䝲�˚�t�EٗR[�5B��H��Y��&;ⱴ�b�3%e�0���Q�~�;d��wx�0��ј7k����#���:��ݢ)�����P#���T"q����h�{�w��hoi���*̾�:T�?��e�t�/�=p�th�	y2@�h�0�h%���]�6� �	y��8l$�:0k�i@ޟ�&T|�� �p0�$N��[�,~n6�l@�N��9$���1u��O ���p)�e�m�|��)N�ii���9�F����x�[��>��#GbӖ��,��Z�����V^H�����Ƽw����a�F@G���3����æq��	���8�Ҥ~�E/��<��&+�g'>!�d�Ă�u�"�wݜ�ذ�[�:z�N�XG~	#b �!K�N٥�W�5���H�Y��?R|n���:�x0NU�&<���봚���1�M7݈=��)��5�4�n� �ٌ����!�2�����u5"o�-(ô�WJ���%K�$}�w`��P[�B��|�Ji�#F��3'�!�a�=�[ڱ��~�s���̴g��!d-V�?�RC9s�P�$� &#�r:�i2ЙHB���Oz��<k��w�cRܱZ�{��%�����%�&������B�EȂ.�xJ���R��� .�!/Js�0$���&����7#�&<&�RH�N���W8�M���	cd�Ǥ�(�bkX����w�pl�sYs+V;B����!��!]�<�S܀r�.�W��5��0Z�Tȏ�B`h�*��dG;?�"���D��d�g�af�9's�E!���,��s&t���F#�m���!�����Ps�7���P<F:�����4ZaW�uٕ�6�]<_�b���G.�\�� ��S*���gΖ\ߥ+�"L�6�E�g��c���F��\�L�,ZL[�Ϡ�u�H(��Ǐ�Б#���;v���t��/%4D%�NJ�::|��o�x�`��(�W�Z�BA������Q�B2yD$���JƐ�pߙFQa.fϸ��_�#�wB�I��%���#���LǧEzGR�3 �.�I��02��x0�$�QAQX�so�����G�{�YY^]���ާCz�i��bA�=��I�O~Ӌ&��h��H�"(]��0�������9�xss��y|�1��ʻ�^{�����c��2R��EO�(�g�/f/�4�p�DB��\��Q���;����x�]w��Im���B�z��`6�nE��}���]x��PZ�x[�]as�`�Z8"*��"���9��è�P,�g��i�N�Ξ���栵�V}�:-�J�,H(��rMr�v�犹�rd��T���Kc*8���'�ce7���"%�T�e�jH�2h �|��������+�Mͭ��}���f�-�ar�	Э[7y�(�̻���Mi�޽q��S��OJ��.*�ч�-M����D�&��H�`Z<ƍf��8N	���m�=kƌ������AP���PZ�w�s���k7cZ�d���k+I�K&�5Ԃ��<g�'7�1��a���V�%sߪ�(��DR�~���a�����'+�7�����f'���C��Z�vD	���2�E�����a_746�z�W���������.V��v�@�v�liv9��5әx��o�����*5�@%<p�=�lç8~p
�N!Fs-V\T$g`"ͦQ9������W+煬9�HJ���	�U�*C��@m�"M#�c�0�YX�v��Jvw�/��O(-)B"F�ŋ��1+!	�y�������!�Wa)J��P_S-�8��&_��g�ѱg?��v�\�F�m��Kڒs0��`����,�"��L�#W�͜���]~z�;�`Y��pU(���\A�#(�Qu�j�J�}=���=��P�O^
x^yٳu�؃)�ј/�r��NV�*艐.)�u'�A��"��HA��C�l�\�����+:�DƐ��2���D��3hFL����Ȝ�$�Y��b��}4Sy�g1k5B��o2��&���698x������@L4�����0��,NlX؝n���8});kE����C���Y��	N9,����%Cq��dbD�~̚>ϝ���[PR�h����%*����"�οO%)���4�h~B��F�h4�¸	S0`�p��P���7*����*9��Y����j��nU��*i�Y	h���%L��q6`�DgBW�.iq��n�y�eÐ�䒐�8�Q�o�(��P,����6P��w=��H\�H{��}�|�rN���V�O�*p�UV	<t����{�гD7���m��i�����^��0�.�8_>�-�w��sWq��aL�/�KA�GP&6elLi�9��l�1�$p�@f34h� X-!�jufi>ɄNƒ/�"���E�&c���<�y`'OgUB�z�Q�#���^�Հ���d������/s�ti��k���/6�
EM'B6
��<�BZ����|r�9|�P�(�V5�:�e��MG�n��x�j�9�e�}��iq�2��>X�'��/�H)�����!7cɒ%�p�]�馛D��B&�Ma�sM��V�Sg�������N?���=F��89|���ֺ���J��ڡ�y�ݩ�776઱�лG%-|W�FN�D@X��Ï�BNB%��ey��bH�5���Gɹ	0AY�x~;=Eh	G��fS��wj��1���?O=���.|K�(��<xu��٭+��ݍ��Yq�A%�=��ό�%��Ͳ(�0��k���Ğ�����=��Y�<�X��:G�>�[B��$�?�f�����@�s�lq�̗���Gi���w2D�].�¸���%����M#� �0wea�����}9�f�6���V�x}��z��1k�L:�����C�#��f��Z��iko�<1��0�фΕ]��TٱB���3J�ր[����!.�̟��R�B�d�QJ�E	ha�Ƶ3�W�y#u�(��i��9����J�.t�&!�G��Os��~�;O�g��/���/�j��ʂ�VS�����Y�y0�������[A���~�΂N�>H��2N�Oa����I����Ce74�b�a���)�<u�N�@B)��(�Q�K���bWj���Bkԋ{��=��0��qd"`�#Im��4)�����Cx��_�b!�$E�n`qv�F����	j�Z+�dX��K�b0JA��B�}�l�]8�/�m��i��j+Lџ�����R�m��(bZ*��p>�5=�U�Ȟ�b/Ĥ)�q��)T՞G<�Q��N6,h�5A"!��s)���-���$��K@�v��쨕��(?�D�jX�u��\�X�8y�J�e��ޑf9�]b>��Th������w��*Q�#h�e?�r��G�K���Ga�i�:���mF�i���U��d�+�󼺂��p0"���YH���҈e3���;�(*ņ/��C� ��"I�"ۘkR^��p��.�7�H��A{H&�/���RLNA�mme/�͐�t��]T�]UJA�Ӕ�Ł�W8D�� /^�ըG6D6�Q�F��x��G���(�g.�5#K���m���Z���uЩi/������r��t�m�59�JEB��Qe��g�z"��`�Ѱ{��a�v$T��6!�)�N�U���)8�V)P�t������d[~f^C�K�B�Y4�ɤR��M��=#�!I��tJ�R����L��^8�D4��&�pehL�I%`�S9W2�ip�I�����k+�B�.� ���z��F�yo2�`6
����4�q�V#��[�S�����#�ɩp���V!�R#��2�q�A��S����6\�'�|�(�J�is"��bϗ;��� �/�:aw6'���gU�N��[�}8v�,v�ދΕ]��$�Q
u�>p���Z�j%E)�1d�4�").��zn�~-V��gN����HD&t��\��kk�k�/�r�jXx�9��=�Mʀ��>N��4�H�V�R2�2�1�Ǎ�R�X_۬V�[���X/��G����7ZZ|�B.�q��P�ȟ�H�@�ن�N�p��+�oB���2�%���(�i����M4�莑��tF�5	��H��/I6��VA)Ā�L�Z�Bk2�S夎�i��{�{��=t�߹�n�����5��w&�����Ν��9?���Ǆ8�	�Nqʄ~B �|A�C�fڴ��/s�B�/�KTLٿ�R�)��"s���K�~��p�d��>�r,&[Q��X�믽=;wDCm-�
�n$�1��R!X�6ѻ.�x�0�y�Ϳm��L*"˖9Il<�	��~r�g��r�
a��/�/2Y�|y�lv� +��Nt:e?���b��o�8��ۈt4�l<����b�)|�{'�6�R�6��(N�ҕ����C0��
+��2�Q%�K�/��Y�s5u�g�3�L�S�f�p~�rҎ�������`K{��F!�����Rى�^���[���#HFB�r�$i���>�Q��k�19�����u7�T؟�ρ����h�aD4VB:2)�}�AH��p���y��7Ҟ�D�hiS���X��Bԝ:#;Sj���4���U
������Q�#�w�-�S�	�#ӊ)�[M=�d�'�j�u�]�x0)R�(�(?�-�ҹ�6��m,DgϞ��/��Æ�}b�y$d�s�%��S"Mf�eq�#Z\ʢ4j��n����(�L6.�$�p:,Hƣx஻��X��b �B(Y�M�>���j�r�������f�tT�I>�4�6��`�,>w�Ҷ8?u���s'�Q��������_BZm�����2�)M�F4�,���C���]�}�J�dr� �y�w"!�]�`*�$�,�fY&���Np�Hɔ����f�S
�%9X�Y͂�A	�\�l�S
���a}՘���    IDAT�PZ�u�>��l��Đ�Л��犀
����Wȼy�b��$���d<�^	$aZWeh�f�ͩ� ��.�5�4>*��ء�(--F��/��qm��*@{k�\�dZA,��-#zӒb'�I�ۻ�ZLV�H/��Eȍ"Nƕ<pj�5���f�ː@�1�{�T'�r��l0�4IeA������������ J@����7/���ܕ�T�H`B�R��4�C2	������f�\H�b��R�Y⪀�-�W~QsN�M�[lɋbs�a���y�_cY�zlv�)�p�,�wl�:c������%(�5��3��8��:�ЦT���c�B�� ˹�.�C��s|'��������!�NC�g�C��5a�?����Ѧ��W�\���Hꎄڠ��+脙x��:�?�.�N�\��̲��$s�;�/�l�	��abVC��\N6��h�I �FVg������1���ĮDn��"�g<a��έ>[��tF����Č��)v�]����F�T��y��1�>}�L��Ӎ�?\$>��,]���ehjm� �_px�s2ƐE�樳hJ]����d6J�f"�ì�SQu�(���3�BL"�QQ�k>`<0x��|��H&o˃��
\�BBlX�;u�s5�b��BdsX�|%�	!K"S��7?�0>۴�tj���p�Z��إ��(V�Z���F�Lt�삉&H��I
�_2N^ �=zbȰ�ٳ��\M���ȮO|�٤)ŐS���Hjr�y��e��	��s5	�z�^/zt���ޅw�zg��0���^HL54����:9y$�D�
EA�)[�-�(��8�Q�ŵ�5�3�;��Xp�|L�:�_D8�G��P�5�$%y<�رk;֭[�4��|�IT�w@Kk�V&��e�g�7Xĩn�K�f�Z��"Ƣ�����|Q�`�����d3"	�a�����F��x�I��C�{��B�t�U�&+�^^Z��hyՉ�*�O�_���MQ2}��P�VU�G�ŒHd���UВ��ŕ�^<�M���E��y�3�/"aܟ�ܹ���p��"O�4i�|���-E2Ō`���p��1��6�C1��cA�LQ����$���<��N5�1u�T�0��ECl[�"]�v�dq���w��f2�����H~��"] d^��܏��b�� i�����Sg�6Ẑ�iVԵ���=C�NKk���7��Tt�-�3�f�\�� �����{%i��r�9�r�����-Z1Zٻ�d��.�^g6�,�r��ڂ��Ƹ���L� ��4T����Ŷ-�p��1��*�"Qٱ��� U���y"��t�:��[�p@��Ndè7Ʉ���� ĝ���$�*�6�p!x��|�k`�¢7
r�ՇsFGn���R�l��U���G�!t���eeB�Kѧ�ꀹ� M��u{�z	0�V�r��_=��DYÀ�D*�VxF�m7�k�}9������
�YgFZE�9^�('t_���?�8a�w/���7�����?6GS�#��w�WYЕ(L>���td��ѱ�	}2
���/7�,�b_zEAgg�7�ZE 	�u�<�9Y���Łfo�xR���%`��_�X:*y[q����m�F�9��k���]�ƈ�c��;oq��2�+�ԩS1f�Xl߾S&�	�'A��੟�,�Nk��/�&�M�� yxHn,+/������:)�|@�,$ƀ~�QP�`Tk�cڄq8u� Ξ8��R��t͢(ȑӺNR�U��Z�����1��b'Š7Y��7�x6��,k�`:�J :v�$i�2��6/����I�Ɏ���Z>���W_���H,�N��ݺc�a�sǫ7b����-Y���T�����˖cۮ](,)C	~0+�vꅹ���I��)@��8''"?F���Չ�L��@ ݺt���7�D�ٳR�Ut�S��:G�[sP�f���c�:A��B'w|�t��AA�X��Nq��4*�Y��f��ɨ��p?|�f��d-Ə���"|��KD#\u�X\�T/���>�{�ZZЩ��((�v���B� ��K�8}�<��~9tｳ�����`�T���� #Gl0�T����<��?U"#�<`�����8 ��5`�����WC�(?mC�$�1,	���z����E���V��[���=���8�4#TE@�K����O�z�֯�6��]�nspl�Y7l� ���fA���F�����<��Ν���cas��O���I!vҜâ'7 �h�H��4��j�4n�e���AdC�%��n�1Cd����gd1�0��A
�a6���-S��*��<��w���i�4�Qi`w9E2�H�@a�Y��V���3.t�p�-s1x@?񌯾x��jT��\����ߒe�p��q.�u?�|A׈pR"IN Y�<�������}��7����DD")q�w�6�Tΰl⨐�H���Z��,⑄�9��|����p����dV��#rX�h�h������D��|����l��(�%���'����˦�`� ���"��ɻ�g�������(N�>#�O�ݻuE��4$d�����ę�p��-��V/<e�Ҥr'���\yxO���*$��c���8�J��(��ot1IeA'\�_&t�����^�o6���\h)��{+�k�en�A��o;�J!�\Y�I���NE.)��+��l�y�DYL4b��}kr'|,��ܮ�Za�x����Q�������a��r�:�<f����Xd1�2�&q{�:q��^=��Hӯ�CF��SO��ƍ"צ����C���~�#|�a�X�q�w����f�X�V���g�w�_�ԩW��j�'�V�����8t���}�Ķ�1r��;p�j��G�)�B��p�U�q��~T�<,�aL��R�)�,aX���e��!�If吐���D�D:��}�7��YamO���_حF�Q:�x���������]�v�%;�|u�6_ܻ�~�i�^&c]c��A��?���D�m*�./�|��窱��{��k�@}s�����%���'�J����SQJg�`H����셫���B��:'��H(�
3�&�(*��$�c��o���9�"gF�f�����+DR�o��C�����	9�r�+F)�|�Z�B�Ӱ:���-3�R�)uF$�A����}	���Ǿ�(
]n9�kΟ�kAm�[/+��Я_?ABV�X�z�<� �����w�ǃ<��Kx���a�Q�L�
�	���.Z}^t�; 1��H)��r���"
]D}AD�ðHE"�e�LmX��#�p�	Q+�׃ӝL�9~���r�3���_�b/�/�	�%���j���՚DZĉ��2�Ns�]{���'~�(��.��G�5jq͔)��>q�8��E�ǵw�]�
[����cGлo���;����7�v7~�g�Q6�Z2��V���).;2�5�p�:�IM�yZrr��F����W��.˱dѻ���9�@��.ş�,|�i����'EO�WB�4D��b,�
�âNR�9LF;.Ե#�QKЎ٩��h�\������vmیS'�a�����ը�T+�R<I~۱k�Ğ����6c�u�9A�xBP/z�3X��R<�~�ܟ�i�v��h�ښ`s���ʜ��A� GZ��*,w�����K��l�":�]ʋ%�(�mCQA�V����M�D��~����ZY�i�y��s&�g�X��Y����Z��"�m�͘u#M����s�
�����qXm�� B�,�PB��ǏÔ��!���T�h`s�%f7�գ��k6n����B4 .��J���Zd8aE[k�~y�q��=:��<�0���I<��m���Nȝzrw���^<�3l�?�|W�ު��7>\�Bs$9;�3k|�LM�Si�@��P�	]E蒓Y��8: ��s��xXX�$}q���{M(���7��B΃����M*;��$�;/(;�
�
שw_L�~�LX��AHk�e,$����h�p-u�q��qĢ��5v^�t��nW�������wP�^��DFjcs3N�9�����lt�v�ڋp$*0��cGq��a��47g�<lݺ��w�w����z}�p�R�KEba��(�(J��)L3��ޅ��g`1jD���vΙ��H�A�b��J+�;JXNj��i 0
�ބ���;~
�f�]������1��JQ��`H|��菹�fbӺ5�XV����|�����c"����Ĵi�0p�`�?t��t��)��ɓ'l���Q�8{Vصo���--���G�r����'^{�U̽qƏ����ט;�f�u���������"���BsU���ƂΟ=K����*�(��5�ń$�&%���"�̄ͅQ
ʚ��E�_U�l�\�.={K�:t�4T+��� Ij����g.�V|�1zv�_k+��,+..�_���Ȇ��u���ի*;uD�^o����c������
w�}/.5�w��fL��fΔ0��;�܍��Gb�GK�o�p���ڍ��d�1�(�x��t�ѐ3�'$��7�F�ۈ͛�J�+s���9F���s�q>w�_�O��X!�ѳ�� z���I�I���-6!Tq2�ޜ����N����7��f\3ER��h��m�#=$�W_���;�yUZ�43���3OK��9W��cFˁ����(*�C��~�G���Й�BX#9ҨS���Y݅(���,P�ښ��TAO(Zij�s�O'"�:y"�Z��H��!o�x1�/<��j%a�ɒ��0Bsr?��ͱ����Ki��R*�V�����$���Bͦ�<�v�{�Ox��?���	����8s��՜CsC&��/��%g��8a���W�I���[�ϝ<}N����~���7q�L�pX��� 
�S\���t�p�%a������l��1슈��:���`��)��n�r�;u\�p��`���@	�p-��ym8q*�02�E��K�6�p2��{�}L����HHrŨb�j�v��4b��סw��x��1�Oo�����G��E���p��I��iEd�MW0<�t�Ut��k���/�F�a#P\�KW�Ak��pXjDSc�DiG#䂘�7Y%'�"�p�:�WX�94+נ��{�%㲇#*e�\yȳC-���AMt��Fb��{��_�yԘ׿sA?P]���E�^l�gf���]:�o����W��t�!��5�G�B4���.�NUI�Q�����cp��X�)�K��	ه�|�.Xѡsǣ1��'q�ÏI�vCs��7��+P~�n&����F��X��/]DKS���c8t�_��@��r;��\�h�LPS�N��@�}Ί����KrC١�Y��%eR�X<�w���P���[�r�'2l�����w �'^-V�l�nU"I�C��ޓǌ���w���s�0T���(9ْ̗�4�ˡ<,�w�V������:Ƀ���A{�̛D��ޢw��Y⩢�A��ʡKw��#�c��-�׫�ߋ�Ǐ�;��= ګ���Q��,ڷ� ��mڰ7�x��V,G�N]d�%t^Us�����5�P�Ԋy���� ��,B,���sS'O��~��˯�wy��]�G,;-[=��bdԓ��A���zu���`��o	�Nltje�]��\Ag�/����G��d�J2��#��m4���a�lޱ��Za�;�~џ�k���9o|͗P{��H��1�-�F�n���ॗ^i��G�����������@C[*�T�бc�� �꛰nͧx�������zL�v*v�څ	S&�K�م��a��;`���%.��n��W6����^�̝	K��ܓ� �<v�����6g��sk$��_b����t�(��E��BX�1�΢bi��}Y��� Ə��C����o�n�$�P_'��O>%�>��3�������Ç�{���f�;v�@s��*�����x���Ψau{p��<t�0�4h��(V�ۿ܃�3�ûK�5��ff�����y���Ƀ9؆y7̈́�f���¤�"���i5 	�*v���8�or�n�y5������9����hA AE�QN��O2:T+W{�?��֭E$�Ť��q��9�"!)�?z�q����F]c��Fc��H.)g㯏=�=!�N�4�k����D�?���_��M^a�-7�=Z�vLfr�xo�x���p��G�W��pɻ�3-�AW$��k�"�����ضe#Ο9~YmB���b�|��TЕ�L)��<����.�2���j��`��:B��Z/�8�_9���̝y������c�`̨a��xm-Mr��F=>��#)�T����l&,g�w܎�����V�=���ko�Wq	�3p��?/�keE�Hn�$�����O�Ҩ�()�B�ȰF�pn-���B�LB�X9cr�����*�z��rAϑ��=�\/�0����v+i��;��S���ﮮ�pњ��#��:��:�K��Q��L*a&r�/�K����	�KI���傮# $�6���}E�H"��+�9g�LB��eT+��q��9��O<�ӟa��m8|�ϸo%˘0X<���ߋh��=�w�4��
֟��)x}����� @��)�D$�x�	t�����ѱsd�*��6��p����Oᓵ�1�$OX�����^:�w�-D;�ld�����~�x�8�9�J��S��4�$t���%�bu�z&��eL�N�U�*��Uc���U �*��ku��Tbʩ��G����!#F�g��X����b$'�%���.����a��U()p�ı�8y�0,��u���
��Xˎ;�����"8��[���O^���=�()+�Ac�=��G�֠��"�y�A�a|�u�X4��w��ұ'����Y�����������Nx��av���7K�a�n�7c��tN��XP&t�ɀ��U&#�6���$�J���c1��Ϯp(8Yj�h�%/��w�u����Eɕ�Vy�}p��Z�m�}�2�t�R�ǿ����T�@�ջ�����C���y≧���Q{��P�	�O��T.�anٴ�ĬY��N��`�<��}��ޯ0������y,Y�
��!U�U��V��&��<��$��$�s��c��DQ�[$�=�+�bZ��a��C�xy�rS��	=X&h�f4�y1e���X�X��&���ŸH�5x�'#�<~,:w,ŗ۶��eG���6�`�'�	���[R�X���g޵k�\�Y7�(�U����}��eŕ�����G+᧮�jø��ѯG,��]�4cF���l��Sg��_Dqǎh��V�a��X�p@&r�F-ҾI�GK��ʥ���Ҙ*�6��RԘ���I&�9�B�9�j9�s�(�N^��r���p��HC�X�cT��-�f�(u�p�m�aŒ��ǈ�`�+1�}����׏~�8T�,Ǝ���Z[ŕ��0�O�<)�����r���3�s�|�޳{���a�§Z&�7b�ܹ8p䨼�{���DG� ��쨃�b��#���a��sf��k��8r�!� z��\w}{BW�;��O�t���l/�Fh�6�COs����,�?�#���(.t��J�NC�;5��ڵ��Ͱ�殝I�[�|��c����
����	'�*���[�:v�q�'��}w!ƍ��#GIC�ɊU��k j�#4��X����RR��	�I���(h�¯�s�}"����X�9�;i�R��7��?�=�j���t�_Zb��SZ��ۤ�otE��ܴ+!wN�,�H@������yLq��C�|�Ť�(e��7(a�����KЉ�`�C��#�TXl���G�sח8|�$lN�**!1$:�������ւ�֋��o������ΨÖ-����RN����@�8s&���W^{�:����޻~��?��g������HA�8q"�-��ZyiF�+�"��?Q���:!�e��FJoV$"�4�4��aA߅ڪS���Ć��D��s�b����5�ϐ���Yйs$�^g0#�j�p�w���Ͽ�<%h�U��    IDAT`���a��O����!���oP�a԰�رs��~�gϒC����Ңw��a�����޴�3aj�3���칷����{4���O������a�+y	�̻ӧMûo-č4s���E%D�X�f�HF��},�Υ̟9�>|g�)�;tq��N<�3 -��\��CV����b�7-m��NRY"z<�ď�|�Z|�s7
i�HB Zy�J~����u�&4�7�CI1.�;/r��.21���K��RE����6~���8|��(���BC�V_�53�Ñc�$��'~$��k׮ƵӦ����߿/^|�ϸ����ȹ��o�jw�C�
�+Gh���Ю�.c&�7�B{]v��D6�NP�$����,-��ݓ�ϙ�\&����mZJ�p2�kn��x�e�ۜ0�\�I��~¸Qܯ>ߴ�.N?�T$&L�_�����QVV�s����&��믿Ɯ9s0z�HT����C����W^��#�**ǻ+�����
n�YU�C^���b�U��\�ޯ?~���%�J�dJ��*C�Ai���g�0�i(q۱a�
dRQ��A�3�˵I�Is�H���+'�+�,��T~%�*�,u��������ڜb~ԥ��q'���4^��V)�l����}������t��߀�غe����q)<6lBqQ���j�p�̹�l�Vlݾ7͙��]+�Le��~�8�KT{��J:��%˰��q8<%��h��ltz�,����a���ǆOW���q�x���m(t{��U
:�xBΊ�K��R�u���r�	�L#׆�'Z�Y�UL_�r���-���qӌPg��r�碃g2�%%�BV�@��s��A�0t�0�<v\�	'v6�7�4K�Պ`4�O7n��n�U�{.B���F\�d�Hۚ�[��1�W4��Bc����-DT�A��D�MR̶��]�1�q�(gz��{A�ϝs�9\r��i��~�,�|Ӹ�^UY���&��gj+.^�zk,;5��#U�d.��)�U���)./[�NF�J w���	).B�%�+-�8�1P�qń΂�	=_йCWأ�4(Lo��	{�Ek.(��ٷ`Ǘ_���N`Q�)B��I*�{�Z���F�Z�1fL�&.%W��en�\!:P:UW� �W��-�j����M2���ޣO_|�~�?�����X�I��Z�T"%S>�Ԧ�����hH���z
\� J"T�DC{�TB
��o�¥�S�Jv�Z�)I�}�s�Gqz�MŮQq$�n��C=�|~htf�]%"�>n<���%˗*A`����FBP�n]���o~�s�5cG���U˱���PVV"IX���yńAGX��@���� :�)j舑�;oV�Y��Kux�W���;Ե�J�B����C������܀�C�ʋ����8p��p���9�-�Bv�ZI�U\�h�ؽsn�>k�.B��Ӱ1��o:��N#��Y90�Y�5���%I��
�G�=^����ъ��9�⓵�}�W��܊�5w;�b����⛯va���?v��>�TW�v��k�I�R�<��`6]++1t�0l��s�.̽�61ܡ��3?�%���ॿ��AÆc	�����+,~���W��>��<�O�nG$�ЗRy����dL�2���0���u.|��{�dc)�dP�X$���|A���.g@"��Ӧ��FJ Ы���XV���[��� �˥x�gSh�P�y��������O�@ߞ=$�#N�$v6i���]�r�mm�Ҝ���?äcǎcҤ��ѣ'�y�i�4s:v뎧~��ħ��ڋ��_�@3���̻�z��r����i�q����)FcK@�#�*�Q�q��W_B���4Q���7���P���v�P�x,,)��ٓ���Z��k��rn�Z���1e����s�`�����~v�@D,dm�{Qdq��?��6"#���1��e%%���?�c�<�M�eE2q�0�&1�a��O~�SlٲE2�uF�8�Y�n�4�nڂ���92�Mҝ`���v9dűt�ǘ��X�~6~���O�&�OY������dN�zU3�����6���YX��Hd��@%��]١+��l�9���&��{�
h�C�9��$H�V
����X�T�&MBY��?��+ʠ;u=�qո1��_{�58HP�����ݸq��v�}��Л�D2��T�}�#��H�ҊO>A�N]q���8�VO����k�[@'QWi)����h��йg/x�QX.�	��s�J�<��[�{���w�/��C�t�.�U��ˬ��_��}��]��x�mIL�A� %$���S\��K8!&vaB�WHq�p �;KA�p�t-�r]���(&j11�<��!w���e���b��	��qd-*��������hhj��j��S/	n�wοgO��;o�!�(�v�t��uu��n4�!v��yd(3���D,^뛛�����8Yu��n��D�Z�����T/����sh���o���tB���
�bP ���1L3G��A}�Y��q+��/9L�ѵ��a�la�>]�7dA'�%M �H���+�����
=���K	�O��"�V�ڀh���}q�u��󧟂ը�pMm5@�GJY�
J��m~&N<�� ��s�{D��&5M�m((��O~�����`h�`0�QSS�`��Z����T��HD�\�$.f�~/�M��L�NeŘ�t��h	.�<)r6���+Z��� A�Z	z�嫳�-k�ɔ��~�t����w�ͷ߅u7K����F��Ɗ2o�]nE�عuF*Ń�K����WZ�#����b�¤7H�4�?�)Y�ojF�Ε=f,V�~�����,_�Z�I���@�Qo .�}��������U4\�G��DY(�.�b�0T���f���}�Zd"!x��E��+��bU�+�����W����	r����Q�v�웑P���w?��;G�N���+��4�L��IcF᏿�f^w������+1��ޜ�&|��Rk��7�����M%�j�,�o���
��0�Z<��/a+*ǜ[�{["�Ǧ���0�1w�l� �������N���Э_�#!�|>!�:m�kT�2~4
�6�Z�v�^ȵt���g4g0 R5ҹ�l��,��"/�w.���.ޛ#Fbǁ8����)�*m��*����g��ﾃ���Q٥B
�?�&L�[�݌��Vcߞ]p���:�ns����7ߢ���p�=hk���ƽ~�\������fb�5�\�n�j̜1�M�.�ˎ����V,�d-V�6L6�X�Fi��bM�f0�V�3�`���|�I�j$�R��v�B����+�t
��ʂ� ����F�n�jI�Qh�iL�/Z�gRbk<�O��б��I���&�gϞX�~=��:�W��͋�ΝQu����:�~�]ر{7���8r�*{�@i�r���/�SP�^=zcذ(�"�W��[eػzڵx�o����$����e�'����� ��'1c�w�.��
R:���ݪMz���zӸ������U���h�[�I��hV+]��ik�O�s��)��҉Kn-B1��Y�{u*�*�	=Ń��:H*�"j�+�����.�$0B-L�I*,Q�3'+Zv����a..��waݧd�iwJ���L2��}:�����%)Z�,��J�%��С#X�z��=�&^5�*�Hw�N'8jV����-�j�|�s�tl�`D��T4	_����n1K�֜g�ENk1&���r�UPz��#����{PW}N�Щ ș���0� )
<sEAg�ć��;'`r��\Eh�1n�u(���+`�9��@�,f$�`X���͞��W���
���_e�Z[��nlly ���x�2��P3�/�%�(t�V�����xG$:�
�X��P�tX���4�Z�FC���f1
a�!��E�D�d�n�q�ঙX��c)���L\
:W:,�|��A�+Ӏ��؀�m5�ܟ+�bի��k��w���b��O%���É�4YŔu��������Sx��7D�,rK�t��(��D]�%���S�8�E��5��uZ��y�|����D}k;}��: T�eFJ�|A�;y���@$Eܪ��Ѕ@�ꡧC��!� "�J%KFZ���y�4�5�HA/'�>G8R��s�e�9SR��we�'ZD3NQԟϚ7Y�,[�����(/U�)\63���~ݻ��?��zt��ۂx"��v"�j�9R�P����C��Ƒ$Lv��#G�b�%�:#����<�Gh�n!�1�7hG[S,F��N]�A�5���fq����l��0:��ۣZ�ꐎ��kmӧ���`�k�Q����.t9e���7��JAϧE�hI9�K^K)`9W=��$�C�.�KCc1#)�E�^N�?y�1,y��3q�?}��h F�CBmM���6���Pޱj�FVEE%8q�XdO�>�D'�T�?�%�|{!6o݅n}z�d7bϾ�����"B�e咖Hfw ��#�D/�,.��e�/@,������0c�d�[���j�ioH�R��T��!�a9dLX߹�Q����M�4zA�x_9�'�z�U4���CgGڛp�-��W�.���~�a��Cy	�'g��������UP;��D\���Ge��6����O�7�Diy̸�z<���(((ļy���](��޽��Pe1h�(pz#x�����r���`u��N�4
J�r<(��g���CCA�Hq����C�z6z�2�+����]��������_�x�۾���(�֕+�m^�b���E�'ɲ")N��N�N���%�P�C�=qɰ�l�����`F90X���#���:�����a ;֋-m��t��<�%˖����0I"d�ӡ��p���P�Pf��A⾎A!�[,K�e���&'��]a���g���;.:3y~������j)0�����L����4���=N���a� DJ^/]����F��Ҳ�0%��)c������p������F
�@9l��T �!��G��T�|6	q��P�(�z:�9���a�5�EW�e�
��YJ��f��f�𼹳D����A*�m'��6$n\�I���4z��3f��!k,Q��B��7[���;gF7yL���Qj1��ڤzt��i���6J�B�O����l1�Q`�"�a?�w�YӦ`Êe�!o�3.��N1��b,��K�Կ
�Iyn��0��$}1<�7G b?�..��{�[���Rk;4&��[r!b��G�=�vűC��'�^�Z�i�6���;";a��M`d��y��&�@�٤
5/�[Ͼ�=pv|�5�رS����6;|�m���:�Dk]�3ܕ��qG��#�)���^�@y������u�-�6�cê��Х�\���3��&��|aOq�bb��˄��
f��U�7��Ye�X�r-�%H����+|Y��[fވ7_{�U���j3 ������I,�gX1P�qⳤ�	*G�U�����Y0}�l5�/[���8F&S	h9E�B�y��R�4��:JB],��bñS'Ӥ$ӡ��m���
���D�Ũ��+W��L��&���Tii:�[�d��4 T>�'9�OP��Ͱ��?>��dJ���;h��4&I���Z�f#}�>���������Ѥz���,�IqA����l�[�ő��/5����7*�fj-<�%�.��6��?�w?@0��7B ��m�����)�.�K~܅���M���چ��"	���OwB摗`��)X�v��ka֩��HX	}|��l�*�;���q�i��>�5,k�:��M6�|��4�"O*MdO���zL�8������W��#
W��X&�I�^�sg�亘f��qO�j��F9/y��y�ر�KTt�1���/�;2*
��҄+�x8)�_�ˌ����oll��o ��V/�"Tt��#W�4:��=:SJ���3���d��ј5Lg����OT
z�R��挟��w.������'k�ecC	��F0�F�)k�(V���{�0A ��4�HEѽ��g�@"��êG<D��ՁX��#����S)�| ��L%L�-*�9�ɔhT/56�b��^T��~#0l�$,[��>t�@C!�0=�B&��zW���,����b����b៭��{��t
:#��H��zR��D�4�BY  �w:oE#(+,FkK�L2!t���Ƽ��3��@�OBCĮ�h��aC�ȁ��X}%n��hN ,�T��Ie�U���K�#3��B�z'lC��H<�X6�� �� ��86O16n�B@�\!Pi ���p�N�FBAWi��D?K�����R��	%�6hIX��%`f�C#�&1��"Qz�G�1،Zh��(��7���5��/-)Gqi�h�i�ASk��y<%EBhj�ѵ['\7uV-� ��F�I�;��B�u��d�c�H�6A4��9�r��4z8�nD�	Ixjl����{�X��rD�Y�p�M�A�4Z2D�+��F/h"@��J{�1N�9���A�x��VY)�a�Z�J�(��/^Į������n�ܛ��+B�I<���m�݀��"�pp��mj>Ks}<.�+:���I\�n�e.ڛ.b���
��G�
)�|�hJt94WL���z۔�rf�s%a�*��|��F��Yi����A�`���ka��-��b���]���{�E�)�>�H�F��(�f�4l������r�~�7\�~�:�*(Yh�C�8}�o|�A*6z�ل}(d�P8�@�W�o�д��a|r\l�[��R�63lFq2�'���n�fz�%(v9�XS�Z�Y%�n�ɘ�&�k�G(�`#����{�9�310��"ItZ���F]{�XV,D��Ks��W�J<����j��=u�xD,s�3MS_o馆fi�� fF\)�kf�܉�0aĘq����q��
�	)��Ρ�iE<�C�(�$b�as�$�ͨ������sv���K�0��bw܅w�y���f�A"���)+?�V+y|�t򣿿^+��4sb����gi-�2��*DFg���B8�AJmDF��ˬ����'��������1FB4�2O+��N�����J��hf�*�r^�Iq��*I�����gc���X��3\��`��a��M�j��3��� W�K�5���ɄK�u�S_S[+�eDN4D�#9�������R��(���>Կ
:>��ThM\Q�`ӥ����O}ˡs=�[���PV?:W����t�QNg	ŧs�;�WgSRЩ��P�B4Њ��М$ ���������F���U��"�Z.6���ʋ�d�e��R�t�ܳ?�M��M^l޾M:!_&�Y�zXxٝ���1F��I��x-G�p9\��Lbeh�
�`',����E9xN���Z&-e֦F[�J����!E��xB e~��Upzܰ�,�AB��K5��G�vy�S�J����o^_CH�~��}�? ��	U�z��a��CM�Y�](3�M3&K	c\64y��?d�e8t��CX�j��E2*)�DLd��&Z�.YYu����/�E)�B<�@VK�0��2�Zz�)�l�8���
3�]��"�r��.�/�0�B�g2H$���HgThii�{֧wO�"A�#!�77�dGLS��h����O�;����Tz������A�g����S|�r�:�\�VV"�Z�PVR�@(��� ��i���/o�2-�$f�3��F��A�h����$������{�$�	�$�1I���i�}��� ��i0���IP���D�a+6�=}Z`ߒ�2)�t#�f͙3�&I�Ub�b�90��9�7b˧+�6f�I�e��p�"��y'3��fJ=��(`�xCs�<$-rb֨4�����0�U��Ps��t�Z�β����� ٺzA�:w�����"��(�>���ʄ���5�I��H�+�&H��Nij���#C�x�ANT�Ǚ��<nA�x��y��(�Z�
�E��<����"��Af�`q�:D@�N    IDATњ�7ͼzu�,]*��H{�D0�H�%v��+�3����Wa����R�����D+R*�X�j�.�85M��i) ���M��1`�Q�קR�`��ƀ]��f�Fm�=��Ϸ�̙��q2�M.��D��&�qyf%�M�p��h�JA�F�l��Q�j湅x�����%%� �N+����8�x��LD�קD�>�����-��$���hN���)Qr�ѐ
*�7��T�$㊽+'VI )@ֿH�=TJ��b3�v��N7�Uz'��fӖ�
�mذ!8s�"W�F�5�x�C�z9��۷O�w�`ф���(��eC B�C�A�a+.Ż�W��� c��Z1k2��H�²�av	�maYL<��Q�%-mJv=����R�LF��1��M�Wi���4ʢ��_��"�V
:��(�w��o������<�q�Tυ+6-�8*�傮X���]�o]����SS��Gm�U�BK�4Ԝ�^�D<�'^@�ޱ�K!a|�kW�`�p��PC�I��\����&�U�hJ��ƆP��dw"���ki�F��7�V�i�P!_%����(L�&�&�!H��;|���`b����=yV��9�7�6�f֣Ki)��틸��Rb�AG��GKt�]5b�d��=�����S(�#NçO�:D��*�L�˪u�Bk���a�(�j$pCR��s?Ǉ����n�����F�!#P^�&{1�}8t�4�*��K��M�s���Ծ�縙bŘ�8�%�2K����}/�b:B�Z#�� w�S���2�nV$�Yes�rCD����,�ڠSkj�O�����d�PP����W&d�������qv�W��u��w\㮄8A4�H)PZ�V��Է�mw[�P�^(P�H 	b�]'>�3����s~7��y��}7��'M73���9�9�`TK��f�~�o8u�0&�4 �߇x",.R��i��F�(�<���{.�U̩�(�HoE��D~R���GEEC3~��k���3<����Z��r�J"�J}�pC���gx-����u�F�����J,��W���� ��b^���~�z���a|K���PH|���Cr��GP뫐���𰬾������c_{�x �n�'~�;/>Օ�6Æ��(	���H��T�t��6&{eI 4!A���CE�y�878�w�o{NoM#"1N��/�6��2T�8keu%I��tN�B&&�����0�7y�h��~`*��w��32E�4�u��]� �!�Q�5`,n�~�
�mf��kD!N�d��p[�p��P_S�7^~u�^�wv�ɔB�$��JɩҨ5!�+}�pӍP�L�y��̵WCoq
\̂�4iN�M���M���'�����`���D�0��F�-Q�Pr�$���#�~�b��b@�'y"�\�rhJ�2H1��(+Û�,|��Qb�!}E�i�w ��˳��DƦV鐎'�hZM9�J٤L�=�1n9�$�,��0;Ki�(q�Q6TF�D��4'��}�il��r��W2H�ek�E�)�A�k\Gѳ���t`�;��\�M��I�b�����ݻw��7a���EF.u�����[����Ƒ3�q��9-FBKC�/�c��@�l��!��m1��K�0<2(�	�)���V�K$x<o9��)� u�]Y_�-(G�}^�u&-J�8,�~��%/�n�(�����l:qn��_�״�4�"�~�	˂Β�	��I�����D�)�{jB���
�p��Hgr�0�+��"I�R��Ov�݊@0,/��D9�J^X~��')�iD�GP�,���޳�����"�����S�'L�m~MFqTc�ȇ�LX
�A#P���|	�����à�*���>!!�&	O�8����҅x8�g��~��pT�Ƹ�K��օ��#8 �������O0y�x��9�����%C?������g��8��p��b(ݛi"�Vԩ�e���F[\�r���AXY��SI�=�؈,���U�8}��}Л��̎Q�mxu�rzT��H�i9Җ{0y��#���4a1��p��g��#��?W	)�K"X$�
$��P�����wݼ&�)�kMd糴�������-��Es���@$��`d/����K�P[U�|&�Հ�Sg�~��k*��tQ�'�B2+"��H�Zy���IFE=�dq��t{��څ�<O�lW7,�D�J:�Yг��A���-��>q���H��
GY](F���� O2aw�GA%aaqF.���Ǣ�ʋ��0LZ�*�q��q�:#�����^s��D�~��(z�>�>���!P��Kf���ض�}�P�t ���{��t z n`*�'�WX�dѓ����O����F�,��n�3�u��Vj��_�੗�����4�PD��^rr4�Q��PȦG�SA�4���@f"6�q2����M��%w��d!c>�N�4Z���/( ����d1aP+�+�N�w��)6��]���G��v�t�a��mpXL����t�"dԳ�/�f�Is$���)azWjL�c�bI+A1FWZ��FW8��H�b�C	�x�3��4��<�_^"B\;��Z��_NH �T¸�G��Q�E��";&Q�͢��6��l"�Q��A��,xz������.k<��,F�����hC�D�M�R�ظ�����#�A]@�?(�S��g�=��������!-��iN�by*�	C9S O�,#�F�f4
'R��ufi t���)	�h�s0A$h��<˴vV��6<�N}�t��J͘g6\�^���Am���%�Ƭ�3ס�B_Fd�B���G�%��ߩS'�s��f
E$7�duY���tV�rO���j6�
W��bJ��,��MA_w�u�+�{5���N��ݣ"m��:z����fW%�Ir4�)f��������%S&bɢK��F�����2�F�%�%�����=X���k�Lx��W�~�'Xp��2w8��F\��:L'Lz�iʔ8��M�eҤY�iI���?e7$��ߗS=��}F$^�:��I�lF$�73���k��G1��_�e�5�"�N�9>�`֯]'��J��~�\{��n�@,�o�����Ne1f�d��=y�0�B.�,������b<�g�~>zH�㉘����5%�N�,�O�g�����[�%�ؿ�J�$Z���J$sj2�H-=C'G�,6�I�i��
�<ti�[&uC%B����l>$Y�({�"���ɾ�)i�Xu5�H��#�{�]���%�:�/��zB�E�O�Z�C:BC������q��U���i����Ahx ��a��@6��jT�p���u9h6����4�d�y�Դ���a�(THf�oD�/�َ�� ��)S���]7�}
E����{\ٶR"=i�Akbj��z/'�q#�T��H�c#Zv�cP�Ѡ���a�/~�C�z�8w��^/�����O6#�J��o�y
�����&ڌ}��`՚u�3pV��A���'E*8�Ho��n��4�B�?�s~&�x 3N��\.���v�����0�atzਪE^g�^Bb��Qs,�:�J64S�K�X�oq1'�` ����pe�d�"���"�H�=2�s�(p�B©�,�bw{͙���&ìR����ttv�=t$��93gHDꩣ'!����1�D�jj�0��V�	mgOc��K,_�̣�S��� J!�ʈ��4%l��YF�2s��q0��tA�4�x+�0i��%��nҠ�6%F0+	h�e�y��0R~'��4>b��xN�!&&R[���'S6�b�R���d\)^Z@�K����DV��r^=�á�N�9'�HCm�B��J�cz;���)SkUm#��j)�kk�޺q-��
)1��˳F�j��dr),F"� ��ZA��pa�+��21�h(3��F�67�-P�<���֚�/�R�ٕ��Et�b�ϵ��i�j�B���?�'���@d2M_��|�h4FAK���΋�U`)�u1��l�Yk A�}ج����8mVe�ֈ��N�\d�p��5Y��%$�uT&�R�s'��::7B��������������Z��dA�t�'Y۠C�L�$�a�H-�y Yԋ9��at�C_�����n�~��#,N����o���W�:o:
,���?��)S���fJ�o����nC��4�����09��[���HFA�]�M�N	�\���9s<TI�*��B�O,w����Q��e T\*ʞ���L����G �J��Z�p��at�]�C@�����#r�i��ȃ���7�l�)9~D�RGO�A(���Z�TV&�zo�̚��K����I�l�c��C���l:�!��@�|��<��_J�"B�� ,�������ko�U�]�,�Fo��SM����d���d/tE6	�>'�@#�vA�h�y�u��D��H�$wB]�ި���t*./����7�,k�������������@G��_�k���ϊ^;���=�e������݅�b��V��(�I�_MQX�TR��t��z=?q�ܷ2�,q�ܜy�s�:n���b	%=�vt�w�u�,��e4�V;���#�,��`��z��$G)*� �r-�Sg�X+:o5��	YӯA��&�H9ir�1�1���n���F�υ�z 6�(��D�\��<x�}}R,oY~������։T"��;w��HFyzT�7 8<�Q��P�͚*A�~�����`�V�Bp$(HQ���Ji��O��K.�T*�׋�6�����	�ਮ���F"hM2@d��YUQ��fE��S�1�%�������mї�I����."�yQ~�ȡ�e��n��XЏ'��n�z"Z���,�{�B;^x�w�bٽc'���*��W�Bog'r�<V~�{�dD������q�������!�WR������\V't�U�$��X\6�U�>i��k���Q���Վ��K�hD��-izTGp_��D�5���K!�q�C���-��>БӢ1�Y#�ˢ�4���R�X&�l��	�5��� &6��w��لT<"����X�a��zг�����:�X��r>�'ZOb0��[)�;��Hv,f��ǂ���)\%���r5�d�qY��Qy������EU����3)Ogs�i�h�>D�@F͂����:I@4����Q��kݴ�`�iF������.׬��ә�$K!y�u�dA��0�J����P�D|X����&���@<��d�̩S�s����78��m��@���QpTT!�/"���\�yR+��I��e��Y��85���}-��̈sB�X���Eq�R��즩�V�B��ߑ��u2�a�si�s�rܼl)����"�LIg�)`wx���7ߐ��Jkȹ�^"Nonڹ�(ْ˯�b�g�~���􆢰��������`8��v��ʃ��QD��Η�hp �0{�puZ����Y�|)Y�����
�F#|���iI���r��?���vlG_OF��d�V�)>�7^{��a���^8��'N"M�����.��`_/
�8~�L5J�qL��������w�vl۾]���0�y�
I:"�DOj�������/�|�����-P��2;1�⭐ɜ{��o]PC_PCé�'�^����v�P�Z0L��~N�|A�T����-�b�����Ĕ	���}���B?���H��wx�K��v�^�L������X��&��\2c._4�]�7�g���g ��悚/r:�H`XvǏ>�%��;�U��]��ف�{�ݽ�C�?8��-\�H&Hv�}�w��tz1�H2}W��tf$r$A:�L�� ��H��4���/� je5!��GgQ�����yN\
�*}��C�@K&	Ij����c5��)��{�´1���m��z��q6m�@0�=ʿ=�\�x�R��tИ�B��p��U��e��d�XpK��O�]9���4�ɐ?���si
�*��/���_V�?��e]�gl��8x씸6:뚐.j�ߢ6ZP�	�Z1֐wL��Ə��4��r��N�I�2��랋���!�6<W�ʆ5�I⺥K�<��ӏC{�#:2�k��K����NE7͜����˻�c�vL=O��_Q�q�BG;>ټ;����p@�A��c�(��}��➂ZMS�(�����0���v��݈��n�/�m2M΍�3��w�=H3�#�m{`8��n�.X���$���S�AԈ�#��3���%�
ڞj%�,"����U�b�!I������\�����2�&�4�*��� ZU�� F�4���o��R�;;�%:�w/>�9ӧb�������p��y��lF�U�W,��jKX��(m�e*��C���۷o���V� �e�^~F��'N(ˇ38{���U��֚�0a
4�JĊjd5f	K�0���˳��g���kR:�p6�Kj�p����I�͉�J[N7�2r���U	�!�O�aJ�N��ˮBh�[�SfNG�`B�m�#���
_~� 'Y�f6[w�ƪ�7"�)�ꮂ��}�	�2�K'�:%��k��JAg�Q���ڃ����ݵ�e����FHq�VŦ�?t��偺XЕIDx�~�Y%�Dg;�&�Y��ܶ�}�t����۔40gz����ٝ���Q�U�hG���S���c$Uj��}���e�0;�0�}�fBg�4`���yx�4�Ɣ�&s���5��+���H	)Ca�}~aKE鮩�d��OŴ�5�1�߃*�W/Y�����Y�%b��uk>ׅ�#��M�ȇ��3�;��ƛP���EuW� ����U'�^q3��03��aB� L�e?u�H:3��"�F#�͝-�9��f)yL�<�.���}���6������	%k%�1���-�ڂFL����l���^��:��9 Uv�Z��h�XU%$I�)�3�؂h0 �+�XRv��t_��n�Ԅ�X8w6~�DK��ı��k���`1;ffN��'�z��!ES�44�h����3ȥ�:a�������8~���
�(H/�}`����je���55�^������̝�u?�[﭂���N���Ȗ`��0�q%[�RB'č�T�{!+��tG�%��g��8!�r�P�FC&�W�59Q��n^�V�F�v��O��
;*6hr9L;���7n=�\Q���.L�>w�ur��/�`ͦ-P�(hH<BllV������.Ǉ�>��-[୬RLu�����a#��MPuU�X�Z���
�>o��Ŗm;�������S׌4��N$2482ʂ���l�d �ӛp��H�!aE�%��Y:�|N�!<S����$aId�7��zz:J�Ë/ <8��3&��z�!?z�:�z�:�Ofp��	�v�����۸v�"l۱m�=X��I�ղ��4�E�hL���/��~�7|�[�U&6B�V�����z�}�lv�j�T��y���1��IHkn{��6m��]{᧲��C�>�Z ���7���JH��^Y3�hh��N�:��� �k�LJ�)�k�0i�h^���pP��U^�T���������X@�+�ذy36lމLA-���`/�_w{�A��$�I���J����S=��6݅��ni"&�jD�ӂ��������QY׈@4,k՟��Op���fP�#hh6'��#_��XKsJno�u,Me�9��8*�[�s��I �SQR,����sCD��OPW��.��Wb*C��Z+)����}��1>��5��+<�P��1FD�~ە�c�5�c���@��F�I�������
a�'O<!�)6x�
֬߃7�[��� ��:T6�H�	�
��5 e��-��)\��
���)��O�N�`��%�4�p��.F,��q�]a��t.bx%N��$ �x�N�Q?���
7�-�[֯C,���E�C����x��Ԁ�d�"���O���}R�����Ҍ`8��h2]2͌y2[�i��F�Y�����N2�XX �x4�Ńx<)]����}���9    IDATȄ@��@mCX8w�L�,��ZR�fN�!Zl(��y��@L�p@c�Y�$;�pW*Zg�/��Dq�cPC�?�TQWUL�d��x�q�F����l�XL1��L,�?���I��Le��k���%x����V��#��c�,F����䪬��S��6�	CY�&،ɷ��g��l@��G��"Ȓ�$`���HG��=2�X4o�b>X�>�L� ��HHZt�gO�_x*j=V��\���P��"�N�̩������a�ͽ��Q����(�����Q�&��'�	cF�_���ضq=��+�Bޔ�Q��s�^фrgq��)ddWI(��g�ĉ�����3u2�٨�[�%r�%��GM�[��w��*�7���̸.@�(_��8}2��E�zh��` F�s4:��1�7���d�[XFb!ͺZ�+��0g�d�kl�O�K.����'`sy$ ��l�5WBU�aۖ͒��98g%J*�����}��8��ކ��N��6�/��Y�!|"J�PdΜ�2���!YY�0�K��./���Ϡm`1}T� �ѣ�7#O�F��v���d�˺�ɘjdɹ((.},�
��v��@�29WX�2 ��>�.�5^'�47�����'�s�,�p�X|�d?�Z�
[�mE����@ۅN�ttbҘ�X�h�X'2i�w�\[7�C2��6 ����C���i:|R+�[�
�s�`v�ȡc8}�����c̘Q���J*�}z�9̾t�<G?�տ#F��E:��i��k�$�6
9��.�l:�^��buB���Bx���y���{\�@,�I�V�0��)22�|:���j��I4�k����`�XΞj��næ��p�TG����;�'��n�a�?�X8�uk���\;��:���ظ�t�?��̟�G~u���;%���-��}�OX��475 
�9..��O&�"6!��c��������fh�d�dU�1qH��0	���:Τ3R�S,�Ez�Sf\V ��s�H��ff��wS���a�ˆ��N�����O>����Q����I�
X�Í��ge�b��Cd��}�a��IB��;��:�?��:�°V5@gqCc�![�I�Q�_�7Q4�D/j-vo$&`1#�}ϯX���m���[�M[�y�k1�~j2���.�'�$���+�$��,��Ka�X����_��*�E:B:�A�B`�-���C�� �јs�^�M��H� ���>���Ã�V}��Wp��]���&�S���d��d=@��~4�pUT �L �nf��9��l5YP����"J.�F�\L�[��@L�8�V�ƂK� 	K<&���t���ȁ����G$��R
Bм�ͦ�ǝD	��d	��I�l�]a�I�*�����$���P]S#�3gNbh�Od(�Nd|��L�0W\�XaF���#��H,��3�ą���+Z�5����� �_�!�̔�l��E��H-x2p�M��uk	��"˔h� �O6+��u�L��i�ƌ���Zy�C� V�\)�|���F�8��ܯ�mc��F�y�I�Z����hI��-�K�
2$���[]����[�xK��J;�*�ܕR�$Sr:��s硩�IҼr"�3��|W_?��44&*�k%3�8�$_)Nq\�p�a���L�D�F��e:iq��B���7��f\�Rf޻V�J���/Dww7Ο?��j��x���:�q�*�u��HJ�Y������@4��@{F1�ˆP�yy�l\��$�Y./��<�r�8+݂��<�Q_�/,�q�'�� 7� ��w��8������/�ԧ���H���N��
Y���Ű����6�c��.���z�X�^2!/�"�!�Pٴش;%A���B��S�'e-a�q��<̈�mB��=i,��CsC%�͝���|6�W��x�pDP�p(��S&`�9ذi;1� �P@�Y����p�e�GĻo���Q�ر{���h�)B��aV�>�O�xܸ�[��ӭB���Q������3Y���ǅ�>4O�����g�ޘ+T��.Yg=392$�r?,�4��]N�gA �b1KS�g��X���BC�h��3���%��ɺФV��[-���`R1���>�x=TF�4�;w�B00��Z��.̛u���>�p#R���t�+@TH���٧1���wlI-M��E%"����`�4��,��<V�|��m�o�^�?����_z���5ɒ%�V��D��9�5��'G�.y��s��\��WT(*i,�oPy�բh�9�5�y��u�Ѣ�-W^!�j��m878$�إ�����P@}]zBl۵G��W?z� �j5�_�&�ӦMù�lݽ�z�)�a��Ac��Z�x|���qBR�I&oq���щ���<�P��غ�����P�$r*��ٍ=�t�sWI�ϒ&aă��@�92�S	��Ã�����|��H7�-�HRIw�i�Ġi&HAw�b��g�^Tx�B[�BN4�z�'iw�]sI���f���XI�e	����[-&	^��$�*����*�0S��`E���s1��Y�]�x\�X�w�Ŵ�d����u��L��"��+�x���$ӓjfUs}���bG ��?����	Z�ٜ�j�j��J��(��T��2��+ΖL��g1�ӅK���KJ����w���;v��'��{*+��Գd"'v�L�Ӫ42�ID"Y�&=bT1�4b|B���Ȅ-,PdDi��e����(P6���z�51��?oƎn�ɤG_**�x��W�	�O�Q������h�))̤/j�I����'�i������Y��1��,��j���-"ea8
N��w��N�`�:�wǍǘ�c��(X"4�D>u�H|�D���Ս������F4/"�Ay -o�V��#I���ԋ.4�\����b�ݨǊ[�����e˖��;o�؏� N���_�h���p�ş�+��'�|,F)�I��� 㖶��%�*�[d8,R�DH�PW��n�bOe�7�ń������%q��.��r�V]=ݰ;�BȪ��p��I�p��!� "z
v'U��f6/]�f��I/0;�4y��b���;"���ϝ{>wlr�x���I��{�q�4
����J��a9t�>�*�O;9�9Fh&v�ъ'`�M�"Il|���P'o��?C �%����D��&Sng{≨�׹�6��'���3��F;�b��>lٶY�.��@D�x>��Q���:<(��H���}��sC�5�bZ��4���$(���(`~�Q�	��i����`�g�?�M��61"���rB�)I�v��)�
yT����q����o���!?�t<�����.�h""J�OoD�E�nj���FBu�p�+`V��vn76o�����e�d2�@*�@�	��,n�en��f<��ou ��Β�ݴO����G�/94;D��t?�&
���x>��DH_g�H���;ׇs	�v�}��,��"�6#b�$J�<,�F��(Fp;�A����]},��@._0{O�i��8$����Q�K�]�|A,����p2�HAo�D�]U��;w!��š���F�I�Nx�em!:�������^�oO�om?0c��ݯ&5�)�RЕ]=�RiXC�le��2��b��uN>�<��CAd�Ja`�hw�D��]�Yv����r���T*�Wz�[<�L	�"lB�2=�Z���T4Z ��EQ!�h00@cC�����Bc]���K��.��%����u�d��᫪����ť�/��];v
,z��W�W^��ko@oW7����N��@��3��f�O$�����%���-�C����gJP�0&�G�+� �3�$b1�fA��hG���a��D&�*�MvE�� B�!47ԡ��D��MwW��N�[�Z�DU5�B<I�2ШM�G�ttob���T5�#�.	얈Ea��`T�a�1�!�@(,���f	\#0�5��?~�[�	O�@<�0��{v`�ޝ���[�p �T�1	���N��(Uy����m2I�J&at���dFR%�f�C�p�[�yO&�Щ�ª�����<�1�Q��$??G	z��G�R�̜,nh��Y�	�q�	����]!�a�2�����)����T�*a��QH�e'�Md`�X�3�x}�]Qp���$f_2�<�p�>����y�FL�2��~����mp���)�Ҙ�W��XJq���'���&�Sdu�N	���\�� ��NQ���i�������{r=T�P��.�i���P��"�N���������������"�N�d����g�K�p���@�D����4�t���9�G��<�B�$�E�C�Ų|���I$-͙l&#�\<u�5صg/&��_��ߠ��aP%���.e��<��>+D��D���U��<���d��8�#B�����S���4a��($�rơ��lO�w�J���J�@��U���A>;9�9�?zkk+F��+���]��Γ �$�TV3���)W�ÀRdZ��+,�2�h���98�Z+g0"?��aFV�|�;o�#�����5��CW�_~�-�l@ׅ3(%c��2h%?�$��XV��h.��d
.�U�"8䕤�A ��_U���l���h�񠷳]��� ��ۏQ����}tblSn��.�^���N������B	�D*�����7�%�L,��	�!�����kE�2։�/�좥i,*i�D���Q�'�a]���cڄ&��PaP
s^��֣�q��y�9�t/j��aB���48�&�@5U5�(�q����Zh-�.D*�`DE�8�6�`>��L��]�a+���]oe��I�g8��,���7j���2�d��C'��_
���}n*���.��(J1_a���y� ���*��j��!.�fL�tǸL�^����A�Mf��T{܈�B���p��IT"8��sfJ�4��&�Y`=�LK(���ӝ���Ì)S���0�7(���qc��X�ɧ᭤��JP�H")�4w�{�ƬK��ʫ�a���2I54�a�ⅲ��n�����V�ń][6a����t�]R���b�C*��!=�L��	�L	��f��fq&e&L��$���E٥�m�w�w�Ȝ��N�â3�5c�\���lhJ�|}C�LrDT�Ö��}��%m����ڄW�؀����4W�B�%�^����#��J��WءJ�F����Z�{mu�'Lf=�;�c���S���t8��pPЗޑA +FCAT�]����h��'D�^�'Tj6 z��V<�)�#�()}Y�P��ILm����j�IcB�Fr|��j���s�_�|�1LY��N��;=��1�$�~�ؑ��Q[S�Zo%���Ct\��/���Q�C�9y��±0f\z	����hlnQX�C~̚=?���n�`�{�u�<NI�b����xT���!�Di8�S��Ʃ}����F�`CZmFQHW�:@� H��i6�,:�Y`��%!�U��dL�k&���G�,ݴ�������������S��R�8�����VS_'�4����т�`P��lz=RY¡Jä<�ji8�{���ʗ�*���A�?�'��m)�� n��6<��S��4p���m?��(E�DF���������$�BU��H����:��u;�dh	I�+���`X��
4�ʦQ�����/O�ND�j�Ϝ���fA�h=�w�.9?8�gUy��`��	��,��������g�cl0W�4Gbv<�w|��3n�9g`�oB�]���Q&˕���o�� %�.ĢE�ahxXxG���[q�-7a��w膏�DV�}�aTT�d���Y��J���BH��0�}� Q�p9b��Ø�Z���ZN���������^Qc}���e1�w�`T�Xa�W�<�� �p�T+δ_@"���n����dj#QI6@�����Q��޾>9���//"d��kV�E�S�����'aӀ�X1UU͕�q��8��c,�:E?Z��[���/��֎:�	���\�BFL5:���r��N�����v�Fw���##,�:d�J��!��	]V��D����+�;u:�`��������[���`��W�:ˤDI�t���B*भ��	��JJ�R�h��Vf�B���Mf���L�5q�)�8�ӟ"���V�A"AhhP|�k��pP>���.<;Җ�:��ø���n�R9�_v��
���������[�����X "���'Na�)Xz�u�s�m&��5��Վ���������0c��\&t����2�{�vd�b�iطu3�;�Q�$�p��:�@�ܠ�-=U�֎@<GU=r^���.;�����-�?��	���2���Ƒ\����v!���v����D�E0�BoO����LR���|��ZO���c�1g�t̛1�v�ƅ�gq��!�А��j,�;F75�i�(��>=� v�8�K]�Յ��/���D,��M7��Ѧ�eECh�ps�� �����уhinBp��%�].�E���>O"��AE�Q��x��ېU`��@�{m�4H���0�P�I�֤f3�A�zz''S�V�B	��=,zar��b��#�f,h^�sfNG.���F4�0����8,����PP�K�յ����B8���N�{O��'ϟ��o~����<��KbaI؝�
S>\��8E���$ch��!��K5�|��-6�u6��D����P�:duv$�F4zaM�*8MZdQI�'1&�щ�dV�k�ģ�l"!�P/9Iibـ[�6i$��G{SNҜ���'o�њ,�XR{�9���QY�Տ�V���n�� G�2����7���ĕ#۵����_~��^��L�ƍ�ر�q������u7\���z&=`A�x�&�Ǣ),f%��gL��d�uU����:!^e�F��tF���F�PW#�	�|��0�TԈ>9���^X��-*�?N��M ���T[/�\�#2���:"�]ND�q���d��J��J13��I�lVBWI��IԱr6pՖ��k=6AD5��؜r7�`����oE}�ҥ�TV�^�W{T֗�>ـ��_��`�y)�D����~1Ꮊ��˿)��d:W"��0�����&W�|f�wc#C���g��󂆃KNt�Dfy6��N�7_B_O?�N���c��='����3��bHd�bR�����H�%��6I�49�˯wy<����nA� g)������]�d3B�Y�-PYux���qt�z,�9]֩�=}�4�Śu#����M|VC	�dL��*�%�B�P�� *���1�D�t./�%3�v/R*#r%��*B/1�D��:K�*>��y1mMcQ�PLª+��ջ��e�e�}���Ov]������iKH�Q�,碬��.t!��5���]:�tRD�,~��� ��c4�bȡL�$�%�q��|�0��A�_��ͳX�G4�td7.�
K�ö�1B�����G��������J��b*#��V�Q<���
TTסqt�����e��e�������Ł�,nL�!��$���I�%K��&���_{'���֍�u����'M��y�bˎ�h=}
�&�����n��Y�Ov��$�+!�+�~�b6+�L|�Os*��Cr'�"�����,�
�CC=B�8���r�r �F4U�"��ͯ�j1��W������~�k�{�VL�,F"55�p�L�B�0fBd�PL�h�7��̸����u�<����G���]�p�d��:�(s���I�q��kP�sb�ʷ��"W��l8ŝw�-/�-�f�XQ�4
��\��'ΊG8#w���j5rH��q%ޒ�zV��^W���d%��,�d�HRȚ��D+�i%́k
�{d�bЫ�z<������iĢ#����[A��Μ9��s}���^4��¢W�t'-��j\y�?y�G���׋��&L�>U	�]���ȫ��Y�0��!!T6DU(��p�U"=�`x�W�@�ؘy    IDATgP?	�0jt��w����3�$�n��08=�$)j�A���s��+��a�OQٿ�`oi��]�U�%����&��=.ӥh����-Y�ٴ46�^����ա��Y�:zT�&ꪪ᭪đ���98��H5MM�5��T8�5k�j�p����-G�xg�BD����ҹ�<�ze/��J�)�ܿ�6m��iA&8���������_��\����cY�d&s�3I*���3|��ń`�/�k��Q 7@ȿc��:�!��֢��� :b0�3�=��8���XW'9�L1c.<���|,��-{zp�f�F�d�����dV�s���`� �e��YӦ�<4�`Ҋæ��ʬ���~\{�X��:l߱5���B7i*=&D�?Z������eW`�o 9��Ya�ۼu�`�F��LbXR5ij� ������ b����/�+]6��1dS�0���F�@Y�A
���Ʌ0����\��LU��Q�B$��Ȑ���i�B`�Bd�hO\�qp!ǂN9$:��ƌ+	�pP�M�]$6�칉��e����	ԌOC�}9.ڃ�3�c׎�8�z
s�,�u\>B����tEŐ�%��(�y�U)�B/�2�i����Fd�"��euϒ�G�{:1�QVL�/��3��Ê����l�bll�����8��r���?�������=��޺�Y�u<�O�;�F2B�D���{�rh7�W�X,���Н�6�E�<��/v~�x'���c�}#3�c1qú����p�Ԁ�{�������nG��#8qh�_{ƍn{$����ش~-lf|n��Z�Z�%���,�Bc��ЅL6\��z������������_�X�wW�GN�xE��n��L'"!�/PuN��:�_{�a�_�>Z����P_-/";�-�n��<Bʌ���üyK��5�o������J�x�`C�d��p��f�t�,�$���-5�d�C���v镸���زi�<���z,��j���`�ڏ�T���}[,1?^�!����عm3���g��ag��V+�Q6���n��i��ՈF?�M��-����6���l���܉%W_�o}�8p���:qUSi�<!`���4���+V܌k�,�sO�C���y�Q�e�)�]� CH�2���2w}�!��n>=x�:� �Q�XN(:d8�ӿN�Պ�DKJ�D��C�n[ 08���qcG�G�����1x$#���RK\���/����@�F��L����g�Һ���Lf�&��B�o@�E�4=�َ�P 5c[p�wb��m���k1}�<��o�z�&�
4�1��"�­`XM!�DuՕ���qx�n�߽�dZ2r&n��z�X}罕"�,�������?�����+o"or ^4 M�2����%�2W��5��:ѧ�fs O��!��@�#'�3����f�?�O��L[�bA|8������s���/��Sǎ����<�44t�S�DP?�V��1
E�WU���`��	�W�p��E���� �?�����B���hu��/���<� ɶ&zz;p٢��d8�g���p����Z(`��ْ"���^��i��� �	��zSyh�^�w����n��i�A
-o�Ɇt��P�l}ڭ����@� ɜ\�Q�b��GKs����;��T��Ok�`��|ᦛ����b�$���ta�}صo���8�zaߎ����1��9��wVڐ.d�t����oo��5�����e�_���t�`׾}��p�ǌ��5k?F���};��|��6An�S�W�F'����ń�,N�y52j'��)4L��9��/���J��i��irJ�:�1�N��FW�BNLXؠ�b�B>�������$�0lV"�\2{�O�$י,y��k�����Lq"��G�Ȅ��(��)�����I��0Q3"Zá�G�p�6@m��K_�"�?�{�0~�X�C'2�d�FbadbCH�{�4������K������3"�Z%K���j-�[��ஒ�!ew��%�_�Ue��t���'t��Y��[	8��z��7�����l��a���3j�8��N�+_q�aV-� ���h(�_�r.vTe(^~/�����p1p��'f�o29�UU�����Y�JHVL?"[��W�s���X���s�M������H�V��ZO���-8s�FUWb��W!
��d��;�t
:�gj�n�]��ڇ�D���Oćw�?�
��R|�i��	Y<�����E���y���9��.�=u
��s���:�d.%��_~Ed^�'L�܅�!�࣏?.�'yJ���+9��P	 ��]�IN���Dor�	�X�x���tw���ʇD,���G���ݸt�t�;y�����<���N9v S/��S�'�u�FԺ�8u� �:��_��N:������j���
[���+nB���ƝǱd�r̿j�|�/�q�0J&R�*52�*'X>���˄�p0��/�/��g��2�E����.ÌiӰ{�.�a�9Y��C��N�,����K��އ�ᬮ�@�C��ƒ�'WD$k��g�Y�����(cִiB"Q�ҳ�3�c��Y���y�V��w�w׭�1y,^���h�̻t����$b����� ���jءF��	g^��4*�.|z��������5k����sl�u������DNŀ�ro-�JZI2�8�A�/�Ϣ���K/
��qWCekbj���f��	I����/�VU�W�[��ڈ0�S?Wh�P�b�d�|+�[:iQ�Q�����d,��jjjd¤Eosm-,���dz�|&����uUX��=��w��`d���o�ɕ���-�h���)��1��.����X~u	�Q��n@��	�&���/��N�F�l�
ҁ���X��n�dbMDXq�uXq�R|��/K|)�(D)q���[���){�s:`2:����G���{���_\�H��@�/�+�э�h|%B�V�&=��fH��Y�X��*郪F��8��Ev��:�N�on��<�"�*2)��,F��@E����ʹ	5ۥQ��]X�ч��͜>{����s୭Ƭ�3��x�s/�"��˔{R�C�����e��\��r�����O�w�FhK98�8��u�c܄����+�q���w�̔e�o�H<��m]0x*�U餑T洲6�����)�J|�ȦZ1�)�g�7�0�u�=�oj������2m�K�B���è.��ѣ�<n�0����"dď-[>��I�C+�Jyi$�;L���%�%6 �X�CQ���?�d[�$����:)��!	c�	S�E��vZ��c�&9�s��4	�5}�,QE;q
]]=�,�R;y:*j�����	��"Hl��R����K�3Lyꔀ:��|IK{�,�bl������4mt��kB��7�m�KVm�JR��Rܭĭ�	t�LEC�����)��?�_�,8�
U3��,�"�L2�A<�sr�bQ�����)�q鬙������{E���c¸1�2a,6�Y�/?�I��� ��V�_�|2�|"�&����`B}=t��Lݢۗ�Q�	g�Ķ�{a�zp�-7a��F���x��a0������B�,��M�ė_wƷ�E"��c�ٸl�B�0J/���{���0[p�eȕ�ذm7N�<���3W[�<r�Q܎��n��IB�T���A�����B�͏<�tz5֮Y�	�`�q���p�{��?~gOCW~��w�u�<�}���q��|�e+J�
�8�4�FSE%T�4��6��j$0g�#�c!,Xv
z�j;n��^�d�_�6���Ţ���Δ�x�e[�e���ٳq�5W!�׉�3�p��Q��g?'�O�oò+���CGN`�Y�i�I���/o��O����B�Nl|�ʵP���������sgLi��F��@@�s������
�{O|�֭��%3�a�;o����������ǜKf`��f���_��O#00�B8�E�fb����f�h290��.��j7�w`D[�]��u�پ��1�b�8z�/���"y�^���$�-�d�KFa7��_�P_/��ك��_�V��[طc*�v̞9O|�	��Ӆ\�cg��ӿ{i��ŋ��N�d��S�ب�x����)oe8�b�`��g�,���V����f`��c����02؍?�]T�l����q��1�p�n�5ȹ��q`�>�N1�z��ВȚɣ��F��p�>����c��͸i��xg�'�v�(����\2�0<2Y�ºf���l,���g�%���sO
�[0m�d\�dv�؎����8x��������'~��?ڄc�DC�+j��@"�yB,E<D6�����+������XƷ4ɞ�����[�#@~��lD_���Mjn�}������C�{@�y����e��+0��ޫ��&��DG�lo��lv�M�����v�DRL)�%YV�V�V�H�Pb/bE! �����^ֿ����s�9� 	L����ק���؈Rٔ�z�P^ַ��-]�m�~���j������Ju��)���7k��������_�ˮ�Z��m}�����=�b��=`G&���/Q�џ�hD��;}����~�C=��i�7+��jEk���t�E�u��)U��z#ڵ���?�7�b|��U$7�F'p��S�|���vD[p�H��D��h��j]��>ǝǎ�4>>�>+����_�VB�]�Ho������JSǎ��oM{D}(��� xU��z�ݺ����~.`hb�qR�m�@�M�c�)�|�R���9u�'c@��v%+�VC�\�UW]u�>z�G�ۓ5d?8��y��� �:�z����l����xZ��A���HW�#�S�Y]��Cү�z�IH�G{?������_;������?_��7��(��N'M��~m� $c�\�{M��ڄ�.�˙� X�7ې���9�kE�&eth�٭�7i��5:��^=|Dw����c���k���}J��{t����~�G���z�aӬ�$�z]������K'������f��η���K��;~CϽ��U�������6�?����/V"�7�2 ��V�r����j��:Ԫ4Ԯ�@�ҕ�]�+Ƶ�0���k�Է��]��6oݦT���zTsK���l�_)V�6��_6p1�x!<`�4�ue#mg�܁��t�e��g
��RqQ����{�z���f,V�?��:��~�����T*�-�G\đ|�Fr<���Xi`�0ɞ�^�:�Z<b`\�؄&7�����_�O�Kz�gԏ��R1�LDY��CU�iB�n���e^���4u���N�4-p��M���4B�s���n���h���k�+�飏kTf"cI�$�Ng��AbGA�K�rq^=)|�v{�[����MW]�Q���?�n��_���=Y��mo�?�y����.�h�����G�� ���?��gϨ���ɞ������/��l�U_�G:��@A�۩j.��S��u��o�^�����_�:Vl�j�'7�v���}y������Ȉf��Ѓ�oܩ�|H�+&�zr�>��Ѧ��u�wj�X֞������X�H�	�]���;�q�vÜk�x�����BH	������7n�Y�/����^g �_|����;��'?TqvF�o����z���i�3Oj�p�v>�����/��N$j5�M�W����X"��h�g�RH�x��M7���o���u����������j}9E��Y-L-i�oH�ڲ*�EE[u�q�-zÍ�����ƹg�����?�������$�/?�)��c�)����;ޥ�}��:tj֊���xz��]��v.��ܼ��RȈ:�7Ǥ�^V�����>�\s�U��W��7���ڳg������������s����m�efg�~�:�0|Y_��t��:��1�=xX�����'�z\��'����gzr�.���[��d>�_<�W_�ڷ����w�ٞ�W}�1�Z�vj�e��eu��ߪ_���������Et����QO!��V�O�R,�ԓ�������?��N�/�s_���'֩�0�]���iG,��ܫJƲ+��+�m��i6590�/��w�m�؇}D^�ݬ�cG^ѣ�<�t���|J{�}R���
�����7_��}�I�\S���h0����z��̽��?t��e�{�'t�5׫�N�^gn���Y}����ν/iWQ��q�͂(�zAN��������7�A�����U�����^]�^�G��ޯ�ۡ����m�@o��}�{���}q37?�t�6��Y���nx��K��|@f�����i-����{�W����?{���գٍ��`��hɉ��ڥVP�
O��¯��?L��<��e���V�*�����zDF�N���W�l���ܪ��1��--�ꁟާw���z��ߪ���/������#�v���Z����А^ڹS��c/-k��Ԋ����kr�:M/���ܴ~���S]t����>�g�ݥ,�H�%T�RXq("�{'��,8�ח����]..i��A=��C-p}_9vT�V����B��*h�z�������8����zص�J���Zղ��zmͺjr��m�b:��l��];t�y���?�_�^z�z��:v���?�?�n�*�q�{Q�3~���<d��|*�!�c)��L[ c�mZ�e�^>~D'g��S�X�F����R�����#����e���&�t�-S�T����^켻:�&�pӍ%�=��G{���q�1�H�X�;���{DMQ�~���^�#Al-�U�HP������Q+��������.rAq�����}��_��箻��}�z��w�w�C_������3F����_����(�՚;�ឬ6�ݨ|4�LE�&t���je��q�7���q����koԝo}�����k߿OS��E�wC��Db?�VR�g�h��r�uZm:��ߪu�6��HkW���w�����k�*�k�ˇ<j'�#��@E궽&���A8�^�N�ؔEO���'�*o��׿Nw�q����޷������U6�ӧ>�W��?�#=���:s�������V���_<�o��W�83�t"���T1K���-N+�lh��\1��j%-����[ubaYW^y��o�H�����5ik��qI�+M��*������8��ccz�^��#�ٳ�E��o��܌�~E��{�דO>��~t����wk�R��W�u�f�A��΅'w�#��Mz�a���J��#o�Ī��6�t͕W�=�K�����.����]���'�}�y���+��/Io����曕j��jسw������<��=���]�V�����ɸY�U]=�g�^�����J[���wޥv����G>�����z+j���ܼWY�F������O~�}Z58��{�衟�LW_~�~��[O��q�'V����kv|�-�k���zf�K����d~Xu:t�I�v���#q�ޤ^��~b=
<0 [�#��n�����ӑ�jV�%ǚ��7���~Ww��=��c:�o�V�i��a���U�^����~�0�*����b�&���� �QA�vS��N{]sۻ�֯���e׽N�0����;��X;^:��R�w�{a{ ���P�+{R�u�y�������j���m�u�e��]oy��Ɔ���s/����R*��Ukt��W��ٯ���;�%�#p6y�*�'
�l7������D��	��a��o���O�ڠ����~~�g��,����F��	�*�o��
;��1���n����~�w<砅f��#sgg�p��%c*�I๋�B!�sR�
�Ƃ�����;u�������GT257��˟߳{�;�k��J��o���C�448�;�~��}����II<��o�]�k��G?����8�d"cp�S k���tqЛ��*FF����޼��~V�Q�c��?0�Nc�ٲH௮6���c(M�R��o��RD�[MM�����`p	�r��CfP�@C�sb�
ڼ���H��_���Ɔ��{��ܱc��Z�q����:�1K�    IDAT�����~�k_Sy��\&�b���z����J}����O���`#�+����_�ȉ3������7��������"�n��}����N�L���Fms��0���H&5<��jq���"�j�kڐлX�.n^'�� �
ZX�"�r���m�ݬ?�����rQw�q��������}H���M^e����ڿ����5=;������z�=�rm��U�v�a���]�f.�ǟ�`ǡ��펷�7ߡ/�o�����Y�i�t��@��t�V1S��� DQ �k�n���Uk֚DD���+:==��'Nht�"���1�yR\�:�R!%��D[NL@([|~4	���	a�xB06�'}Dׯ�(#�o|���������o}S�<������X鋟����|��w� c����=Af��0 �7@P'_9�d���⒢����\���e�\��.�F�|�3:p┊�fx�i�Yb��L�<�C�a#����ԕ��1�v����͟Ս7^o�ڽ?��|�<��d��,���j�Z7�Ӱ�zd7��~��5���0ivw��ؘ��}�!=�-�{������G�z�
��ͷ�/?�	]��<}���{�Y�ݻG�g����Ȗ�4Wm�P['Wk������@��{�C�"5=�J��z�F��Kt�;ީ�ZK?��>��/���)e�GlJ����P\k<7�iC7����1l_za�����v�|�cҖ�[��/|�l�K�y���:p���:�X2$�׬B�������\�48sAB�\��c'��s����;��z�n������������с/������ȧ�fbD�=��Nς�X�`*��\V�_s����-4���1p��z�gu�V�Mo���ц�.Qax�7�3���^سǀK�5���'����EϪZ�~����jP_~q��<�+��]wi|`H?���z�-�j���_����;�������}��t���̔�A��}RxV]��С��ɳ��И��1�*���7\��_[).$���GS�JKU����=j�ǃ%�p�����]�.��<��]~���x�3�^(J/9�TF�&1��}i��d,��@u�����J��1�?���i�鑚�Yqqa������z�a\�C���3�	ųF@qA6�=����"�R��2�5�#q�C�نNE��!:ڶ���ҢU�@��X�&_��Җ�B.�� �Fi�gh�2�~�zND�8�3�N�\������N�,Hl�y�@%W�%����������~z�M�U^\� I�N?�v����n:��L�3�<����C=z����:et9�P�p�~�y��Yp��dFD�L̱�G-i	���Ϭ���!\�{a��Pho����1�ך���bH�V�]�=�_Mꡨl�1ѨV]a�u�0���\ ��u����_���GGL �p��|@��r�n}������v�|ޅ��Ƞ^��48�g��UW]e݂�/U>�׮�vi��M��;��K{���1�x��U���ku������}WO�ܩ�R��Й��/ܗ��8��l�A�Ĝhw��!������L�f%��S	�M��ѩ3�b��#��u�
�.�@E��i������#�����~���Y9���~����oi`hȜn���?�>~�G���{wk���������x�|�=���+�4�R�Y觐���M[�̵���r긊�N�-����:����\/�;`�`/VP���5�2I�'�x~�6 �81 �����i kA��ȉ#Z�n�Z��V���?ʕ	ډ+���v���B�,y��x-��օ/��JD�����?�}Q]z����O~�+.�T/������m�������ܾM���}=�Ѓ��..��|��P�dB�x\7_s�F�=Z>uF󧦤HC�VU�fE/MS#�W�ʕZ�v��z�oj��m��'>�G�١��E͕kj���r�#E��(;��_�-�V�<��fqYÅ^�.��+�a?�bŤ�Kz��]��cx�:-Ԛ*�X;�5l=
�$�v�#dάG��2��,6���v�Dh�~���M'�T���������k����c��7���6�^�����瞵�#؜H�����L��m6Փ&��Lݣ)��7m��k��+s���Ϳ���	;��/|�oL+-�.�[�v꾆��OOO'�����ܮ5U:;�����-6j�Ν��K�~�����nf�]���E��e{�^]Z(zʄ`Xw�n�7��Cn�`��F��F'�/���˻n���/[3|�M3�������pӣ�_�\+�^W.֜�%� �P�(\���^r���ht��&/��B�zu�N
�t� "�����܌_I+�ꇑ���c��پ��I��9���Z�ұP@����F�Y,�]uos>�Qsz������/�y�	!�d*���N�W���N�&+���Q���B��#�F�R��=;��HZ��-3��j��_!�=l5;�]#Ϗw�el�=UP���e7&�l�Y�9�0� ��OŃ4.�h��z�ra�P�(���ј>u��+�N���>�񩓧Փ���' ����N���h݆-���'�aV:b�E�Ie3����֖�XA�B�ϕ1cJ�k�T�m3�8��Z�E���K��vq��|�NP�P��)�����O�:���5�,��9B�:"ו�c6_��-8���U-���J9x���yˡ�eP)�5�;�=��iI[��KEN:Z��c&&W�壇u��i�bz�N6�G�bvP�T���oc�i`!����$��&R�(�-�\���8����b�G��?.xB��@k���]��E�Yr�ĄBg��1.�Z�b6s3���VD�e��(�Vq����o}�;etϙa�388d��#G�{�r�[���[t���zO��7k������sgT!�fҺ�o���
=�ȓ:~bʨ�V;j�(V�\b��ړ>`s &��@�\�1e�u!P��)�+�u��jE�i�q��Z�|��=0��=y�z�kǏ�R��J(�1��nڴI�_~���D������*�<�:yT�����ګu�W���~_�y�{�ן��?~�Q��<����>mZ9�L[VΌF[�Y�Uz����*'RZ�~�r}�����Лn�S�����{�\k�Tk*��%�c4�Ų�v�iG=h�L�j5����Q+��X��Ԍ�Ku��i��N��z�XDY�X=���am��L����6,*��Joiv� bk�xo}˝f����wiy�M�w��M=��c�B�>~ؾ�FM���M���˞m�u�%W����R�b��r����׬�y�_�}'�뚛n�tvq��?��0��Z��W�&
WrN�_��))���o
0�Y�r�R=9�����������invi!�4'��v����c�IeĎ"f�*�EӠϦz3��5���u�����N���;?z�#�^�\#�Y[���$a�(U	�0V��Ԯ��kp\7 u�]���tnz�i��\��M[+�|�H�$x��r�`���X(�F.�LB���'&0;!ƓV�*���бߵrՙi��2x�$ul���$p@_�WP�����`�qӟ�����Zu�,�'/�	���σ�#�����>�r��7oYZ���%�txx��`b�I��7�&�\-��y3�+L788�B�3�/�fM	dl�ߗS:�PqnI�$.u�r���3��{*IF��~���������
W��cNx��gĸ����<B��@e!��s���BW[�_i��Jy�z���q���_�(|O���%ꌃ_=Y�Y���Mk�\:i���gRh��N;��\�ˤ�M��D��8��f3��\�,-�Y���HR��A��Ғ*5w�UԢ
�jU��a��wQ�Z�@�U�����x���k�+=rG�!��&hV����$�}�Jc��P��4*.B*��U�p�cO"w4�{���$t{-�"��4�]0����'L��� (�v��F�RV;�R���,�4x�+'V8��9;�ɕ��s�dsδ�+����D@d`�_��9��e��;�-,+K)��>�f9_����6�Kx|��t3Ʀ
c�bD�F�Џ]���3�tf�zs��I�4�XT6��D|�:���9a��vm�ZIk�k<K�hL�E�2����������V����&ƴeդ���/�ƛ^o�VX���O;�������^�TZ;�{֚K��W���i���r��+��V+'תpL���/��g޶ҕ��!��ҼPoA���4ծ6=��ݕ�@�0�v�e"4;=o��v4�����d��z�l�R=��e��q�H�	���!.z�V[�3j�.����{LRJŢפh����a+r�Ӫ��tۭo�����W_6cJpO.mUɹ�3*��m�fڽ���4X��E5�R�7�E���.��*���R���G>|���UO q��!1��4<�E�mm�q�;�+b6з:ĸ�F;`P�'������53��d6��hi�Z-`�j���!�{�a�jNOΜбRuB/�������o�m>�ku������]?�LdW5�XT�����bT��F�\V*V���E;P�bW\*Y:��B�'��x/�C�8�˽C�O���aپ�(��n���X�jZM#�}*d�*�M�=���C,fԖҙkE7[P�!)i���ғ$hy�YW2����J�����/-�+E���ĩT�AM�@��?��n5�v���Ξ���9�Ӑ�D>��)BLQ�>����RAE/��a��qw�y�s�ĉNgB��K���4����<cܶ�2�ܠp���ƶk���xA��_7��{����0�k�� ��U�Ɣ��MYo��τ�%:�r0�`�a:D��g�û�k�{W��L�`Г�p�8�Z$I���g���A9	V���@χ$d�J�x�Y2I�����pɘn�������q�JuED��2!��@�b���R�<��	�8
��2�%�)�NY�pi�+:iVY��T�R{�Ҳ*��b��6�^֏���" ���N�o�����kc�B1Et����-�l��l�)	ۖ��P<��V=g�{�~1��l�}�<��<-A(�↿0Ao�3�J끮�*����+s�9�$Y��Oΰ-U�(Fl������y�fEu~��)]�9p&��O�ծ��%�j`�۬��������\��P �(��is�9�ϜTŷx^�
�WHw����3��=k	�<��b4�V�Y��Ч�((��Y��Ɩ,��[���i�`*���K��l^�\q����_�R�hE�D*�͛7��>;s�]b�IYM����^�5��{�V��Z���4��F�B�eP��&�d+L�"A�)ןwB��>{�%���*o6�*��F�c�곆�x��:�g_����aR .��AW$�r���h�xwƆ7M�2�4� Ī�Y-��j���j�1Qm+I�7��z��QQ�>d�N���}��r��щn~�񔦧Nk�X���#-����<�!~uX"fk�E�F�"���'f,P���A�>��ܢ��&��	ɸ�-��x,�t2�8�ڢg�!�8�Y�жG��XS�Dki�H���r�e��͓'~����y��O�9��f<��m��Z������x���\�h9l�'^*��Z���6�&�w�0��Q��j��d�*��^�����n����ț��Z��P�zq��eͤ�I��E�{��C�H9-O�NgB噌�G <h\��qZ\֞����̬R��N�[g��t~��o�x�����Z!�R>�$b�.qp�	$xZ�-�F��펌���G2eS����E_��1`��wQ.���Ǩ|"������'ب�V]Y ������d"�+�E����\�0?���(��hg�D� ��tlzZs媲CÚ^\��j`x�E�"�R�NTA90�;f�|�X�B�������^��r,ڴ	�58�q���=1
�4"�z+ ��E��%��g�M��:8Y"��l�Ht�
5��AC<�J�����f�O��s�؊E�faT �r���b��N&ѸA��^�&쯾@�N�3Pv+���}�	�u"�ix������պ��W*6��[ӻ�L=��	�Hxu���j�N}�^9�w�����`���l�#��{��7I8�pI��vTlԭ�X+���݆Q*l�Ag3�m��蒉����X�_�aw+u�HF�JǲJ�s��-U[���|�����{�>P���a��]L���b�^v��:8���sG�ǅ�x@��_&v�wA�E�A>��J��ê��.��ɤ�^��@�m��Vrq/z�}Z��S���d�V?|����^�-]�e{�/���91p�`K�Yr~>�
��(�4��*ͅ�N"t�ݩ��@�㬃��HU�d�?$��ꪩ��`�FGG]О96�v��vUQv�񄛮z�� =VLK؝3��p��&�5[���� O�?����r�l�<��p�d�<,"'���<T��{6!5*��/@]�12�w�e[v>D'�K3�QyD��T���o*��YB4��E�k�� G��ܚ�	"�������	�m�y�si��W2�����&Ec*˞��
9�R	�k�|��Ϟ��E���;L����{\"�T4^W_J��Ɔ?����į=r�����[��{诚�̪F5,�٭�q���/�Î�/�� ��
�V��WW�n+t�T�\Ƌ%�t�G��si����ٛ�;wP�� ���\RV�:o�:]p�fmXݯL �:��P��R:a��7���O�Y�*�#�=�=82��~�����~�{zՊ�<1�í�T|p�!:x���T�`��X�jj����U�0�|*	Ϗ�Ex�����^%�DՓ�9 ��x�r�0N�.�9�GH�w�U'��V���C��צ5k�y�*m\;�`JGK�P3��3e0M�5��4��N�kH�;���o���:�ei<�}U��u�n�̻�vht�q�FRJ��hp`�I�t���E\JŅ��X�`�Ze͑��N}L�3z>�_��	�]��*4?���>���H:&�Z9�|�f�v�tN�6�^��+�;�*�0��Z�.`��� ��Ɖ/F�$`�y����v;��G��od$�S
�}��=��"�������p*LV3r�uQ�e�'���'�y�L��g�c�<��.+� �Y�9�g�����wA��ȹ�U��ja:f�09�r|h@j��nǗ��й� e��9��	h`�����Z(��]Pkƣ*R�$�j� ..��J�MYo=�ϪQ^R��Q�t�
��Uh�	-񥯯�σ�Dǵj�ɠ��v�.�;ŧ�	�"09���w4Tl>��5r���̒G�q$� 9[��Ҽ��Z�t14(���E(N��Z�?`Y_�W��G<�S�iK+��d"�SI��x���С`2�w�̭�[V�L�.���ug��{�h#`6�H����m��(�a�|��؉�ot���8�֒p�t�����W-�l5K+�XB�=������,UUo��^�?��S����4?$f0���z��dK��G��k���GH�S>�8��~&�TV�fD}9�b55�H-���!e�Ǵ�Ņ�Ј�I�.,�j#f��dOB�#��a\,���'M.kAŽ�s�
E��n3AcJ�� k
��0r��R�y���=s�oi�'6�ur���r�uu�X��S���7~x���z,�
ak�W�F��%Wڑ&�~mݲ�*SP� �T�5'v�7�RH~r:v�!�lg��ś7c�Ȼ��� �	��/�+;;Z͆z{ԛMi���Z�r��Z$(F4"�E���!�����QS_n����`o@��2��lF{��?���-��wc\,��1��h�R�d�F�݄�e���|�ctvۨM�L����ic��9H��G�t�@���w�p;��:����uPco�D+�=���jE�n?_kV���7\�u���$�Y"c]�`����^��s͎�Ƅ��;`Ҭ_(-7�����_�[ڵ�Z��r�^�R:S�5�c8�yW�۩�@Mz�8��>??���RqW[�L҅F�De�P<�>^�pN4�<: g/�,��f��C0    IDAT���mg�`�=�,��"MEaj䎬��ѳ/dҺ���u��t��5қ�"�'�}���*-���o��t�aM�&�p���9W�y~�~���zn�^t�� 	>�л���;n��P,��ϳ�.�k��t�%�()�=�S������Z���Ḥh�ɼ�xR�L�6��f�T�~6�ݡ�Lw�Ic8����%���J6�R�����&��_���i����#�����#S�g��T�+*�%~&F�����9���ν�Xn+���MQ�hםTu�U�M�V�SV��f�Ng�� /@п3�S^0v%&U�QLS8����@�lu��7d��sc�?�#��ƙL 6�)��{i��F��l:��(��O�yr��媖��hrtܠ�,L�����0&u�3{ЌƄB�fc�V��E�ת�W�T,W\\�&��ʚQ;�b[ip?�䬳�.nM����|X�9(j�݇�]����V�17:.�	�&-���Vhv�y�������=v���+;�M6r��*�(C�a�%���E0�)��I�@<�>&?����&�L��`��Zk�w�B���f��F|�^�D:S�:�(�z;<;���\�h~��x&����
ۡ^�x��.1Ź�"���V�)'�^��?���'/<ޭ�1�aJ�D��4TH�_�z��p�埽rea��j-���r�����W���L#�^٨�}^�Z
��z���՛�q���>*媖KE'w����נ@Ƹ+�+�R�~��K���$>_�X���0��4� ���զ�+ '|���8H��)�\T��*5�f�V�#(��1bK�5��C��q����ei)Tp�O"�@�c��ȩh�?q�;���E2���V���uWߨF��l���yFPܠk�)�A�h@��~F�\ P���žn��m_��j+�qE�2���y������U��q���`��\`�z�\h ��aҒ+�Oh���Z�7��T��*�M����g4�;Xl`=�@���B��N�5N��GhvnJ=��ѮO�5>�Z�֜�nȓp<�w���4u�\l΁�G��P\�y�3G�>ߌ�Q��e�Z�r\׭�$��h8c��Y!�Q2����
F������;M�9F\�hڗ��lM��٣�?��Y���Q�ZƠ��t����I���_my��,_���ME��?:��.����q,C��#����;O E���0��+H�azH�g�t��dT�^�U7^}���?�<u�9e���z��~:J��$Cq̠���?�~Ҳ��/}^���A8zR�M�Z�+0e��9M��Pe��	��n��3��XS����ڛ�U:Ōq>oM�c]|��V��c�v�����D��D0����3'�nՔJ"�$m߼^�_���߬��+�43��\�w{�Sv�m7!$u�y��6#��x�\����hi��#�ծ:p⤊՚���y
Ua�kBV;�R�M�+A&pT�B�&V�����SN���K����(�u�+�U���-rB:�	�A�Ŋ�I��j�s��=C:B5�|��L}ym߸A�Hۀ�2S�c#��Y��/�\�O���w6�S���̔`Z�Ϋ�pX+jo �e����y�bʔd�%?_;�h"g��H2���A%3Lq����3��P,y�ɋ|��{�s	�k�@@ָ��F ��+�¶5������겉B@��������׿wǳG�|�M��UA7L��A�x�����K���g]�w�������3:u� �0�Z�=L�
�o^"��@���(��*F¯2ꧻ
H�0~XC W�R�X&��q`&XS�$B 
����)��@7�b��1�eN�s�EE�)̀Ofl�B�uw�|������Hn$t �*�U��N�<�'�v:�0�`�Ԭ5�e�6���"͜�?7��e�J�i�� +���dRC#����\y&�d�L�K��)��DA+�%`��	gM��÷��l���rE��tw�I�d�t:��#s��X+��BA0n��x��2�̄u݁G�@����5-����M�I
��Q���=���h�h\�}c�X��/���k7��G@�s���ôb�A�fCו�u�E��6ݘ�����X!Fm��W�Z`52��4�$u�,G�@�m���Ixa��!�=m� � OY��Xc�$�N�cY�Ƙ�ǘ1$� ��Q�`���:(�����֑Çl*A��ؽF�5�����70��r��i�qzw=�}j���
�z蜬�P�]N0�b��8TM�.3ɘ�KV�Z1:����Jax���U�ݸ`4���v���h �L6�����<����]����fg�¾�:~zZ�vB�:S����U��nP��-�-6�
[
g�rX�F"�/.'HO�b���E8~���;j�[\j��e��#��@�h?���1
�)�Ru��W�ٙ�ŷ���>�t͕z�[�ä9�0X�E��d�-\D6]!W�tz��:��R-K�(��,i�$��B=��v�t��N���{m7VHF|v�x�<�Ri�O*�9�Z��	���}2c��œ�S`� �1}A�'��G)�T)�]耆����?�9�띜Ac�fm7V�:lVi�XO,LM��o�M�\{�֎�(֨���{�ȸ����in�!��(o�N
w$��Q�];��KKz`�za��g��`Jf{�&�0E��4*�����cRmzA�xD������j��C!FB��:?#�V�	�$���a
�ҝ�ᮄ{�FJ��{.��mb��[���S׎���,������3��D�+*e�*|ӕ���CѺ�K�/h��LOt�l~���ȝ�}��1�|$�x��l���્�+~:uƁ���E�F�*h9�S�A��U$��}�EhP�cl�!c�ɞV��5̡l�h(ۓ��;된��%Q� /
#�͹fO��b�m_�Jg4��KuF1�#��Z�8y�F� ZM����k||�������l������,/Ag�wuv��Q��3�@:���	�.F��/("x>�Ғ�=I����DA�<U����pxy�Ʌg8 
�}	ٍE�HK�e����y��,��Q���ւ�~߻�N�����O*�ـ�
9U+����u��Kڱ�9S��_�J-�q]xѕ��._�N��y5���$�1uح�􆎄����m�����i� ��咘'�8�F(J۾��"v��f�����H'Ҧ'��j��۩����P��%��V�@Р��:!h\,x��p�� �D�#L��@].����zq׎бw�!
h7��MʱV��? VO\�v�z0n�"�j(�˹�(..�=#�hL�eP�ժ�h�7�_��`o@r3�6>��]�t�� �L)Iy�C�~�خ��(�z�J���g���0�$�`Xd�6�&�m٩�Ϗ�bة#Al`>&��$�X](}��}}ށ>�裚���
��g�bz۶m�HFɐ�{e��o��ڇ����2�L�`11A�h�UJ��6�b�=�ۧ�\��F3��zz|&Xg2��$�n��]�^8��jf����K��#�t��I-,/�)����A|_ڊ�"~�1�3�#
k�t�5����ݳ��˄x�i��`~���8�e����q�}:"6F���9GG�D��8��5�8bC\GCT)/iÚ�ھq�~�]wj2+-��5�M�;�5B�ׂ�	�w�Ͷr�Ġfj�R;%����_=�C����i�9��<+�H"iV��%&��
��4�}v�d�0�����ryV������<����x`�0P��V2Tm����I���6���ѩ��_K��hq�������⦵#S�V������-;���d%�^Qa��Z����o7#ںi���љg����yYНN�>(i����]t.c+#�;��kG[�L��C���}���1�*�b�ƕA؀o�Y #����@��\�`Fǖ�x��Qx*)��h��Τ���hM��ۘ�#�qh�rxG�0�jB�����I9r@�j�����Ͽ�T҆M[5>�V�%KY��,��Tq��3g� �W542fkE��FۦX0be�dlM�0"��؝Cqk�S,-./Y��/^ʽ������~�p����+~��9X�̥��`#��A�\^�3sA��Q���DU��-_��]~ ��Eg�:�1{:��SGu��+ЬJ던
�m�r�2���N��6��x����S7m��9�X.���T]�tDD�xڡC���ZS�TU/�:<Z�����Ōh�cCx�\��X��������)��B1@��}D����h�Ր���J�]�K���t �3�3�&J�"h�2���A������}���KO��l���U��9�S��E���}S�St.�/wV.�4D<���e��_�{/�E@@qᄆ$NPu����bi	$��3X\�tB�$���a1K���y������X4c��
�hХ��?��<=�e���2Lnx��>X�0A�I�L���>��U=��c���q���ܤ`H�m���{��qk
D�~��9�����E�(��Ңi��=��LyPDC`��4�|*�u>� Ͱe��z�`|H7�օ1%C��u&�n̚r}j�"����{ݔ�)��h���lXǵToU�xݡ�Htɀo6��������ʝ�J�n04���N=����Uiv���xO!�d.�Ig2�C�5�� �IZ��Q0[p^
rT���c�,�ff��P.k��skU����.vh��{P�Fb����
	M�^P,�R-��R����}A/8��bM��� am`ݫ8��״�0�@��l�Tk&v��Cf���%�3\@w�#磋G���{����\5�^0!�{�T2�?HK��Xi�����r���\�jկ�C�ÿ��]��?�܎L���7z�͂���m��)�Ψ�X��0��e6���,*`��ʤ�Oa�'�t܋�;�nr�R��J� $��`I?��Պ��-'Q3
r���	y�#�H\A�^).{w�Tkhxl�t#�;E��R+'� (iz���0��
ϣR\�T`IY���l��@�ة{��6t��a{�:|�\�������\��{s)�u�͠j5�&�[�T֝b8���|�/���Ɲ�g=���5'!�4௳G#�x:�c�6���x*� �"P{J���k�}yDU��T�����nS9W���n��.��w�z �0	�?T� �����(�"�����޴�y�1͜>e�։t���Ƶ��M�L"����e�촅}L��޽�."�öڤ�$�\�P����Uݡ&t��Ǯ$x~��r2�F����E�(s�����+z&��{k�5yƞU&Q����,��#x��0*a��Hkq~�@+��
~ #	P�R��qf��ђM-p����� ��'ۯ��q�Z������][�
kꁶF%�(��9S�`Z�Jf��a��y#"$i���&�^,f��a��Te�+`Oa@4V.������fc�J �=�21�ٝ���e[�WfҔ����GI�+�&���;�
�ѹ�~?�z���[�.9u���s�L��g"�b�ʵmG�|!WP.�P��;���<�
�(^���H|�>���NBc�1��L�6��N�T@����{ ���Hx���5(�0��P�Ìh�(��Ҙ�s�n:�+�x(�cI�k5�&�O�:��]�\-g�W��He|�FG�ur�zz���r��93�x}�CJ��k|�Z�Y���>�� ����-0�s�e@/eE�
��`Q#�V�)M"n�?�/��#�b�`)MB���Ϟ�ɩ��8XE���x-�R�qv&���ye�;������ !f��(h��r/��L�p��c(��`ʽD2�-��ǻx~^�*b:����A��M���.&��cj�M�Co�?+m�ܛ���7m\y�����՗���g�?V�D��'����g��X��B�mڦz��p�2���A�N��+�͚Zez�d��6�^.>sǯ- Ż��J��؁2
J^4F��I�T�>���^��/)��7
�:<L]:�4���/���v��й����� ��h���M:|=T��ޙ0p�ЙϤb��$�����u��[l��
�*�Ֆ����m����+���[ޡ���}y�[���^}_��4�nb" sh��y�V�:�{�oѣ�׀�����\:c4�����;$i�:è�L�g��9��LR'��#��F 6=iY�(�k͞�M<���ES�̅bɀG�#�]�r��"�Aq�6;^�M�Ui��f�U���Y��������z���]���5�L;b<}zJKs^=�rY���0���g~�O�D���g��5�i�p��#�̄&}�{Z+48����z{{�Q�:P�#���>�K%%r}�Ǹûۚ���6�Q���2�</D[��O^B,	�E,
�>P�ZA���2v��|!L8�h7$u��!|�%�[��-�].W58�B��am�t�.� �Jyy�#f����05�&''�����F�°�;3x��>��� (�|BR0'Z�����	=�h*M�<0I.j���b�	(W(�ʦ�m�����z�����lZ�gN��P"���"�"�����B���"K� �r��)�ɸ��Zo��˳z��*��ڇ�?S3�D:���.��b�j%�x��V���D�=���왟�$���aQ�j��7��:�)]�D�3q�Gu�lIh�ag�A��2�W13R�J�~�덮�נ얛���FI�H�Vej�3j�)F?�p����r�4�^��kOn-�k��SNR��v�xF�V�TE,v������F'V��0
Db(��.
>�ȂP�@q䙍���N���1ϖ;GC�j�O=�d�W(���D֤f�t�{�G�w
8p[�1H��M FL1�9~��#��?��3�;��+H��썽JRx�9���c#]6��m8�j0�2�رc.
��>XX���4;;�^x!���I-����I�lj(]^?�����Wz��K�D���Q�j�o��u�V�Q���T��$�䊕���98&�7��F<��d&�b�
g:�B�\?�d\Y��"�Rh���Z���P��O�/}k��T:�c li��'g��C�_��������򡃖5�NG\cv~A۷o�Q /��wE��&V��K���uld�	�Q ���rM�d��!�'��Q�Ssyɂ��~�=�F�W�:�� )���v����.��jcj���š��[d��8��*�.��Qj �;]�ħH]Ǐ���*fh `�,����&����j��N����j�Y'M~�i��W*���1f���e߾}���_}��?Lrz47����pPK�y�O3�2ɶ�l\��^إo�I��e}�K_ե��dЈQ�u�ɃX�W!��]�;�����'G���)�`Sg4�cL��t�AD�i�{9�fR$,��(��h�?g����J#�GNu��dZ�8iD�����Ӫ�MN�����N��׫�����.=y���S'�nƆG�=:x�������	=�����W���`�:������������K�{���ګ���:��ӊ�M�a��s� `YX������l`$Ӟ�A/���c'�z��t앻�Į;����h}��O'�&�18[����I=�!/C�J�v�(oZD�ӦzK�t��I I褧#M���Nܧ�Ų�\�<�MF��x�KQ����s'�k��]Ъ5�tz��f��)����a-��ilh�b��ٸU����]ȓ���KnVo�Y	SV)##c��,����{���g�ǹ�Z�r���"\`���3�X���d��2��wŝ#�t�8��U���)�]  �4+�<L��v����T3�����܎x
 �ެ�#�N������C��/k��W�3�j�㊥{�e�J$�^Op����}��4.�cnbܧj`Y$bA�k��7l�PL�'wGM��a`a�C�y���`"�E���+�zi4��B��f�V�Z��G������@���ȍ�jtb\'�FD�    IDAT��P �Nk�r����4��$x�n�}�HҢ�I��U�&44<���S�r�����Ǒ��4��,o��­�_��_�C�����{^�Y�X5#q�6��%�Cg;I�^�0v��r�:uJ������=�I2i6=�dW]"�����#T�Xm�����EE���$^�y[6��I����:o��/���Ċ�L�9��iF8׮����������ץ�_���viמ�f�]p�Ez��gu��1݌Wq*e�$���E�ګ�����ƋY=���Y�ZS{^ڧ��l�O�Iŵ�cZ:{\c���|I�lt��lZ�6mW�w�`*.�z����D��g��a'80.������/C���n2�>�.H��ե�Pd���(�A�cV7nR,��c�?i9k����a�AQX7��~�J#�gNM������;��P���ˮ��O>��6:>������:~���
��[�j�K{4}fF�''�fr���>����L\���s���m^�~�mܰYW^u���_�y�\����:}�8��N��@ÝW�^*�+z�t�hZ[��:	�#BB��S���f��L�㣎�\����hݚ	͜���[#aqV;v��R���	Ɏr��J����K5P��SO>��l�.<�~�Yw�8����hǎ�����Z�ݻ��^mۺ�v���Li���V�ۼy�=�O��Ҏ���9^P��s�u��7��﷛�M7�Ng��T�F��{542�R�j�+�n�!��,�Ύ�"����9Ǌ7��	+P�b�\��J����-���T��T�}�F�ǿ�1�T��K)��
�T��sM���@�4�*θ�(���Q��%4�{����L/8$n���e��؄DT�RE�\��m�To,�˷k��=����߯�z���t�
��#��(�M:b�Ͻ���&��0����n��3�5J��}���UN�<��9 !u����1�f���Ȥ �8���i�@�4f�
�C���o'��*��re<�&��Eۚ����ϩ;j?�� 8�n7Cw���₋�x��-�'�<^�O(G1���nتB���>&L�(,�x��i V�fgq]{m��Y;�y�2*/̅�R-�vR�XV۫$���|�V����m�"� &$t�05f���\ß���o@��D09�T+�������%u���ۜ
������'��	n�d�;�׺���w�>��:�
�O�Z��ГѺ���҆�/�v��qÊc� y�y��v;������-}�����d�v��}syCB߾y������0F�耊QRw�@0d\^��$v�٠�6(�e�k:�.���ڂ餫2^U��J��B6����hphL/�?��v�������$��K/֮�3& ��Uk�httX;w��ƍ��:6����oՑ#G�w�^w��^}�v�����'�"7l�e���nW�KE0u-Ͻ���<�H���^�'c�ӑ�E��x�F'-��e'���1��g��;�0�s9h�s����O��5�w��LM?�D\�~�ͪ�漃���t���Ǖ���2�38;}Z�&�t��Ͷɬ-����%>���|�y�>��CA�V�UW]����;tn��F��s�>��e�X֪��u�eW���#ڽ�E�hU��N?�ᾜN>��w����ĳ��r��Z�z�f�.yO�u vd �}�ɋ ȑ�F|A�;��Bw�͏��U�s �;2�`1ZU�Y5��[7�7����x&&W�_�B�ʵ�z�F̓oיf�������q=��cbo	���k��9}��gt�u�ꩧ��VA�:�ַ�M�>��N�<�[n�������gm
=
�ի�j��-ڳ�%�XT'�ҙ�ǵjŰ�cY��g:l;���ç4�z���u��MM�9׍@/E_�eB��ߏ?̒z�+�؀!���68�"hD �%��㨫��ஒ�������,�dzꔖˌ�s^Y)�1�ծ+�hk| �v���Ц��k`x���|ȸ�L:���+�ʡ�j6�ڶ���[֡��Փ+x����Փz��u��)]~���?g�Nx��k���飪�f�q��zu߽���7ݢ��y��Y%�������Y��#�2#T
o&[LT��:tȝ�E]�8�.�Έ������~�A9���l��O�O��s\�z�}b����� lFNw�,�A����iI������L)����8����z�Y�s��l٣��Ii����df0*�U�֫�Z1֯�S�Luf�?�P��BM}��\�d��ZZ\6��&��������2rB�fϭ]4b�ݥ�u
P��� ��; 0&N�4 Rq��Kֆ�]�Ž�0K~���O�ï�*�l���k�A&/�;�?q���]��\��f�1;?#
���<.�6���dz�ڽw���@��0^K�bJE��-�]��_�Co�����˿���3���H�:	�~�Ahr��.�r�z���ג_�������C��t�`ai�㢆p��
_>�μ{�I�f �R�V����#�i��u:u�~T�.�X/�yI;^ܣ���0*v�Ht�UWh��O�� w���.����cOj���n�:=��3��H�Xc��klڰQ�ׯ�/��Pe3"�:e���׽Η���R)��%�M����fOTq�������R�/i��d��_���s�};�8�ݓs� .��e*��G=����b]ei�rQ&�2���.��lZ��K.��� f0�{b�L�o}���X�Kp�V�v1n�������	.628s�:{�P%��j�$Fȉ7�ώ�=�r#c�ZՄ��p2��m�l�|�C��"卓6����\恞2�cţ�N`iy�)�L��E�=���Ɔ0=1�g���>=;���~|��Ǌ<�T����<�_���pN���'ѯ��;[ے .N�S�y��l�N
��5x�,-<F�����|�]��iL�����ŉ���1k)K�͂���������߃��8%�$���ڍ��b.��Ő�P�L���\V���#T����/>G(ҍb݄R����P4t~bC����ސձ;�����/>1���s�X]�A����~�s�A�̜ѽ��7�y��sf������3u�Z�x�8I#tae�Ԯ�c�˥O*�;>���i!	�^ѷZ6�d�K_�	ܘ��ÂrO+��ǂ��'���e��R]K�9T���;�}(�)ctbrlT����I��O�<���*B�J3NJuM����~7Ν�����q�#L�����]<~�W.\@,�����	wrf.O��x�����>L���q�ŋz�'g�z���=d3T
�%�ez��pjb��8��Ý����n._�P�i��?G���DP�H�F�Ln�!�'D?�S3+�G��O;��[y��d�`���s�?��ŭk��!��Q���,Vװsp`Z��i�� ��Ƶk8:��7��ƻ�+�#J�g��tk^]^�����ȸ�/���Y�بi��\������=��I�,��͌�I��-v�P+�������G���7�)��6~G��K�b����A�p5cuc]���Ŷb��@��1��$a��c��<�8�z`��lz���V<��X;,H�1���4�e�d�Cmx��H����~)�/�<f��9�o���9�ŸkgXy]mO�*�$|;��芠\�c�ټ�}Z�2��^�tSa<���\��P���/��b2�u��Øп-�
���詳8I3x�����Sb����G�Y��1S���C���<�[d#ڐ\����'iNBx��QC���X'���P�$���clm��d�#�!�M~��r�ʤ�87=��g�p�HkH����e$��䍏O"��it�V��	����X�O�7��/���K�u�A�a{gO_<׋ew2K����X}�nS]ݤ�H�ۇY���.N]���#J}�����ƥ��A���d��H���5�J���z���v��}�N͐���x_X�|.���V�&Og���l`�ɠ%L	��������b�S��{�E"�966�������~��G*4l@~��baaAr)�Ft��M����5+�:���`y�*�7������W���Y�>�˔
�2�pH�4�A|5K>B�z'�$)t����ʗ�˄o?��m�u�����hR�h����Sc����ß=��a�(�t����%�q��v;��4b^;f�FE�"����!�6�4��y>5=��!M�<T_�|��pn=}�����x�zKO�k~��Lc}m���1?!�ugA�;[�Q�028��]j68<Q�M	
%S�FE���a;m�cWn�Y��!
&�̆��;-kT�y�ZREB�<�h�C[9,~NM�#��8y�t�DM!����-�$�9�����YEGď��|��_hB$�r�λ�:<��˯�����ocwgC�2��⇿��XY����Ο?+t�������x��(._����5$��^�g����=\8;�'��*`���ѯV�zG� z�r"If�Ţ�[>��0�0l��s8�Ε	C:�Z5C�I��n��-[Z���Pww,�k�`ce}]jP��>W�-��ͻ�S����o�@�� �{�1�G|OWV�pt���kW������rh��{�|Ag3��N��9������#��ӧ��۟���'�KG�*�#�1�|�X����ۉH� \��Nw��nMDj|F��O{�P�͆��-�Zoo�~���o���&�������G�����U0��b�D��h(1�9����P�!VKea��ljP����o���ɦ��o�{
E�r�����k￲.r'z���Y��UL��<�*���\+�o��j��^���e��O_���)?��W/�:'��O���\I�������-�N����&��RF%;xNJ��ܭ�E9�m�����~h�4���ً*R+/��N���| �pE��ՀS���8��C��54�f�
���
ֶ�d�J�I%��܌i%���(Cb� �n;A?��VDʢ��B.^Dgg7^/�`[D"C[ʗrrl\�<w3���ƹ����6��#	�%�v����[KO`.����v��c��m�FN�X3�6�����"�\�#Si,�F�ԊmCʭ��wV�ͥo�k,�\U�>�3=5��.?��#؝���6���	�/���Kx�)s�F'�4��ǔeLt�����}�;�!����k��ؠ|��t�.�����1�BN{X~7��-v��{߈���0����rr���e���qz�	u������u��TV�[[:Y2m��Ug*��%�{Ng��k'��2Ku�ʻ������z}ƙ����|zS3t��z9� �N��B��c�V���/?E��D��E�Y>���!:�v�3Diܘ9sF�?��_?0�L`f��-j�W���
�b ]=F��k����� �J�FM+��Yk�g��gP*ftP'Ѵ��7|
]}���eg�Cz{��t_�7�x2�f��oH�F�9J�h:�.�bMӜGV�TV���*�i�ݪ���Cwַ����'2�X��ӹ� 29C;�8>č�gq�����Z�ޓŁ.hl�/��řS�x��c ���i<�{�Ã8N�>���^<���t*)5��Q��}����x4���K�q���f5�Z!+�q�M��X?|�(6".Ur0��"ֆdu1�����S�w$"R���Z�Ri�[����Y��kxI���v��YM��#�`�=�I�(n�\	���٨����H'���<:"a�?�^�|����b�J�u���MO�
-�����۷�s����_�*����7޺�����s�����za�M�V�oo(��	�7���i��n�A�\)!1��񾑱��,�R�}�vD�o7��dn�I$��B�����8`#����#� %�+��q�B�x���\���o�F!5h`vfZ�ܣ����i�z�������K��ӳ3jLH�	�d�B��8�<Z�S=����w�>J9C5P����׉B����j���p����(�5���'�_,���o�:x�H��y�\̬ԝ��w:pv���:r'F���t~T��mE�	=Fg%�G���J�P9�
>7��6�K,�2�ܒ8�q�r	~���n��(��v����`NЀ�Z� ��VSv�0=1/��lf��	ary���,A2/K
��u����<��!�R�HKUB(�1+�\�U�a^/3�	�V������R*�^�!���������{�,2Ŗ�H�0�[�$�,%����T�Zz\iˍ�^�*-�@�W�?z�%�0�sM;�Q�P����=t�����^.���0y�����b6�j���F:L��CWwL2����z�(�yB���;��zoo_ ��P ���a�Ãu��BeJ�QJEC� +J�X|���
ɸ��'�Rӊ+�� Vg@iG$j�d�J�sjjO�d�K]�4?Z
[�W�!��T@!E�3��u�E���X�<�V3�"�bL��鴡imh�?8����s���]9QmrK׸���}v�9=*��H�����Gs�f
��o߾�L��/^�!!A�(���ҊlD�hUE��Ή���+F�&=�SN!��!R�[��Z��\Ewg�'�!�L��G�n�d�wT�X���Ъ�l����̆��fG�Gߏ�<�GN���V��	M� ���j� U��>tvD���E�ؑ�5M�P��Գ�0��kQͣ'�õ�gP����@�i��'��͌��n��t�s����sI�Nrl<lx��[j*�VWtVPC~W/���s�5,±��._<��YD�H�+����4���;C��'�fO���q���=��H�S*�����EI��VL(��v�mPP�sQ����h9���f�Gz�wؑˤ�0+�+�L���<IzY���(�G����.ɣ25L&<~�����5�~�g'x����Q�y����I���b�e�� n�|_=|�cB��4+X}���6\(�xW�@�aF�g�Sg�u^�;~�6W�}^	ml96��r��1���l��0�vke�O;��j�p�[$�3�"ܸ~�r^�qks�=}X�9����u��̗�J�Fǆ��ۃ��~���/�xGGƄ:�d�:�׌����������ʿg1�����T*�X�C$d6^s��Aux�E���X]_QDh����T̲�b�׬�';"���޺��n��<�f��?����������P�M�_�����IA���y��dҹV&�a�t+�<��J�sj�q��g���&#&���o���e��))�jtN4W����nC�l�B�w�H�I��X����s��|�7ܺz�lB/*����(r��N�9�ٯ�l���-;�Hn�� N����khdP/,�uh��Pr�*� �X]���s0Ӡ��C(���Pw�����A�d�;"����m��3ӝ�j+��-�QT EW�A8�NQ�z�u混���!�~���N�˕Q�6�H籵w�kg�$	"نR��LZ�w~�!*��|Q�6ܻW2�4O`C4���آ|9nݺ-	;~�z�d�S�E����X�d��0vU��5�MXL%,?����&
�#�X�D����w>��Tu�=o�^�i�J��ei���Ǭ�������ª���:#��V~��D+>���Y����EP�Q�\4*�ug��'���"��KY�<
ýH�UL���w�p뺍�#�I�C@�{��7o�o��cCcL�R�JV4!� $������0���p$�|���K��`�5l��`��\	fW�����i��ly�;�i^�!RV=Fz�S��/�{{�F3�I�S ���ìz�ȓň�/]�dLزR��唜�B�M+���Rl�ߪ��I�W7�wL��#���
̵�>�X��H�h�Vװ��Ղ}!�1���b�����%`��p�͠�'���Qtv��sPjiu8q��C�����K���8���4�7�yI�z{F��F00y&�9��0�T���~���PCK�[����Z���o@�<A��n��T�1Q:IG���{�^��� :�!��no�bim��ݯ    IDAT�&����}:Mje�j%L���3��>ϝ�}$R�I���zE���g'��DRZ�?�+׮k��I�SW,�ۅ��=�^�E�M$ɐ�"V^=Fr�f	��E�j@�}���nm#,^�g"amΏ�y�s�i�JS(��j��p5#)��<�*��7�I�
C]��0�R(�'��� ��}�i����ڣWEm�Yᮊp$���Aeq����̬P\*�8��z��~N2��_�)����
Q�=sF*u�ŉ^�,�t�� >��]��ˊpԏ�b�˯�Aϖ
pѰ���z����E��ߺ��� .@ѿWA_n6?��?��k���k �Hȝp�lf�
��aǹً*詤A�o?��	[��Ҡ��m9��Ii�AAo(>4��܃v�{����5x��:"!I���L����v����jz�!N�!¦��8=>3��.'��V�wp(x��T_� ��)�c�l����'����'48c�b�������g�Uh,�Nv��9X8M�sG|(Tj(4��p����)���W�p�j��ѵ��q{��!,�0C3��~�/]�� �e�IH�jZP6����J���5���H��p�Ú���̥V�����(�^�vÄ��޻�N�5�MN��7�͒�X�$"ѣ@(����]�)���/����&�
:P�Q�Cj��Xzv��m��D�+���ޅ�Gw���m�� ��mm4�m��6D�.��>�Q#ɩ����g@x~�[;hI�l(��K�bK�e���A�Vݤ�5���� 8�ǂ	d�-N�u�embO/�fv�uHR;��?��Dx�+M4�ɯ>7,a����R(��~�p ���ȍ�?��n���"v�[��RG$Bo�:���Ff�	�k���	��Kr33&�o[[�C����4�D1(��XI6�b�xW��ZSS��9í�Q-)2t���HXS'�>�+���o������@er[qvbPzt*b�=���oT����0}z�A/v67O�=���k�p�ƺ�̀�V�F &ē	��[w9�����G��xt�W@5�2ar:���0u�,n?j��G:�1���gS�i�l4��������n4=�H�`Y���3�����N�4��جp;,���E�'B��g@d�0u�L���H�Nt\�WTЋ�$Fz������\^dAQZ�����Dh�	t����95�����abtB?#��Ã�)�ml!����$ӛZ���`k	�jɣ}�Gl^C�c����`g�Є6z�{/��<5_xc�h��8j���Cw���G�Aə�Z��΁V~y��G��AO4��hX��n������Q�)�|l��=�&=A�:5)t������e6"S�B*Iv�57�r�~�+�;b�����=��'��1�^W��f�Y�*�!_Y,����u#��b�&�ULw��������ܹ��U��6����������k"�.�|@�Z�v^�M=���)��C�(����c�Y��i<��l���w#�F��S5�i(`�R���c�x�v��F������~_8*�P�nF06X�*Ο�D1�@�x��(��N�!-..#��W��px׃�ɓ���iD!o@༙�Pϝ3:0t=�����P��`��}��K��*�Ŧo��}��,����L��f�/@[On/H&a��mAW
�c�>�t"N�x#U�����x��9}��/V�����k��TuH����A?�[���ȕ��0��'�~��Hvq{�o�	~��ߗ����̃����������MK�)��io�YMc��Hn����2���\{v_�BM��f����;�H6F�6&G����=	�:[�RN�l�H�!��`��)o�猝�F	��T8�JX�(�jx0�[{i�LNɮ�-P)��,���Sp[ G���� �z{�w@H�����d��=��I�]i��tx%G��f�I���ŋ��\_^�u�T�f�?c$����֗#��V#��S��C��x"�r6B|�r{wh<o���*B��`!W�-�6̌�k�v��ƨ�=�jW0��)t��yJD�8��b�V�j�p{�� 6����J�4:�N���[��*��G;c��G�HJņ���$r�#�nm��+�����\���&��r��Ш(�9`��9�^Z���1�� �5��Y�n|��_�e��V<�iS$ڇ�1L_��x���T�G&K\����Y�a���M����C穬�������V�;/����T�B�ac���ų��E�(�2BD��"��^E�ʠLvw 0�0�KRV����6��bBV�<�jT��a�f�t��I���_~%q*#r�2���03&�RP���O�x��P
Kmy[�/���1L�rٸ���r��1��^F �+U?�kֶ�n{D&�КxX,��^|N��`v�,,�D˗�=���.Y;^��2��!�t���h6U�;<���M�m�1R��t��a��W#z��r%�w�g0����E�'���������Hk^��ilΉ�q-æ������sUɷ-�:ba��������F:2�Nzf�ݬ�'b�?��ε���� ���������r��*�4�]9�2��^��cu�¹�8ɕ�NQ�mڕ����`����.���c����n��UH[�c�P�c���aGgG�}��'�z�5B3v��n<y�
�/`rz�4;5	��Ts�qi�4������8�I�uQjF]���Y�䄥X���eG�}Y�gj3��13��3�.�u���r	l/ϫ�[�w^�!�#_��7.����5)�I��7�]�D�(����·�}�ߐ	�8��N��(��H��v| ��:���N�����7y��V��^�ӗKh�p�E�#щ*u�7/�G�������G
 Q�i�� ����ǝ�]���k�6�h���j�1����_���^��:�T�ql�|����)�%i�|��:p��mtB�ljި%Zp�b[\���d�q���hIq%����Z�IJC�/;caM�\Ӹ(c��)�=�S+�B��WK��;ʡܴ�Դ���6d���@�딿 #]�v��L�Z�,�nt�t)p�S:�%9E�"��55�w	�m��>Ie��G���;�6_a{�9
�m8�5�[H5�;08y��!0��-�1��F�?d���F��H-#�R����d�(�+[�2D<���q=�R'�I���|�Z�S�@_��p0*v���:v��ȔDB�IiW�^[A����w����I��֖�p��9vw �<BG$�"�)��?��T��d���ƕ�����X_ߔ��iD�R��>�Ń����YԄK����{p��H���N���q ���a�o��:�j9�����g��H�x��u8��}0�
>#,(Z�СSo,�5��Vd��p�������Z�L�2��[]�IvsA7n\>��� N����;��nŭ�7��L%�vۅ�M�����+�,:A���F��"!?FG�t�T@��]��jI���+x���*�����(T�P��f.��чMfê��s� �F,�^��>�P�"�ÜG9�v��Na�s���N"k	A���1�P�3<.�
���!�Z����{�g�P>�1�����a�n��נBga�zz���Xd.����P����,T�ߓ�6#:x�y��3B~u�̣ !��0��+��I�+(��>�5O��&t��F%7���o�}��WA�N���?����~���`��M�p���Muc���q��t���:�6��S�:}+�$��&j�m��_MI���S!J�
xog����|��e���&.�����6�b�+D�Ꮅ���`�;,8��D4�D��ĝ;�����_I�/�D�Ϳ���8���#'�����=�XF�$���A�%Ə4�Z��xObg��1,�"�J�|*��W��!�=c(�����y��(̗F>u��P"�	������O��ѼՊQ5�zC�H}=1���!f��H^�Ϸ�T��bB*S�'���.��^��֚��4,����Z-��M���ɴ�s�ړ�#9��7N9Z;�t������d���N�j�3�@���E� ܃[�U�J	�<���޺�_�-�B�;1u��
z�L�ծnY1�*:��Ŏ��Um#�� R0��A�����+4-���P�&�4��(O�^+������\(W4��?}�̓�Hq������
|�*��4\V��Qf�]@"]��GsrBd1��,�uǴ�#�����jJ"�ag�H+�U��<N���6w���U���߅��%l,�#�����
����w���ju� �I�6��pŽ(&�Q5$����;L�;u�ĬF��F	k�id&������¡�]yV�Q�[,2`Ȏ��KX�9@�p{�*�	�.N6�{��qp|����8fsm׮\��?�E&����G�P�A2�f�\Cd��&0�V��^2�DF�	n�G:	S43z�p��1P)p��Ï��)���ǨX�8�!J>*r��Y�5I�S��2q6Z\�6��N�j#IB&H�bSDo�V*_
���z�jcg��	�����P�ӗ+"�R�Q7��K�즆�xm�����ry��<y�[�{�}���rȳCԍ:�?�G"�����{�驩1����O?j9���O���׆���x|�3X�9���P�YT�G�/"�9���-yY�i׋6��}�8��k��,��7��ƪ�MA��j�+)q�Nm�oG�W�Bn�	�œ4
��5$���Ϥ-*�qйx��� (���$K��G�d�İ���?t�$g�Y|�����֒�{'�)E����H:�[��ܬaa��ڊ�G�!ɷ�bA���߾v�'��X���I����������/�,.��{Y)�����نK���0����8S/}k�N�e�Z@Y���=���m�r�wX���,H�2�Μ©�Q����VʣYe��!3jt���dӤ���.>}��խ�n�z���q�y���`r�^�<�7�D�!)�ӵ?�����Ә����!L��z�V:=u��qloo�`D�	�^��.�E���JUT->\��t��j2�v�����nc�R�Ӛ���y���5���!f1�D�&��Nc��K0'& Z�AD���BJ{u��� ���p�jV�a8��k�`�[+�ij`|�!F��]�=[�;�Ǔ���k����0"�y;�?��ˇ�R6C�c���E�pO+����9�m���f�T����£/��Y��R0��QX����ސ|ܙ���h�vi'�����]ħ���Ҫ�ԅ&$����Ѥc��/�EOw����P"����}�9�ސ�/�AÊO�����l?�sj�2I����c�}�:]r���I����vhJS�D���Q��yuu�>�t��{� W>m��+�X$"�{sO]�O��@�pKϿA1e@�|��v/̞�N_����g�ϒ�z�Z��	#<GM�M�J2Hnt��N�j"�j��g����p @ii,*�t$��mG�ZD�����lV�W,�g/_��W(��+�˫�^���Zc�1D�=���\�����N�%�v�pz|D6�$I�����jZ���C"��A�L"5Q�χ���*ܡ����B�.�0k�7�������fs#[m�G!s�9Y��}WK��8�z
��k���ӍU��G��D=Hh6�bH�y�v:�y���<p�V�A�q�&3%|3���
53�N��C�_O#�ވ_z1���rkkW��뻇H�9c_��ę�@d�ɜ�=�����V�X8D#~<�H�b��C��j�(߃��O���'p5H.ʅ�=@R��E�{G`uzu_h�Ky{���1o��:�x���F3ujգ0�7��<�l��bԛkU8��MD�X�w$��\��U]�(&���뤧��}]���b��Ǐ%��{984���^�˭�ߋg��{����t����!��w~�w�'"�����a�����c��_|�P��ɉ��VA�8-p�+���ȟ������
��q����O��D���e��Qo2ЀTגA�P�-�4Yq��UďNT��v�<�f't�ktIoZ�����"�8+q̝%LF1bQo�$��95�<侮��m��[b�nolJ�p��#d�V���1�_��D�U�d�O8��L���{[��r��N��%ϒ�r,����SII���a�-_�tV)#��z�2:���\��8{���u�,�KZ���a�Z~$�;Iq���A/r��
���~�@簠2�����"E42�x;C^Ik�lAu����R�LJ���:���`j|Dp'�����eӂ!�=�G����	�QA��V����s8}!Л��
N�ǭi���n�Q�#~��t"	ꓳ$����S�%�'f*Y����2�mլ�L��E����C��K�_�;�)�@ H���^<�����e5U�p̾(����'����++��}[���m����Fa�r5d�2� �C�Q���N�ܺ�:h�I����6R�$�v�Ս�C��$��c�0��Q�h�(���a��9��%��px���~�SS���W��Zu��K�ˊۥ�͚D�kyNsb��I�9�_|��B_D>u���^y���⛂N�#�7���k*�ټ1q{�����vtg䯱a�)���/�ր�A�\C
�w",��J��	���	�|���N`1�9"YT)����]M��VQ�It|o��F��/#�j��=7+�]����3,,,� vF�pXMRt� Wn�p��0�ץ�Μj��R�Z���ԉ��I��ww��>y����?�����g�:��0s�-M6�F�9Qb^�!�Qa�8�ƛ�{����p�%ɘY6T���&\v�B�������d�K�ר��>I>�z4ة6lx���OJ�U7,��6��{bn�Ѭ�3��eA8闞������@_�SL�YD y���'�0*�
���f9��lM���� �d�!��%�],>{���n�E�c���k#�/ �?�'����Y�˾M��&S/�^l6ݓ慠�\j:oA�$g�X�"=����R)��C����:�&	�M���71�����bd�(��W�(s�n5���J�{��RFc�#�
6"��$9�V��ښ�¬w<�E���j��P���9���$�EH(�ō+��/?ǹ3��e�=E�aS�*-�]�jn�#�g�y�������r�l'��'�����x���B�io��O��^a:NUD3J*�&.���㣌��$�]%���b��+_t%�٨�����"�-��5��f��9U�0��sB����i�.^�x�ˎݭmA�$԰�������W�����wQiZS�=9b�B^�ۧF�������M��%�Xxax���ɂ}|��Wų�2|wm�r�"b]�Ȥ�j���h�x�^^����R�j��������cXWNJ5ԬA\��t�\3:xZ��g�_�@�+�z>0��ǲm�9<���e��i@O���C�:���HÜbBx�C��)�385:��It�(�tqm�_.�ğ��� #S\�=�b��-���Ȱ�V�d
[�8��jw�̹�`R��X���|�D�ޔ�MM�����0#�̉O>06�GO���Ҧ:e�Z!��g_�`����a���������ac����M*=T>.�55��tKZf�*�)��aj�"$Ǳ���P620��0�w��8<�}&�9�����h8*ȑ(��_=۸�4�i^
�g��u��B�33��]�5YY���|dl���?<D0RJKVt���.c``H��SD����1)����+i�Yc,�*v7_c{�
�-!"��O�O�{�k'E�#��B6���ioe&p�]�I��<���U7�;��@9���w�ܣ*���Usg99<�Y6�N{kL�7Y�%A��)��**�@��/W��f�q��?�LM��M\����i�Nrkw=�8���=�Oʈ��ݡ5�]֯�p�\ٓ�.���`�,�Nn�u�^I�������^>�B��M�ݫ����/�zO��}�Q�&ţ���)cTEV%�]�}t�4����Wk�Z	f�A\�y�g�Ҩ���k��Q��_�&    IDATI!�F�Q�ʜ���Q�CB�;×��c� ���T7��J�X����+������0�	Y<�nl�N��@(�H���Pѹ�О�m~:"ď�z��~8�G�c8�x]f��������(�T�������IL���h�`w�B�`���Q����N�n��9��|"(TR(���d�Y�sOĭn��#C�8����D�j��XS����
�3Z1V�f�&0z��*[�֌tcrlX��|�J;{He���Z�%�7�$�>�U��p����� ج�a3OVg��F�T�i�?6܇gO�p��5��n��Nj6�֥NTrc��?�����{��|�����?��?J��NN�M|�aiJ�)��Z�o������e� �f�'��DQ�Yl�����Y��D��i�6�S�g$ǵW��N���t��vv77T�y�x3B��L*F{{u�,�`s��^)$Cv��"?����835�ŗ��G�d+�Q�����[q�}�M���o���Hܛ�؀�(�O�<.7r�v�,~yjN'(RnF�W)����Xy�͛�N�/S���_��C�{�QP�D�4MݰY�arrL��g�qNLL!�����:<n��{��0[�Ʉ�:�<ҩcَ�r�I�@o�֦�`#'�l6wt8Ǔ0[9Ҝ�*�po�:��(�?ҟC��/>�%�GG���/�&��WVp��)|��H&�111���>�y4
B�ꨰ��a��q!H��BO��9��_���N�	���@.�z_��\<h���D����Nܾy�s��H���/��X�å�4��*�2�M�}�.}�r>'�7:LQ�C�@�G�C~5Zl��n�dO'�:>����;Ϊ�$�>x�ޯ]� x�_/`sc?�������������:{��KS�[�o�/~�Dt���O
�g��S4�����Hf+����Y_����(�w4!�9�,�����F�+��Q�hG�V�f���y;�3FrVX�ܒ̑O�i�if��;��cmQS$�,O�ZWϞŵKcHy켞��!��X�Z��Ԥ���7�gO_��Z�M*Z�桭z	a��?�Wq�H�rj.��*�� zz;�7����Y��\��.d2I��u���4�[g���0^��� n��qՒ:�Ƴ{�����T&��(�]�S�|�=9��T���dC��Y�c�T�I��3W$u�Vc��BB�,b�|"O�T��k�1��-�N����{�JE|��)B� fOO����	�Ͽ���1�\��H�2��%�͌߿#d���s�l�ɩ��<!g�ݝ:g��D�$�1��LA��D��A����h=����de\e�����s_�Vˋ�FH6S�<{��A��k�hq��5�ό!�������0섵�hG�j`a�J�u�6`|lAbѐ�����T)Tx	�Aqx�X���Qd�=ձ���ۚ��LjL�?N�L�����!^�\V�Zw�	�ԗ��>ӛ}usK�4�?�x�l��p`%і������0���ˍH�#�⽝5LN�a}{_�ϣ��j���2
�hg�w�����~��|��3~��{Ɂ�/��?J�,�Y��^G�\n:�����t���q�mlo+ŉ�S!3g��×l���|^$���\�i�/?�B������p7�\,��P-����uw���Ȉf��Λ��#Oܢ&�rx����K�����$��<��%�uubj|LG�\Ѥ0s�,6������]$u��v�1 (;��o�	�q�����_
��e�(�s�Q�A�	"�������R,�R�j_�-:z�k5E�4�j�`�:B�|�v67$'ʥs853+����}�\tS|jK�.Χ�ul��	�09QLͲ�űh�&Lf����Lн�oЍ_~>���-4,F!E�y������gd���G�-f���<y�����r��	2y(�Hϛ7�+j6��ޥC�r/8�?��]0S�cj��Bo�B�Le<���8�y���]��UA�p�ք�h�S�TA�\�a8:<���ט����:�{E�{�`�j�� :P�+�Ӭ��K��U�	�du+���c�Q`���m�I�8����u$�e��"ƽ7ݬ���5�������	F���O^�u������JgU����{߿�@��؄��>�n�(�zxxP���D�zSh=�����^��)�Ն�MAt�	)B�,aN���5I<^�v���CHݽ}����;��%W��	�t���m2������V����v�LJ��L<��\
�Q����gc�p���zM�B�\�0%ӫ�밡3��@4���O��������~u�/^��p?�����E��U,x4���qLL����0[X�ZY��IԐ�2����9�!�w�U�Qɡ�M�����	�"�,��R^+�!L�)x��V*R)��=���w��XM�.z��,�G�Ь5������]�I��쉞�����yvx#���<vR�1~�F�q�~�33=:�l��t\���`�D����TZg
��G__��k+�D�J��F6WF_��X�l�N2)8f�VI�z���c�p�r[���Ϙ.Y���I���w��RAw���1C�'>�9-±�I6ID�ZkZCn�d8���t�h�f
4�!?�_�'��GY�Ӓ�����(�.Vk�犘{���L#=�(����_M�c旧3y�l�!��K�ʡ�|���	�y���upo��o���m��I�L
=���jyI��d�߸z	����1���b"Zj5�3O������n����*蟬�����?ʔm�Yn�V(���{�bIp��������i�8	���t8�H̤��̞����Y��<����݇FN:=8L�eF�.�b�R��*��f��,��p�oV	����"��7J%�F�9:D:_���!��&
ƶ�?:Ӟ^O+\$�x�}�8��%���<4:f�p�������+Pۮ��nss?�+W��Hf�����,S��Yl�����DTRW(A�&!�ț�΀ �78�z�.�����z}u�ߺ�J��WK����GOp"箆Lsdq���v�(脟:B~�QD�^��,u#��)��"lT�X��Q����/��U,U5��P!O ���#����vbc}��]��O���#���f��ʕ�XZZ�ÇE~!�<(Ǜ�Ot��z��SI��'x���ٍ�I	�:��v�}���tA���~�ƻ����	=���K8�V�h�{�92҅O>��}m8ó�%��>�u�T���A�%�a&s�N�cx�_�44����C����[�Q@i##"�j4�N�(\�PY���Uw,��fOO��Wb��������C_?fϝ�*=��b�]8�?Դ©��KȧsX^\[w�LUmT�����{p{}t��Y���6��jBwFS�^�� �N:��n�bȣ���u��U�sY��x�^�r+k�^B V4%Y���R�G'2�lH.�[AC�Z1�g���K!����V �[$�U�&y��x��B�^�6���o�d���(�zz��F��/?��ߺ-���7p��Y�����@�X��sx���|aQ�I��q����6��+�*�� J��X�5>�E��(���z�K3�h���_��.�{��e{�$W�Ȝ쓉�Yh�IR-W"n�_��_��ɴ�ʂ�ZX��l�$�+'����ֺr�ˆ|&-�$WV�O��ĔY�ۯ����@�6�M�B	m0����^�	4+���w��Ɠ|������X
����sp!ʳf����]���(
�"hRxa��������%]eA��p��S���S�LجN)��Gf�Cu����,x�hGe��ߣB�9IKN�v���e�Z���`�s�s�6�u]+B�t�d�,�r)/ΤӲ��ŊgK���@M}<�*|o9��������p� ;{�*�̹h���a���7X���j,��J��皐;W���6ӵ�AEY�Y�H�K�:�٠�tE��A6s���l2��3��Ŧ��,����Ox��~0:����v}��7��dʶ�0�t����kR�nG�Dou�m��G��Vq����Ӏ���j��u(������Y/�Oh�&;�N�o?�2�	�p���G������=v�bLg������>�JK����(��y<�.���V�ɡ,��1'0B��˒���^Y[�~��U8j���K�����KO���o������k�q���T"��3������=�R*�7P��ϱ���tZ�`$�"�bO���<A:'�����'cth�?�ѻȤr*��1�ۛ��¢�!Xp���|�gH5D_�~����$����[)�I���A�v��s�ml`� �?$X����ӯ��{q;6sdb2ئ+V@!<�!��O*����˗�h���?�5��ۉ��ettD��88�ë�/��[�T�c�`S�Ӹ����S��9�׊)<��78�}P�dsrw{5���A��b�M�J����҅s2��~�+�ׅ�E����B;P��}b�
�3s#ZSAw�=�N#H��pP�;U�<��%ە�d�^G*[�Sw�f����� �q�I���Y)���pjj�|��Ϝ�A"���#̞%��)�+���_-b��,��{�����u���+tuu�����_��ܼ}���KyBWj<܀��o
:�ڄ���
:��Z�y1����S�j����\pZ���pO��l맹o�G<E,S�[FO(�ӉSc�B�(S_�ʩ�)�}#��iI&�7���GI��63��J (�֥+��Y|�e�*v�vd,C���c��C$���!�?|�?���"�:eR	5)����D��;a��i�����^����ͪ�jrr�t�}��{Jp���a��!�un;L���{}~�b��
��s�Ɣ�M���.�k����3 _3z;����e�������y3������m�I�T�ȳ��^`zb#�]*l\{1����K���o����������5���ܹ��?�TH,Ld|�E�����Y���0R���	)A��'����
���PA������:����7rQ��R�{P*3���Ӯ�mz��6�m���s{n4U�P:7�׋��fp�b��	�2�֗q�N!�g�w)���i�:N���{5-�!7���:}K^��Gow��26h�b�_-���v�(�͕066!���E�1�?������=Z�l��<S~����V�D��F:<����&r�4B�1�Hr��(��F%?��?�}�'l�G!w����'U���;7.cvp��	��=8�(���}��8Je�eL}�_�}��,&�����B�����<����-��w���9E�k���S�ܵ�;ܓ�	w�4�WG͂�4�AG�4v��K���$���s�O!���1�ۋ��Y���}�h^�><i���Nh��-���ݼyS7�/��/E�D����~�?���*����C�fq�Q�b���_}�*�R�2�� �<@�ݚ�}���?���|0YX�����eG$ܡÞ�h�|��&N�ǯn��]�	����ō*.�N+���4�=�d���Pk���4�{��a<#��?�'�O�@��?����:#a]s�W���L���K�R��="�ϟbbl3�O���'b�߾}s��`sw����	�66���2�.?"��]���q�����[�1xB}*�VW��4��`g6�pr�F� �'���6<:��T
K�[���N�R�ڤ?<��RV�L.�Ya �]ݨ�xx���
gϟ$΂NB���;ҹ�-,� �A���bR-ᴙ%�t�Lx2w�C����g�hpjfZlޯ����s87{F��=$��o���ҿ�������=ّ޽���z�<x�L��������'"ŕi,C�B�&����	��$9$NƢ�s�-��q�����OEpd�9v�[:�J���#�É�ZA������۰�#V;��[N7�ֺ�#/U�l�d�BSn� _.	A�}pS>�#����R�Hbѯ�*(�s�|���\��aX�nēY+q��$��6���������Q�?}��xR������"���RV�h��*�n��b�j	��q��1�ҋ�T�.��z�d���k�� O��V���L�^�YP19t#<=9*�1%j|���Q�`��>�/a'���QB9�l��J�<C�:;���vj핈�01u
_߽�0���~ĺ��f!�T���Ww����{�b�I%a5����Zaqe�| ��U��r��K4ƄNz�l���9�>�`l �O�FG�UM]���!S�%���4<�>���=�GLwRڹb$4O�X�nѐO��J"<�b^��H0��?�u���X�/ ׿O���t���60�GU��8-�rv��K���X ��Gs��?�T��pKKK�˥���5����e�����h��� ��b�RS�U�����X^Z@6��'��~��M�(8��m��+��X���;����*�ml�������&��Tʢ��� ���µz�W^6�!S0���p�`���b̃,u|(���Ex�It�<�<Xd��%��m�p1Y�dU����/�x���5��N��Դ��c�.�GjM��Bt�{��X01�%����u� �_����U�/-� ����c{����/02>�ٙ32����S�:<҇��,�z-صk�����T��=�K126�gx��J]9w���v��p}��#zl��I�lktw�Wf,���HҲ��(�2*0�<ٕS�19u�\K���~��n�}�@"Yѷ�{_g�ݹ����_}����cr|B�:p�rx�j����[;0�]2�ZF6������Y�-�V�E�hhlP��/�&OM�Z<y�T�ɛo�FoW_|� O��[71:<�'�s�d���<�^�ϝ���.��P����Q:9)�xI�/'ttB���(*&���D%�Ģ+^&q$����B��Z^������r�Q��������)��V��7�\�@O7�w6q﫯Ő~��;��ٌ�lǢ��T����s�?J�\�F�Xk��ŏ02ث��=�(�,�q�-�����]5�.�G�#�B�A�4�I�'�&q���'���/�����3�<7�{+眫���sLCr��5��׀���k�ba��M��d�I����3�G��M6;�ʹ+�U�n�a����f�F�����]]���{��9�	?�/N��c�;���ʪ�����][�������^�н����+;t�y�p�ƕ]���N%�U�;l����^
���s����I�K��"6Ni&��������(������v6R��i�k"��H�cb���ݐ
!)h�i6����hO��n5�O_����ު*���������6w_��g�&��������bzz�xwn����.���p��;Xz���N���doS�>G&TA�
)o�k��N$�DX"��TL���9ׯ�G!�BSC=�ff��JajnA�*�fY �w!�>�.JB)���r���j^r��[jq� ��*��
��l���4G��@���6/�ԏ���[U��I���P�´���Z���S����+���$��
G�@/�g2rѣ̍�����
�b!�h"�3����� ��f�c��= 6��E���×�5|N���{KQ,P��k��:���-'F��D���4������w$��㶩c/�v��PDR"�d"*u
�	\N���d�����U�������1���ՠ���:�j��)�����ń�������_u&��5,��ɧ�1�4���k^zoY���a��+AĐߣ���)�������>=B8z��s��C�XZ2v�<6<�tr���O~t�������?��_��ɼ�Â�l�Q�����$�|�Ｋ���$�G�a�8��pJ�J���"���cQΥ3���|��;Ex99��]�G�1[�݂~~tg�z�����o�=T�c�;��|�����W����u���1�UU�&\��u�Y�" ��=X]^�A"ᇇ���<0���~��g��+���4�    IDAT���x���r�OD135��s|�<�v0�������*�ౕ0��Sm�#yt����N[P�˷?���JM,e�'}��
AaW���"p�����<��#���xe:gQ�킞��!�bMFN���=�q\�zE�JB~o@lOB�����;O����ɋ�E���h*����'�������� �#Oh���֩NILOO��;4��O�u�o]��6�V��{�������!y.f(�#�����n2e�@�ޚ�7�+��F`!gbu��l��Lv��z��������J�U��f1�Hf�ߥ��K�gE��3�jŰ�܄E-����`Ƶ ;@ĿɊ�|�5�N�zv<7����BWL���Q����f%3�$I�ɲWت��w8$Q�C �>���ˊ
�pk}�.]��e�����q�8���2�Qf��X�:A�u�b��]�)�#ɩ��?���eH�iG����ו���	!m���հ��������L�![�
�X]�����z��ө��dc��Y&2l�������P��u�9�e͂��1�Z�0ε��g�ξ���+^LϪ�p~\S���4�;:��7�̓Ͽ��h��-=;����Oq��E��>�y�׮�����)��zl
�x�9r�X�4���r�p����`��)D\:�$����Ѣ����[����z������&� ���V></*H\/�s�qO�y:�W/���U![��c$����N��~�c	�H�:<�#&Y����	��Zi��X�x�D�@�LRc
�����PH�|�����F9)߾����/?���P�Ǐ�օt�����7/e�M���c���K��Y�\cY8���=r�C�*蜌Y�I�%��w���ƕK�������!�}i�Z�܈ť�O���:���h^�Pϝ�(�������cQ�}��J���s�����`7���AH�.����w��a�T��\2ִ&#�5PU�p2�4}��a�Ьk��C��Q5�ˣ������ۘ�|�H�w��R	"
a�$��R�1���(����x���S<��PA/�m�	�
��@c�O~�Υ�nw��?
��bq��?����0]���}�)�@�`~�cW�i�͎�h@0R�'4�1|Д�PBD���#WY�H.#s��h��K*L�{�q=�JS:�z&�R��t�7�Q [��_�DJ�����M�7���d�p�F�i�ڱK�!ӝ6�t9�>����Vfr�Ғ�:]�H�/o�	�V��c��В����Õ/�q��S_�l�#���So-">��L'��5���.\���A���)��)x�έ����R1�s�?����o�P��	p��I�21h*Qɩ�����av#:����@v�5U~czq	�@��T�5����s���&��Lr#�
`�˲�Aș�(�\�s�A'͊Ia/*����.���`F����uM�88	�4A���7�Ӆ�
z�t�|\d�����]��	��#�.2#���P�s��e�2v���H��Hf�*��*���fGF����evs����|Z��h�ˉ�N}��Ҋ2�Y|[��j��>#M�r�bY�z�삇J�bQ�����*�p|A���C ����w9����P��J�u�Me����(哂��g���
�a5�2%���n�_��Ӥ�!�%�K���f��"~N�tJ���Ȱ���xz��2�u�� ��i�K�j�Pq��>:�[����}.��ڵ+h�jC�1�\�х����X\^��W�(�V�2ÄR�'���,�2:�T,*Ҡ+����s(X,������ݼ~	3ӓX_]�����1��h���=�r�<�.���$��l0���ڜn��iʳ�������O�T�ɶ.���;{I�<9���oa�S%w��tB��|�b�>�� :<�">1��ÍD.��ɦ;B��%oEX��i5���w��[���7��q��M���A��L")���h˛;��>��@,]�O�e�ݝ��l���O�B�{�]�7��Ž	,�^��ظ�6C���i�ȳ���DbQܸqC�ﳧ���M�x���:���������,jB_�|���gȄ�a'��bS���u��j�N�QA�T�\Yȣ��	Ã��Y%W����O��>w�Ltq��%��9ڦ�[�Jh?��ނ˗.h�N 	�l�Yę��»��&���'�.?�4�����P p�A-�Ho��6���������l���x��K��5�,-ʞ����WU#޹{G� WvmJ$a���Q�\�7��ϴ�L\>���X\_��gO�g e�$�M�������;����C������/~�G�����L�p��zjj59�U�ʏ��r	�܏iB�v��w
d�߾~'�CI�����)����V�S{������9��v?�,��;���f�j��4���X2|���/
�t�^IJv����v�ʸ�N�9}X���[�_ePC�*��,�2"�����T|�y�y�a FL,?ĺ�j���ʬ��(�52Y-d��CX�����;i��������+]!2'��ouw���R�}�	F|�rR��ki]j��r@d1)7S1��C��Դσ��!OV��%��V"�KƂ��A�OdMˉ��/�gT��N��W.�������5MX�`^0CF�2p�DI���k��z��(���i����ew����L
��
��/�3��M
	��No˛��:�@�0�d�;�SNt�-�����f2\C�P/^N���Y��G��i�v���1�=?��{�Ӝ�^�����)���	��-VOB��4 [4ɇ�P*��4��|j������X[5R-V���d;J2N����]լҜ�t����U���v��/�=�i4"���J<)�L헏�@>~ s呛l�������F:W��U��T,���*4�V���@�Y�]=ݸx�~����t��O����ޛ�q�Ʊ���p_�{�T���V��rBgq�EMD���(<��2��KRo�d�[����QH%�L��#/�`��2i����� ���P9?{�	&����f<��p�ꪑN����������i$�L�S�.�Y:Iq��]�ǰ�������]��E�x�<�R^���a��T_��2J��hO^M�dw���h6<h��xNB�n��̺����{w��P�w���_��qH�I�)�޴*�L��v<~5�əet��ZC�yo�����>�j����@$����*zŅ�����C^D(��000�ё32D������3#��jn�xRrp�������<����\�hJCd��{���VA��Ȝrq6(��U�{�������~��.� �b����B.��&B���d���fѶ��o�Q�\i�)�eSL�ۍ�8O���J�t�D��i9���Y�T}ܹsG�<��<��#Ix$O����nЇ���G�028��sc�|5���u����Q��_�g�s	�?~>!�;ya~����y�3�#Hr�:9�����Y�:�꯯�O�ܹ��SA�����?����GES�.���2^7�j|dM�:�D(����	#�5d�e2Y&�γ���\�������x���5t�l��索�O��I�	Mύ���]g}�'G�\&/��ťyu�L����E��yF�҆�,�ʧ�p;m"�0˗N=d��!T�b�T�J�E��g'��Η]f���J�5Z�~��޽{X�؁��Qv���=UJ�RA�\@6r�����fԴb��{(٫au�������� �a7��{��� �[D��kh����7�$���{�ppӀH�i�kZI,���n��,X���gE㘇O_h�E�_$����V�]�pO��L�$'sN��5J�\[�i4��0ZZ�5%r'Ll�Q���ɻ�/m'9I����G]��}������sA�E�l(1��͜�����	����B������B���m9�O�#��_�]2��Z[�(y�t8�l�M�!NE�R�AO2�Ky|p���h�Iy�l<��=��Ҳ`a��'���itN_,�4� BŔ/��?�{��\�x��``
�R���o%f���r*g�O䅆����٥���_VŔ���,)���X/�x�n6dk��v��Wu��?��,�^-f�������?�L��2��qR��3��̳Y�;��K��0��Lِ���]B�2� ��0�g�pS3�B�<�Z4��cscG�*}]�ǘ�ˢ��
�FF�����#o�`q}]��������;���q� �J:d�Y�Q"i��,�w�iv
D!��b��H�;�^�ҫo�dQ"��
����	��B�ȟ�(�a�t��܅��^�mo
=����֎������I,��^�l�R��0�RJ2$�ARg�4�~���lR�^�,���7!����Y���7���^M-�b2!w�',����2�6D��Z$3M���ѭ�(u�kJ%�BR��wt�)�A���C��Ze�Ϛ���������_ai�	���(q�9k��nt����� "Ek*-$�� �w��]����X���I8f�h�Ew�f3������ٰ�S��ۥ`�h���3hj�����Ul�{'߆u,�3x�bJ�`�[��Jf�[�872"���D*��?�H�_~�@+���/H�����U��p�<��/>��OKB*���,�L�����B����H��J[������ �\�|Vt��,�5N���򣫗��͑��r�����?��/�c����<�&�4�0Y5�������F�4�P�{./�}�'vRAw{��K�t�I{�B�{3/B�Q��fV4��x-�.oh*��"%qoCR[&��q��u''����D]}�a��p�RK)��dh\�Q���R�0����rG-9z�l�<�!��	~�[Z[�p9\�0���c�If-_���~�.̋ȕ&$���P8mn$�GX����	����갡R��_� w����ݔ���2�;62$����
:ڻ�x��?�/P���C����4hEPNGSj�ل��N�uu�l���,�/	z���D%>;ꊏNO����a��՘�'���+u��&��k��9�1c�/=v��e'��i�]g6��܏;T���uǔ�Q�q��]<{�{�C�dst��q<��_>^��B����r��L�X%ަE/���g��̋���'�0��8�F�tR:S0����f�|��f�(��������m���(��6�b�XX���Ȩ��{G� 羋DM��j�z�tJ+/C�ò��͙T�Y��ɉ��Y�����!A*��[��z���e��d�s�#���0���$v��:�Cx�+}���7��Y�$���<�~��s�YtQL��hlj�W!xJ���0a�P�d�K+��_�xEN�#��r�~f���/$�gjwy�8)���Q}}���I5>"���t�������4���3��[�n|妅RV�M�Zz�c�X��yp�AХ��[��ex��ळ��j<��Y�)��:���ծ��:�m
f?q'hA)K	,�⳨����?��t��i�ꏝ�}D�,�m�P%��p3åh"%ω��@w�L
wo�@}MN�V"�N&�������p���C��у�P;�Z�����f�/�Po�B�8m�5�N�k�(T��G��c|�Dٜ���3d���|�:#yfG���NFb�I�P���g3�i+b��},M>F!~��;�+�Q�5����P�ԣ�ε :3x߹�.�N��8o3�;�CC�������h��Lf�g��\�7�}%w���gG�ക�47���1�������He5�7��=�,����!	kBg3��!6)���h�"CA45���u�	��y�vu��~��4:crE����TTW�ww�f�u㺆�g�^ ���r$Z[���T�@�v�3Kx4�J:I�,�uS������\��o���O�����~���o��䲚���������.N�YdM�9�����!���չJ1&~�C8>:���+״]�����.���L�p��d̂΋BnNԫҵ���T���pOɆ�RN�,zkk�5�S��t"w(�7i��EOx�;yf�������CIX�{����%�o2�Y�yi��L�#��Hle���tA��v���q��>@pc��x�7������]݆�`D?'Yl��K'���E� �3::���0�_Mk
��8	rB7X�2��0�I*2��;[�p�'�GjN��y������:�j��Ӄ��%l��kjax?g���Y�
D���<�V�I{f+<�����[�Đ/Y��8�(�T\�9���ǋCz˧�"2�3t�2��L��v�,�� 6���:q���`��(��s�K�S�P�>��ɗ"�tv���C�X�{��٪F��8�ʩQ�e��S	/w�xlP�u�gv�U���������G��=x��$Ɋ$��?}��D�XF�%�7�2�M2��^�/8/�X���jjj��P���-��Uz�ّ���'���Z�"ћ����3���E,N=�AA�,�,��Y�m��	�Z��ѱ��;�i;��w Q��l�ѿ�M��cCHT���E�p:����W.�C��.�
~�TqO��zui��f����2�����ٔ�%�I��I��v�.X��c�$�\&'$����b��ҰY�p�)Ob�I$���������/5�@��P�l�h���\��������%�A�Y f7zG/j������(��Y�	m���U{$����A��
M�B��Ag���z��	:�-�LF_�ǭ�W��ͩ�I�����l�J�h3[�9�i�h�;�IFAg��Wc_��!�$;�AMOO�X0���ן��*x��&��w�g�1O��N�]`sEy���!�-�`kk�_����Tfa����2)Y��]�k�{�t�秤��́cg%�:��GH�}33��;���7����]2��}aSDinC�WFdm�2�!�KԘK'�2��煐���܎d���/'p+�������5���5zw)�#��0x�T1'��ih�����.6|��mA}9�jj.O��!���\��#E��fq��ň�N�&}���X�\ǳ9&_�5��S�0������+��w*�<1��g��͟�R}-Mh�Υ�H��c��+9�p��w��u��"�$��n��Y�F��@O^<{�*�uu�=v8�X�ڃ�D3�%i�OMi	id��]
sx�җ��VWk�&�I�s��O&^>�!��k8�����9B"��rRLR~��4I�х�v`��E��x8���^ւ��s��qQ��鈐Ӊ�u�C@Mlu���3#X_����<U>��c4#�8���78\�Մ^)�$Ž]�C�1�� _�����CwG+�}�$��������sbz^(��mt�*OLo��Z��8�3��y��<
��	E}m-�������� x���kڟs��y����oqUA؍&$�T�����7���;����vN��e:��+���^���T������6���ƕ�ek��1}�*�6χ&[-j��T��&���,�\u1f3��l�F�t"�����	��슘�l�H�!r����4���g���D�5<�ٔ�I�#��X�t��ۏo��B�,c�^����]Z>�]Hg��7+�O�C��t��ڢ!���y�&�m%��!-$h��NE����.w~~VѢlTΏ��v��ꦲR���S��&��=UA�9�"�_���Y2'�WE�B1��XP6�?�'�Da~>��m:3s�b���ErP��hP6�7�:�ِND�Rg�)K"���]6�ѻA�LU�� �9f��ln��,9���i9�v�M�3��݈	#D��*SB2W�{ix���<N#�Uȕ�ɜC8���:��޵��ƺ�b}S��uN��0��s �)�RA�L蕂N�7��.��h�hH�0\
���O�/E���Yg�L��ϟ��U�qN������~�"�{{?��dMD���ᓰ�C\W�xT��d-["9�h���jį�l�@�L"bL�Y�Y��Ar*ItٔS3�YȩZ���gC�HZ�̓����`/�^N���X�+�Dc�
�ܫo`J���K���AY�����Y�%ߣ��{����i�w    IDAT�`��͍�Jv���J������aGM�$�4�1���HqXcC�[�T�wISM@�H=��8<�i-@"��o��8�?@�9�Q�O��FO#�/���R\�pvpH�2�{8	�@��h�7��a__[��(���|�M��"�rmE?6c�䩜�*�n�����;��j�<Ø�}��/�N�	|z�K����R��%����߿s���]X��tr��~��O��+Q���,��{�b{z/�=�-PN)��H�K"��f�N�4,�	'��g�� Ty���Q}k���$���F�92z�u�Z(F|��¤D�<�tT#|h�C߸vvSNP�ᮾO�X��Q�S��H2�҃H?�S�=]ݚ �_#Q6�������_��ʋ����y��\���07�`�P����hnjW�����:!���T�9�{��7z]�0.��P��iB���	���.Y>��[�vw�������J�  �ǃH"�Bd@�\Yχ�>
�tv��}i���x�bA"�pX�l�Z��p613'�I;k�%DO%!��=5�T�m�z�hZ�g:L���f����~����I-��ޞ-}���1c>����.�ׄ�|j
�'	x�A��ȡ w��YЉް�7�����qnG�֚���=��)����C�N8Bo߀�,VĪf�Ȧ�Y��W��;�r~5ϴ��\.�����?�ŋQ_�E!rA��WO�aeuK�v��Ryd��٦uC�s`7O�^,��$φ���[絩�kk�"֨��L����'�e�A�a�t�K=���e���#�͠�{���O=F1q�ð���o��[}-2"�J�ig6�G;�T,���A�^\T��Ј�.�����/%�pN�+�I���zB�l��f��$��'��Lb䙓�B6��s��P�Q �ޞ>��w�a�x�����@��EP���uOU�N�i"GB��{X����"�}�2�a2��G�+�z^�����������}6w�n�K���E�<��T�P�ې;z���btS6�$/N�U����8�w���G��r�׶�Q�؈#�l�������l{�U�yz��U�TG�b�=L%�
�{_~�>_ '�cY�Z�y혉���[��a��7T�q����Ai�dxWX��P�ɻ�Ѽi��%5�<��7���ߣ�3����`j���yv��M=�k6*��(��>|�
:5պ��ɜ,�|ɓ"�L��G�,������X�$R3��;x���!����k�N\�p>�Eu�Ѻ�&��)��)y�p'Md���M-UFTj��t*�R��#񄉕�8�?@0t�v�&y�]����#?4��¯�7H���Y�Y3�¢j��!e��ȋa���EM}�qx����L�,bjy��tS����/~�Ε��nW��?*[���S���_����|�S.;��������f�"QnV_݈��!஝�h��K��,���\>]]�["�,-�byuS���D���U�SI�tv��c�c��r���
�l��	��Ə��N�T���W_\Y��֖�`B��4�d�I��{wojOE(��&,�4�`g�i||��w�&������_J~��&����LcccK2��=A���?����}����\v�b7��zP��������7#'s�P>cK�Y�i�H����NM4�t���B$X�� ����y���(�,�d�V�����*�tn�{��%c}~qŸ�|�X��*��r�J c�^T�orjV�W�||?�}����b1��>8���!�ܼ~C�qL}�*D/�Ê��4%}��`���l,`��;݆͖��i�U��sT=�f�I2G�.�l��M�uB:�Z�=M8�h�W����.'2Z�2���)'ϒy�N˥�{K2d�P*Y/�e���E��sFr���m���(d�$�R58�ܥ\���iM?Y��LML����,6qOo�\�|�~�l�brz.I^Q\�rUϗH,�`y������?���HJl�h��6�
K��`J��M�f1mp�ub��MX�M��(j�����*��7�^E"վ/�(�xd��W��dkw��⪬t6�
��/'�F��w��f������ܿH$J&�8�j������	M��L����Ѩ��|m����iL���ldID>c�����gCC�j1�߭�hvv����S�İم��큁��I�N?VA'K��V����+�cAg0�U�M)�F97�8�Z%�{���>Ovz���z�l��WU+%��W��pB��	R�Ն�鱦1�1��D��Ã#�}�s"���z1���H<�p"cL��!�A~����P}�xќ��4���� ޿*`~ȁ`�"�~2ѳYx���ˉ������%	���~\��
�	81��&�|	[.&ȟ�_�h�}��MԵ���K"\��M�T<|��~���k�u�00��<��l�I:��*�1qT�ݧ*�T���;
𸬸va��Ɩ9=�~|kg��1q�kS�@�]&/R2M�T�ڒqGRa�͉:
*��P,"�����`��&�h�uKT�j�P=.�⪕���H��a�g�(�-?O"�U~z;�p� �ǧ_}�p�<��� �j�%������\�7w��CA�M���_�Y�`�����Y�{�n`���� uE������)��<��`����5k�q���:e��N���Y�f/�J�dcCf$�?�{v_"=pω�f@;M~:�����pM�������F}l���Lm�a��C��î�_��$��"��d���Mh��4{;��و������"Y��Hn�u�lm�Mx���"	be�>6�^�ά^�au:�]�ԏ���>�y����fM����%�c�4�"E"w����ojS�o�����6R֌�<������\���x��3��F����he���%,�B�	5��J�`�����c����U�;-��������,�^�� -_)5�$Nq��)#rEKk���}�w��=c^+�#��!S,�ѓ�Z4�����_ z�CU��L����1�����Ȼ���j�Ć�ڕ�h����ޖ�qD^�����{$�㊇|	R7*�F�������"�3`�"˼� +���G6�.z,������^xDIx��׫�P���i�v�2��ڢ���H�H7���Aխ-�:{l����)���}h����}��'�"�p:^_����S�2�*�<��UM��r%g ��A$����$���;:p��%]�4��;I-�����P�dE2������m�+��o���g�6�� D�<��ϞAo_��#��4Ǒ�NN��1J�H�"1��b<�L����xѡ���+����s��Ӆ���2�����*L<ӄ</_���3'-�0x��D����x11���=��.I�V^ae��G[��ED�V���K>��M�=�|~څ�=)d��ނ��V574e�}�/P���M鄐5L�АJ�u�x6�j����c�sŝjX��=,/.�$H��(nߺ����#�z@"��y%W(�<� ���֖&45���/-�b��P,w�%��l���Y����>��׮i��d6�}8{v�KX]��3v8Ͱ[�{��Ö������);��s#o�S׬$L�
yy��Z����8u���,+����i8�����c���ɥ��!5.�L>�dpҶd22a�s�9��Z3ŤY��K�%���'T�n��7��'ǃ�+\nXK&��ڪ������m5E�(e:U���	�"�tо?��P�u[<�Pݐ:��@�ښ�08С �ٹ)l� m�H����;̙��������X�����gZr�.�D!�i����$]�B��W���m���9@�̰Nٔ^�I���Sik�����ITM1��,J6��!D����{�b��JoK�M�E���/<��L<�P�X,/w^>n�N7c����.��]C��̀z[�$-�]8��bcmS{�_��g��psZ�����Ύ��gΜQ؈`�� \>7���Bx���%��B�
�^}���p�D㭂^�<����E��⨕&I�u*ÍK�N��j����*})'�`���n��0K��mA�6��Q�9��A��K�l�8��W"��!�J�Kv��.l6�|�Į�e��\�鷦�Ul:RI���>Zy�*h���GR}]��c���/pO$<<B2F�@��cY,�[^i���m6!�����_����e����}g1|�=��nu��g`By"�	��}>�UW+AizfV�9Y�"dfd�o��/�rSD�CNc�B�z>�E)�~�2s!�qiOhH��t��^���뚐,����5U���N"
��!�Q~}�^ t0�ڇE�A� ZZj�fD�9>�-mveAq��?�����2������I��
z�qcW�A��C�,sIa������t�g��R����� ���.mmٸ�31�Z����5VCģR���`� ����Fnmt�#^BR"Cjv�Cp��zD@�:�P�e.:mi���A��f�N/��[16zF���|$�@�U(�<�dA"��ϓ�O4ǅ�WKf��kH�ی��i,O~�dxWa)�"�gղ/>w�&�jtyl\���b����nom���a�i��z�|+�bi��t��U��J5�U^�m��3G�3���D,��M���,�Y0��ťMA�U"9W��́��p��8rلк��c5\K���َƖf5�V�He�x���?�v�Ȏ�����j���R9TWS�>����̻�a7
:���L��׻��@m�0��j5�p��ͬ�-� ���F�����X�T6��q��{zv{GG�ͦ&�����h^���|N��&�������@���Ⱥ�h!�LA;�jԨ��Idse~O��S�	E��Xa%:h2��y�K[;"�:���.�Ww��������>�[h�?��x&�,���p�X$�ϊd�Ύf$'X^�E$zo}�LTA��ݚ�o���^��ont��;�7��<�?����_��'E��b�\�i4(�d�$� �q�X�Fpz�`��$ձ�m͂��#�[Dm���eZa�;�����S3���U�ҡW&t�����l����d��(�8S�M2��n���u��թ]]�<��S�� w�h)�*�0��Ӳ�I�Sq�Tl�ņ'O���V�dN�\��QL�,�Hak�P� �]���	�b�%�W'`�]�[��e���Y�˗^��/0��p�����rB�����|�v��o�D�l�f���ߟ�%b#�Q�j����I�ϐϔ/�;$ei�IJA�$��?S.��1f�b�Z�e<B� ^��\\�X��?��$t��/�A�a(�����ڢ��F�-��@\�9O�T�&ҰSל��?G�tO�z��FG�Fο�"5�44av�Ū�i!tVʣ��	-��z<pRS],`fv�6At)�*�a8$~�Zp�����\�r1WagL(;�tZ~�	�N�C7��4�]T2
���kdx��j�+�y���h��׵�gIM9�tf�����jy�\T�gį͢O�Z<JRS	'E2���}^�o�a��p�bp9�}��iX:\~t�|�����&c��z�޻w���#����tg�)'s&��J/7�:��`A���r�,h�j)7�q��񼑀f�+�"��=t�2��؄�l���Zt^xdwv�v��ssc��kB3�;�����(\-1�ec���+�!�䬯n������Ԍ���^o��s����ۘ���clΣ��@�d{SЇƯ#U���Q�p�<��0��>'��w�?�/n�|�{{0Y�0�ܥ�R���S��0*f�WJIP�8*��W{����7qi�]�����7-�+,N�.�߅B��83܇4�%'KH�3Z{���ECc������b������䮾�~◿���:RvH�{~��e�(B��6aq�L>�K:*��&�:����d��"e��l��ܼ~�Љ+ZԶ��`?���!�>�>�L��J�� }i��;M�h(V�6���j5��g<��� S��DI��|��=9��$G~Y�lr�J�4��z���j�k1����pD+	��R;��֎���fҲ����OG[�Hu���q��Q�ռ3�f�.3���=����lB&��}}G���V���l_c�_������;�?�r��_�{����~>�M��4�K��^P��>�!��w������q1y�k�P�^� ؏fkc� B�G'��*���⑰o�ԥY->�w�@kL�|��xʓ%?$�r-��v��u*B�;c�.k,�����	��s�������
��Ȉ����Ο?�߳0��?�l폾�1�Ǉ�jm6���+^�P�RDbqx��p���X3Ŭ��]o/��9vצa�V��eȽ�}���")��E�ٿ#Q��&FPR%pv���NHa��H�dZ>R7��'�`9�E����&�m�ƃ� iCO��
�d�����T�^0ڐr%�l��*�l��0<8���}I�דX�JOh��!�P�A��aKs�����Up6-���m`�g���]��E��e�����O���b)�К\�8oL�f� .~]=��|�gGpnt��� �SӒ�r�Ν�;�]�h��v���%�.*H��LV. NF<7lR�}�����9$a1�&��Kȝ^�t��o�v������41����p��=ǯ��Z��w	����Ù�_��f��9��9dRy*E�9���"�&��-w�VA�"�8��W�yS�y��>>9Qz3MK���ꧬk���^���@������g�a��&9��6�z�p$�#�_����J�� ��ن��F���p��"$O��'�2�Pg3��˩	=K�t�w�φh	'��pH�i2F�`����������{Z[W��qzH�dsj��2��+/q���*�]�d�A��E�]��S�
�?�i�HW.��Hf�J<�P�e`�9uL�;@�^��~�O��(����6cA�/"�{�*�����d*&�QSs��K�y���K�j)j@�Iޅ�M��kq~Q����(�ojj�Z1��J�sp�'�6����#=g�{"m�r�{�jǡ��6�ǌ���*��TDֳD�*�;w莪z�#��]���'����k���濫����a�˫��܂��|���yJ�5�|��b*�����{��O�����A:]ԟ����+t�dɱ��lwj�@CO��� vV��gB�˹98kj�����jP\^]�>w��W��¹�X?x.y�Y�{�z5�LN�p|2��Vd�a��q��5���������߻q���߱��(b���L��ׯ�����RtzǢ�4
�L$��30��q������DsSv�CJ�b3�1h�1���z�t���r';1��*{�l�JA'��Fr�����z��]]>Ɵ�"��润#e��Sa##�/w˼xI���t^�v���+
�p:�8�"ͮ�d#���~��������)�	O�K#ăK$�B��L���%##�;)SɊ��^�~���9X�i.Jf�zs�9\��Ds&u�4a���j2Asm5�^:��c:.A��q(��㕵-x��˺VÆ�ߛ>�2T̟[e!����4�6�">t���H��_�0���D}3�c,�dm2��2<��f����S������]����V%�3�s%�I[���5=o�a|�m�ҡ�iĒIe�o��SY��З_�
���VN6vd�D���*��T��H �������)����dm}3sK��	�3ԇot���*�*�z�(�+%5urڔ���%��I�7D#9[Gs�l�-dw>��У��J#��^��o��g��w�a��h����MM�Zi��⟗�屵����ETU�"���x	�˘�| s��MAOf��,� ȑ���gB�.����X/�)%�������.I��5�
D�������Rf�Ӟ��93���nB� L���2�݄tB��BG�4/9�;�ӱ��������<�z)wcb����z�ݝj(ɸ&3�s��˃��:]�ܣG�1�����6�����ח^bs�)�Ǜp���t��7=Iӟ���d1��?Nj�k�}`�OP6m^7wv4��P�0�*�+CY��    IDATĦ�b��oh/%cB��)G|>|~����b���#(��0����Wբ��U�'�x�
�z��z�hnh���{�-�q��Y�B�xױ	b��Ĕ�,ו�r���ѥ�Gi/���f�qt�2ĕ�͚���#L�0
:�vvr%'ʤ8��Fg�<����0r944T	�e���������!��dԍ-��F����}�!���V��
:�\��������>C�]�	�QW�U��6�ǀ6�6�\:P������L��͒n�-/���dBOs��l�{(C�K9[��D�JD��p��w�S0t���.������a��Ncx�W��S��O>�n(��ov�\�Uۭ�ކ�����K��;����/�ͣ�l�Ռ��Y =@¿�ӧ�.-�b�T������H��eފ��cu�Կ�׷L�LM���nZ�Z�?8$���g�p�HJGʽ��N���4�p{Rɋ!������ˇ��zE�l�b��D	��" ���zT���u�֔e@<���y�	�� �`gJc~ ��%�������@Jo��L�XDr�L�3����"Lɸ�N艼m}q����(Z��$�����h�`�YE��-ͨ�����Esg����d4�N7I�=���zeb҅*�e�ؑ�-�ˣT��mjiVe'�ɞ�X�]�.6M�?�<X�9������Q�6'�c=߹�1��kt���}����\�ρ��Ei��&�x"f��(�pJ[�jf^M
�xs!�xx/����Q���5��U���%�Q�/���Q"��GŐ�g)�2�C�z��j�z8f0�����]���!xr�G�0���:/a^���c$��H��v�� øY�>�Ԓ-Kn/:c�3��,_~Z�q����~��sy����#��{ﾋ��u���g�=��@go>{$d�F;D��6W0��+X�4��g��vAg>�&���m�EB:k���h%B>�������4{K��S�����Q��C�;Z��ߚ�59k�Y��2Ad�l�N�Ő0eT�DBf$y�d#NbS�O{�e󼿿'$d��9tvt���~��O�jm�9�އ��OO�RD�Mn����(��D��yt�4�׊��6�`oc"f���s��	�ۂn��h���T"���!����"��Q����i8%�V�%��Y�Ig>@�@�ʄVʹ*��u�|��b�&��p_��8ܭ�����Әtڵ��z�O8��>���n�E΢39gMLM�N������"^�r68TI�^U������G��=�"h��� ���o����1i�i�J|�3�n���PN�;?�@�%��rz�Y@"!Wqt�L9LFG\�d�{��@CUbx�HrFFz� ��'jȿ*��T��$�qPr�"���Q�0I��s��߀�l�C�,��_-.j�OC�$h�h�W�F������z��$�V�qJ�76��Aǔϣ�ևt2���5�7��T�?{����\o}��~|�ҿ��������Ͽ{r���^����?�Ȥ�H���ڌ����O���'O�"b$�0^���ēN���ᒜP̦��֮˕d$�EYݯ�ܻ���"c�JwZ��iZzâ%/���4/	K�&�h��cM��%����<�)�e�({Ԝ���AE�1u�,b��)���ϝ3�:�9�{��o�<O�6���dؿs�C�������j�i��<�N��Q�G��x΄��˸t�c���(�jJx@�Ka�_6N8Ό��p��	��$9�Α�;s����oC�T���m3������ǃT]UkX�2#�{˲)5�|iy	�`pH٫��T^0�"�R�b���z����e���k��]�tk�X�_0$2�z��186����������9ؑ�<���7]�d�	}h�]��K{o������ę��/1Wzvnk[��?P�;!��h�m8�����Ɇ�X��i�Hx����B�t�IY<VEJ���>�������}��eSD���R����I({��
Zo_�������4�՚B�70�߇s���ͧ�6��iq�p:=x����ٌ����W�&�<��ܱ
:�)��ɀܯ��'�T�x^���f1��	(��0!/���V��2��k
�̤#������W���0.K=�Mz�8:8T|���FKS��)���}�I$j��
20����q���QERJ��0Z	ao�@�K�Uɭ!3��,A��M��e6������XD�z}~�.,b}g�,�4'��$v�g���L���J�&{�ot�-��mu"rt�ˌ��z|�[��H�[X^�͉4t�:)�K]a�8P#o��_���uғ�"�r�~�n�")��F�*"j�}~?����ж�5���ϟ=��A��:m>~�~�}:���G�g�h�}�cs@�[M@�=�z�y.6�vawVk���}i�!'���y��l����ѫw��+���#��5���Ȥ���S (e���}O�T2��3����
Ht��F$��E*�B�2e�W:����͖��S��J�ϲ���sg�'铀&%pM�mpz]r̦�hk�G�ӎ�����r��W�_�\���6�G]c6���r9:9V}��q���Ω�$�ϑ����>��%C���&�k���?�D]} ��>��}���=���Ò�m���ߺ�?|�������_?�`A�$b�X������lFkW�<���k���!R��T�~;�X4$�۞�6�UUk��%M���/���ň��L�bn��	�%ӣA1����m�\&-~���CIƻX��
e��E.����N?���-d�"�t^,��tV1��P����졯�W�
F�K�_�Q�$�]�z�L�3S�o�-v�mcy��
z1{S�cY�s�
.��)ؑ�>�	�����>k}\�0n0,-&�()[���#|FӐU�����W�$�{+�\�R�W?�"Yٌ���N�c9���r���<	�S'�:�7�|���.Nwp'DM%�������⢱������ &&_	���֏�Hw?�P?��ʊ� f6!�Մ���{��P>��C|a��(Q*h�E����Ӂ�с��d��{�ꕬY����"���j$�4��t�{^��J�!��|�|�Dnty�S����ɤsz�����l��K�ͯA���sa��NY�}x��wp�ԅ�?ogsKύ���6�o<@M�J^�tKdC9:6����H��k���*f_>ЄN�m�OɜU�C8{��
�1�[�N��6�YM٬���ϔ�-B�߸���Щ�(���%��*�|~���_�as"c��B��D?w�4:�YW)侰A��T�'x���&Ԑ`���q�SY l6O#�.����q�v��/�>�r~&W.^й���6v�V�08r˫��_�ng[��X��
��!,Y�.o
:FR��HX��yuq�u�AM��hH�;���.=����W|hG�8�~P���]w��lFQJ&bB�����(3ޝ*� �U���#<�DXę��p��(���j6س�sZ�x��084��I��-��ڪ�yMm����~���kuA����n�m�b~q]=��R!���ǘ}� �LT�jw+?��cg/߅��E��%me�c2����062�?�`���;
��9�~�L	#�5ܴmN����RE.?3���Ap�h|E�[�
��)��Z��Resͳā��/��hniB:��K(;���̿2�":�����.X���9q<H���n\*�Љ�cg9��w�??���S�ۈP�p���ր��zTU�����{O�Du��t��x�ڿ��۾�N���/_�����[�#t�)!���	ζ����f�M���@�yV�`�;m)�2�!/�1-V��w�"vuvʅ�nP��<\~�.d2�+;���^�2+� =�h
9�HH�S���<����;$�M�<�8���Op��yM��S��4����W,�`�&���dP=��E�
�߳�ӵ�Տ���GsS'^MLbcsݸtbI�#GX��:x����#Y������� w�/�@�[��<M*�:�P[���g�X��;��ڎ`$���ؽ^DbI�Q2���6���I�'&J0x�C��I�6.���}�A�Y0&��ݤ
b>�)���s`�:��$��B><
�;;>������.N�\Yp�A�!f.�����YM}u�`��V��?}j�'�Ua~꩑zݗS!w��
]�1v�{8�3�X�O�f�f\:7&y����n�?;:�l����-��2��{��������r��:
�)�ǅ�X̲L��>7B�V�Mϔ;pB�ULP
������s/�sԯ��^Ng���2E�w�N����u	n�C�:u1�%�bzi�h\�3��W^am�&t���rRy+j��`�����<H��[�E�F�r��έ����{`}s[�?��i˪t>��sOk<�
۽Ҁ�8��Rޡ����0N���QP���q4�~�<��.���ǐ
�O��y~	��Yr�E�u��@��\|���yWp��UZ.�U<;2,2�ƝbB>W��~�݃ �O. ��lK��u���"6w�v��cW�y�D5rg@��m���nBC]�
#�?:.�kk'%�e�8r0�j��d�o:5��]h���a	��lth\�g&�?Ϧ��D<J��{wo�m�v����!���d����W�]w�����:�HDcʡg�a,-����ciqE���[Z��=���䢔�%r��}q3���QL����fsr�Fm� F.P�ޮ��Bw<_3�z[��z����?��3F�<?{*���s���CN�����J'��lܧ[}0l��؆Ý�N�.�g��۵v�;���d�l�s�9VuUWN��U������p8$��}��_|�v�l�A�&��)�p:ZE���e�
r=4��\Q�WZɑJʵ�ZE�fL��NJ(|����6��ꗅ�Po7�*0��v�6�[<���M=���V	2��5��b���3פ�nLH�#�ϙ�����p\��ވ|6!�Z2i�)������^l�l[���~|��������G7~�h�O�p�1٥R��ίQ����O>���Q�b}q��Q�m��C����ǃ��t�blh ��3�lmn�ࡥ�C�)x�e-[���.��wEތ�)�I����84�!�$����� m
�pr�`�E��W`&RH������z%�h$b�j��§�L�(�l�����NC��z���!N<����yh+�_�x�����L4t�f����>bY�:XV�-����f�uwh?�j��4]=h��ă'����� ^J�%�A�8���Ŏ�nLCD{�X�d����j]&l]0��eGˎ�#<B��	�i��V��C�7���  U�u
�T@cХ�;u:Fqd���m�ײb�����,F8����)���ˎ��UL<�D#�RB7����u	CW�G8�U0S!Cf��cRr�����������P�}��2bB'}�;[>Sɾ��߭v�"��D�☝��A��6���^�Hx�=c
�'������ЉCOi��_'咂�;��.�ħ�{+�N�:�I�yn�S���G'g�� M��E\t���42�Oԡӵ�	��y�7�A�D@av�Ujx�3ĘP��TRee$Sq�wvcfv��G����&�jdy�7&�R�e���aB�q	�65��&���,(l�[�t't;�Z���~�*�^��g��r%F���	�?���B��9����p�^D��hmjTw�����	ZSSOB�[��>5���d��_�tw>�"࿕��f�T�=��IM!c�|�f\�2���*���q|r�	׃��!�5���Y�Z�JSJU�MC�v��_���L����{,S&~���W��n��������8�e�J�{Z����cem݃������<^��Sqr$KP�=o�u���_h}�I��ܼV-��w��}���%"��~�0��>�8,�r�:�5���.߁��I6�.�w�$�KE��������dz�᯶�Y	�����݇"�R��<-���sF�ա�XI��dX{��2S\F1����ɼ�N����{�8素�VfC�|=���=��L�����8:һ�o�:�ϐ��TI��ą\$�>;MJ��Nł��u,.,�!!_=p���	>��|���#$H��Ѭ�(��|����˟ܽ�_���X��������_<z�V�����nW?�w��&�47���^t�v��q����������$�|[�/��jA��@Y�{��������h����vg^Z��*]��n��ɩv��bQ\����͈��N١'�R�aB�^��]Z<�,^(��g@	x}�*�\t�V�$��P��s�YL�a���r'�{������G8�](�2��̆M]Wp�ݏpJ¤*�p	Ka�@Ķ�z\�|I�q<�������G8|��¼y�É�"�K_R���j�j/4ꩩn�AG�����q	jL�~d)�J��|�X|���&��ύ���R��dJE���� @\wҧ����
�����7����l�像5r'm��t�����.���E^���g�i�c$��:��+t�r��L$�x55�}�>�n!dK�7�7WEh>o��j�+�ݿ��D���O���gRϯ�*���1�c
�J��s%e��^UU�_#���#�/�42�PGK��r���?'ւ\p&t�׏�9/�&*$�3O<�{�%��Cg������u�7�A8u�R#cb�4���+�}S/��K1%����#��Z�5�Ƽ�B�bd6ޜ�;%��&�Ϳ��d��Č��\�$1lL���ɪ�G�L��u��\�~A]M���Vb����s�E����fm��$��2�k�Ŷ��ahh��C��xW\#�5r_Z�Swτ��1���qn-������Imb��5bK6��pGkf�_k��f�������	(-�Lў���FB2���$����X��ZH<P�P)Ԅ!g48��I��G�WG��h����㒩׌�U՘����b��eG$����*kq��Mٌ^\D��+#��W�T��r�FH���������(�Ͽz�.ݖ�)�����y �W��W��e�&��A��YRE�:�U�h���\A��<�D4N��QDQ��a`Z(|U���[L��,��'<Lʼ�6�MkN��|�xF	�̗���5����E�M&	=�9͠? ��Y/�/..��g�ᙖ[(%��Y��`��ό�l��xEM-������PmmPE5G�-��x<�S++�ЙЩ���r��_�ޭ+������ߚ����~��'O'�����iK]>x�&��c�l��s��wޅ�����>�c�����Ywi�A�$��4���=�`���v��an~Q�$�9��Jh������V,	DC���(�4s)lAa*u�'=�7ݒ����n *ͦ���
��<C��M����0jT����u�2�v��y�x�w�70xX1C
�A�/H��k2ga���e��Eq��:n����J�]v��,������l5�hinT������:R%��+�{���\��~�����31٬�� �">'&'>7�S�`H[a㈜ܕ�C'Б�� %~^R���2ق�ϳ3�ΐSo�n8��j��Q���wvz��E�dV+�n�Ά�c7aos	SO?C2~
�n`/CK�e��E<ie��	Af���sۭJ�f%e�#ޅ�e�r�5�(��v侭(�YJ襤^��K	ݠ������$)_t�"���u�D�F�~ҡ!C�ަ��ɾ�?�s��Xq��?o��"����lGSC=�YT$�2��6��a��F��J�I��չ	�.��)u��Ͽ �\�����$�UpbA��,W�ą:��.���]tM�m~���z<}�R��r��rCj�9��d��w�(z�yCn���i�[Ԯ�h�W^
�f%����*%k����L�Ѥ%�Q�K�o>>�Ӏ�;�ֆ��|o�`�mA�MQ�2�e�*l��4��z�
�;���[y���U�X�f��^���K��u�b�	ݜ�����
�5A�,��`_񄫲���.��صڽ�P%<��m+i�ӡ;������^R%��FExv(;=�y6�Sq~����р��\P`���.�������Q^Q�4Q"    IDAT���x�b��G&��<�? ����0�g��g�{���]u�LNGF�ٗ�5r7g�!ot�5-���6��F	;�j�4�	����W�8L7���3r�ŮBR�,	��Ɗ�l�6�Y�}+��޳A���p�h�	������ Z����[���XS���VX�9M4���0���	���WDю�c�5��MX]Y��⒞�;o�������FA��+�Ӫmh�f��`�݉�r���S��?���n����wF�~k.�����w���w�[�kB������=�\��&���/���w��a��&�������C�^�A(���O�At	�:{{�#-��������xxqi��*D����"0G��b�2�H�T�FB/
�P�� 	�|�ҡ/%��:6V�i��D�`�*u�D���Y�b0���+] ������*$��f�?E'9��Y������^}���9��2Fn�ÍӋ4�/��Ko}��I�j0��:D���5����ݷo#
��ڍ[�=<���*�O�G�ыbB*Ip��Q����h�f�<����<t|�G��\#��Q�w9*������1x���Y�������e�]���'��1�w���ʕKn_D��aGK�"�tmV%���5	�dRԳ7h�L��л�n#��:����I )/,(:�ۅ�Y�{��?9	龱{�ۋd���IZ�r��0�ݡ�g��E��xRQ
6�״�Eϟ޽�(N�a��8U��hS٬��@��E�|A�9Z9r��g@:�]~6&\"���Ƹ� C��Su2K��Ƅ�I1���&���I�ɬ��71x���	���(����2)�=���{w���$1R��VW����0�ܑ3)0+�
WR'��5���q�JS3�k�g���C�#a�,r���3tz��P]C�ٹ�1;/�;�Q���g���$�{xt��ǵ�r9��(e��^�_��'�F��;������`���^(%��ٯq��� ��2&X�uh�C��U�пI�2�%�b5�02؃���)*sp ��p$���_�$�c�������C�[�b�R'�w[�T*��j��b�����dR�%S;����hc�ŀg�[�!NQ��L�����ʑ񓉟�w�g��������dV��A��5)@����p��(��<y�$��kw�*o@�l��?������6��ڑ�%���hh�GGW�ZL��#��jz�3��.�W��J�ȶaYbD�-�@L��0P�L)Я��o���Й��P�D�|��{��8Z�l�����Ů,���@[S�&
++���nm<��[R���d:!�a�o��>�W���@SS��}������O�tr��`�P�9_��-��/~���?|��e�&��g�����?��< �x����������h$�Lށ��(�C\B�=�������s{}M�?�$��,t���]Ѯh�t&��-�]J@'��H�C^�TJ�bL�&�¹�.Uio��"���jfL���Me��y�*#x������L@;[�2�ר��C��.�p�14��MU��@5�ĻN(0x:!���ϡ�Ţ�p�:��0r��zg�� Z���B��\!�k#C��
�Y[Ç��@`us��_Lh�dq8 K	� '}7)�Y�2ZJ�F�R
F���?�V��LR���K�N	A�X_�`�+�k�59��������V�M�\�
�@��F:�T�˧��d�O��+`�p�0ʃUZ!L��8$e�|
��mL<��L���^
��:+$AJ�(��QR3����b�%ed�}���S�j<}9)�m*k����"(�	�ԉ�C/���WiJ�gc�YcL�w ښI�T�Q�]����rdhX�TvP͍M�d,�Ψs⾐&+��p8����V ��z�.��t���}Fr�����;�X<��OIЂ����ݘ���_�:G���]�L��iC��i�j�	N;G�簙���f4��beeY�P�����{�����t�vB�%�kQ�,Ǆm3��̖�g�n�Ϝ����Q!��EĐ����8==X�I�,"�%MBVd6��(�d��`�q1���_�`�7ơ�L��B}�C	��9N���>V�whU�<� g;��m�g�['����+�rgB�a��ڊ*��2_��|eЋѡa��C�]$�����ܾ ��:t����E���W��t�����D�S�(�$ʢSS�����%���:�+;O���i�{��\�ѽ��Cc�����2����gw����L#��=�h�XJt��n���ӯ�$��l��u�L�βz)52������TI����Z��N�������5���(q�f&s%�	�7҄E�˿���5D����q��Љ�$�2�I�a�4�K����t�CE���^�mE�Sc�{~!/>cG��H3'��M��u���Ȍ�i�j2F�m��;t�͆�:��4~��/��������C���Y�h	������~z��k��&���_���O�7�O�������>�}~TY궽�..��w����6��:�\��J��`P��'�``pXA`ec��
u�^���.Z�1@+����1�+rZ%.c$o����S�g%C�J�UT��~U�!�΃\U�V�ݪ�hY�$399)kJ\rW�n���<oy �R9VUj�'
��6����	�`B?�[���O��1�
GV�{I0x���T`%��A���=��9j��u�@q���x��F��>�ꁂk�|y���E_�AH���*V��8�/=;�z)�B��4:�o�������5��҄��,�M��� ##C��.���L	��DSx�� j���-���M&�@�#�6���eը�����^LM��̱��J��=i�r���C�����[{�#grkU#z��Lc������{�-��8�ZYAOO�.Ы�,MEx�,���z���v7^Z]�p	z�4�`������V�k��D�#�q�ƃ���ȝ���?�!�^�c�Eu��:���Ā�,-�8 `��e����I$2X[����!N/�Z�0"�b1�쯽I��q%KYQ�4���!ar"�3����?%���s㑐�-�W��gbr�G�g�q��GM�"Z�A�k)�#�k�Q�1��0�g��3�yh9!��v�`$t�z�W�� �Y���nt�Ē466��_c��������1�|yI}���3*힩ϕ
t�������#2}�{m�Z���ėHF��T*k��S�&��:t~�g@�H�������wVsO=Fcs#��q��1ڈH�IX&K�s�z)0���M����k��)i����8��y<��҆*�MH|���,T�3�zt�FL��m��:�N
�n�8>KC�tD	�ϐ�,�+�?sy�bɄlK���ă7��*�fj[���݁z5%�k%G
����
�V\�4$@��yX*����\Z݀��r�G#�}��ʧ4��f��"�$�z(��n2(�D���Gm�<�4��4a��*PY�ǩ�A�/�S(w5��8�����%']S�G,2
z�_��� ���Æ,z�W��l�Ȁ��6�;<�(Q��4Ѫ�2�=���p�	��R��h��\��{�o��n_��oM�����������h ��m΢��
�MB֦L9%� e��8��`1���v�kTH�U�(�Iu(���<z�瑈�e�M%d��`�ʛ4�l�٥8�+ڦ��S�<��еW��=E}��A-%.v3L������Asc=~�W?GksƟ?C� .]�,�h2��,G���	��`�ͪ��ni��C�����&���P\#��hWC���,M~���y����fy��@��]���Y��>D�#�l>��,�_*qϠ��\jv�f�S(c��T T$+Zc�'��,B�7T����J]�:���IZ�K4]}ilD�'_?�?rq���v�=lmlK%�&4 :�Js�>$]�U7��cÆr]�H���d��%/	�qm��`g?�1����bBK�`�J�]+'1�t\��L��x��&�mxx�/_���"A��:%NExƸ6<���EuBV�~�hl���3�3}������x�D�r��5y�4�H&qixX���ϟ��d`�<vINkt�����4jfnV�"�h[g���a������[k����@={!�si$2\{x%C��0���q8��ʠ�PN�8&��p��F3���WVb���'�u����qy�S	��/L�T�"��|{�'~��_cO>@c�w���{����xa���׹��:��7��PB!����ԇ�=����*�U���UG�V�4'�^�膌���%�����'��g��{�W��������X�9��jJ�to�Sp~��Մt�#�z4w����i;J@���E�,�)���&�w��ٓG�riL��;�Bj�l�A%��Ɉ)��˷��q+���u�F����2Ϡ��?�1�d�	�0���+���gs����}$`5��j��_�y���b�K`w`mmE,r�9U��Hk�a�
�M�B6s˛8;k��g0���v��B�L�S	��m�����(�V<,�l\���:��(�������Vl�ak� &�C �x�9�2�(~~#?������]�PV50\s"���˨)�'��?:F,�VwΘI
��\�Q��6�S?>o):&� ʤ9��(��qU��ڊ���NN��U+L�=h���Sj��!�`*�-�O�b3!k3#ʆ��F2K�U'|�,��?�{����O�ք�G���7����pxk�T8,���{p��wz���Z!S���9���1�+�v�@��	Y��H�d-�Mhl����"g!��4k�u.Ot����ϴ0 �
�ؖU�����U��Ob�0�`�ȕ�蒴'6�,<w�.�1��9�U��@�=m����7��u���KU)�Q(�ïC�^�L�(� 0`�mDO:p���-� v6���';�s�NIe(cv�s�6����p�=�U\VR��[������dK_�558�ݑ /%���i͎8O"XQ#����,�h�w��)2�i��u��2䉲�7��������C��A-�>��SuU��+��{{��3�oi�}#;N���������#)x1������Fow�e>���}��!�`X� ���v�����0�䀴�� �8�^���tޅ��+��.u�|�*Ŵ�EX�>���������jgh��uQ8!���@eE��x~(Nr�@"�ci�-v�Y2�>��B�C]����I6�K���\���&LL�T�2��N��h����@7��S��`U�:���֟㯵�w���M�^6ZZYDm]����Ƒh:�@0X�d��@�%t�_#����X��=����.�&uJ}Wn�*�9�%u)��bS�J�G�Ν��0F���y��T��q���KD��'�O~P�Ƚ�}Y ��rb�^��jο�7�7��I�7�Z��.���$��pd#؍�AD�/���,��)����_b`�_�$�"��3&u\, �|�˂"Stuu�A"Sk"��䔻Q�A���p���噯>�^$���lAS�Z���C�mr4����4rr�2���F@��Uc�~��������.�_l8!@�u��qz���(̻��)6	�C�[ʥ121(��5I ظ��^�&�=>S;��D1�ʕKRZ�[����dsI�{UT�����d�ϒ��_�`�R��O����֕�f����spZSX|�T�9�}q.ol~Դ�o�-��ME��?o�)!��*q�҈@e��7��b}k��s!�3��d���%		q��"�S����0�*o��RR+��?kL,�ȥEڥINk�����0O�9��'.�
���XG��}3ڵ�+�E��D�H�,2��Nr�*V��$�

�0���f��k��X�l�F\���`��y�K�vsA�M��߽y����L�����~����4���0����`��~���|�8�����WH�(2���.�*�a�¸3+�ֲ��C��,z�Z�qG�EE]���w{�K&�<��8�V�	�1ِ;�����&��еR�0Db�=�"cg�@��$��R/���ET����l��{q�8�x�w��Xp���xK{@&t��hLR�ǌՊ�����]vZ�T�C������2++6��	�}�6�.�A,K�LNz�S\#�2;�.8�n��W�C�))%�FTTD�I���������A�>�>WnV�J���'�P���U,rύ)�q����Ο����#f�3���ʘ`Ee9�~���0��Q=�z�.(:�g?5�`PmVz� :E��֡�jkr4\( t�j�]��Ɋ8^L� �$�?��;�S�.�{�*�I����|v�K�K, MI݊߃��J<F�9\��p~z>��j���w�ս38���ǋB}s4ƕP�`х7�qY�}p�b��\	x$ ��	G:g�H=/�#pd�x�8�ݡۧQ-��p�L[ś�n��ubqis��C�x��[����,���Z+�p8���-�noj�g�H���=�x�)����X�%2V�2{.�B�l34�Y�ҹV8�Vdb)�Ic@�$a��7؏��]M��n���o���˫�n�T�5qߜ��1xfw�V��tdw˩GBL���r*܍�u牎�ʉ��P�����������MMx�b�}�JB�^j��$�5ٳg�L��F42��qz��8cR��*O�Y�ϋ����X|���v��X�@�
Ɏ�1D�99�1�2u��3��wg[�\���"vv�q��u���a|���y��TN���h4$\i�C����bV�h%���Ϣv��d�`,�\�.�?��pJ���!��hi�g��Xw�B]c��oo� ����O?Cwg��B�w�6��4Y��}z�L!U���Dï�5r��_%OJ�Z
X�~.��B�L+�ف�ū�N:z��T�� �,��l��W:�������8	���1��.�Y.���f4m��SPMS8�}:���STÆɜϢ�E�8�3�t��aN�:�Ϟ m��wa�Y��nE��/쀯, ����v��5k�eR=$�̝��a�I��2p�����˴n㔃�,��<}a���	הy(?L�Vv7qF�A�'�S�A�����o]�?��$��/~����4��U3w�V���0���T�����=��e��8��p-�ϛHO^<�9K%�t�!����ىk{C�\�(dppx�}��ի}q4U]S'�:C��H��A��*'+9������)*��Ғ0-R�D9�t&�Ŝ���FOg�4��W����q�B�Z�0I�����Er���������R�!�A*~����*�N�}��V�o.cs�z��0�o)r`r�k�.�Go�l���E]h��ĤD9�)X�)�Y�y	WT��5z%�|iyA;��~!N��}pt&Z��=�)C�۝"�`�*6��!=�
�����]-�]e���.?�GcC-��AZcyu���v77�|�z������p��'O{]��Ɔ���<�l&���64׵itId�������-9X�I�O6�CϦ#�|���UB�����CC��j#J��0��L�8��<G��t�BZ�d	Ѻ���LC�����>��1Cf����Z��\�,�~6^Tk��h���XDZ�nu`�|��@�K��,<v[�u:����/��6v��K�x�t\�r��%�x�'g��z\�4����/1:؇��VLMM�dr���3S�;ؗ�)�#��x���L�(C�]|�Α�o:�j��Q�!�n�#�;,X\�EeMP璝���%]N�Da�>{)3?-vM9%qi�/T�Yp�C�bF:g`Q���؝+�bb"O\�LJBAE�����щ��6�����_�~���G����Z|�,�yO9�g�纞���	�%r^�gtfL��+�2�ll-Ob��W�'°[MH������;���+J�en��`�w�,�t*.���yH],;����2��'��($�.�E���o�z��1�e�
�!Lb؀�{gS���A�U$���-�"m��Uἵ��Ǎ��h|O/i��Յ��f,-,
�D\9�L�/_�B[{�l��~�`:;3���ke�    IDATx˂Hg-�٭|i�X����S%t��YH[k��+�e�A��d&���p�ͦw qW��19~��o0<z	�lV�S>?�k)�ʢ��E�j�"�0E��a�m�"��J�`>{����Xy����{PQę@�m�*_�?��h��;P&���GW�p3s�3ڙ3Qs���������"m�9�`B�_�}b�W�5g���
+c,l9,m�!E&��&���2%tףݹ���t��;�B�`�G��?_��'y���{��` �u��C��U����k���7O`������צ�]���1�c-���!	Ɠ�t��a{k�M��C�*�����'OZ��h?G�
���)/_�l�5�����Թ+�z��QB?��ю��Դ�&��ۻ:����D>0;��>�H� ;@Ŀ��g�w�=u�,&._�g������5!��I�	x��^���CCq�t&JR����D�w�1�.�K�H�3<�U�;l���y��칷.'�0�Duu%::۰��m�Q�v���EG�FRM�MKW����-���[���:�aq�Ʉv������]��ш��l��^��"|~�$�����"���s�{��wv��u�&�?EkK�|�秖4����yX��L�~�E��g��|�9#�P������.!�b�u�{��m�ŉҦ��Y R�X�E�!�RQ����m���V;�`y9VVWq�"kva��V�G3;n��J^V;��Qeg��G^�I��Q%*E�S�A���'F6���MF0�ي��zu��#�V=�|�����fg籾�%]��w޽���U,�,cxx�m-x5��G������(��S�3��S̯��4�ىG�ْ�{�H'3J��ev��@R{wv"y��B&[����9dQ�������ORV��ޡRmm��;�t�9v��5��q�Y�04�j��%��W4��g+%Y_%y{Q�8�R!I�T2%����`]�8:>���ԼhjBCc=��tx���x�u����D͜pUR�\���.��BD[>\����9���	6_=�:��9tY&tN�r�'�jV(1͑+��\��Ac�"e��mpxD�Z\ݰ�cܣ#�;1��W�fP�F����"�3�:V�x�ƈ�T���"�8_ ��Z062�/A�tG�J1��\g�V̂�үܵG��MW0;Ae%��3[9NN��H孊�D���Q,�z��WaI������aB�vO�2�dZ��	j��ObLq4�7{����Fj����:���s����������&@�dKbOT�cqS�0a�Nf� ���&DyӇ�;N0M�ݔǵ�A�bcmM--�]\ƽ�}�XR�����CL�|!3�g��p-����"����>��bLD�p�.�G:�ֆ47��岃ċ�	L-�HȦ@Z�Ʉ2�	-ף�\���w�~{B��џ��0����SV�lO���X�ю^�������ɼ;!8]^%jL3�@Ň&���䅀S�@�C����Z�Ң����M�l6�]��W�3Ec2���¨��:`%Q&k^ R�K⸈���I}|���s�ژ����u�
��<v6V���]:A�洘�r�D ���:LR$�޽���(;������eut��,���
���5۰�����_UB�ċ�:L�7����Q�F�p;ݰ��t	�rzF�\m�n�O�iV�N�W�F��G`��PV�UG�ŧ����]�}R�ĩvDt����{,�!��عh�n-h���-U���ֵ��eI�'j�s7Dm��n�D8t���=�U��wm�%�^�˫�N����,�ff���#�������T={��5*���rg�Z�p����0��g_�TH �H�ᡷ����gɔ���|��ۡB��Ƚ]��PYU���|�AuU�hN�.`��=�n޹�}��W��*и3G���.��;M�J��!�2�կ;����Z���,�4�3Y�+��A6AW}5Z*�Ng!Kdғ�n��˗���e*2p9�n��H���'(�v�e�W����k����<���N�Ne��Ϸ���չ@�e�H"�wH6�;��Ձh"3���������/�E�ș�b_�XX���~��ei~	��}hji���6&g�T�G�M%��Ɲ���,���E���8�j9U1Y>�_���N����PSU��&��uܸ����Z��t�y�y���r�1==��@9�ܹ�$O{�>�P`�����1���T��æK���$Ώ����Uw��=����Ǔ�������tj���Zu���?���	H)v�����W�	%&�P}3F��Ψ2V��o��	���"��K�vዊZ
���C��8�G�? UA��:��o������͘Z[S#�����e�bdO��h:�;�wʂ�������e��	��vZ�$�0�5f^އ9y��HxN!���NB�ũI�fj"�b���A�^/��>��Ҥ�B�͞�f+y��)(E�!�	��h抒G;_Mw�;gQ�.��EҰT�4��*)�rmKL1���e�MP5�\KG7���W����@Gs�
:�v�<���OU�s-�<Af (��E�e���^�$�k�*���cnv
N��LY6�l�8�*�ܛ�\�~����[w�B��_�ɟ�ݗ+[�;<��f@�������E�����D�y�F�WW���)e���m���agoWc
oY��r<��Ҿ���������x�'2���ӎ�^���H��x��y��@�H�V��%������?�M� .|�V:.��^�Jw,�C����%h���Np��!�hmW_gXG��a�Ɋ��R�<0���e%ɝ1j斖q:�.I[+�X�}������:(����!;���8��F�<<$72��v��z��;w�T∜��T*�Rp�{|��"�ל�]�J�
n/�؜6ax�����5PEЯN���;Bz��}Cm�F7���?�YUPp����\�
�.F��B#�D4�J���V����JA�U���"�w%,S_G��(�+��m����@%���p&t[!���y�~�9���1��}��	��C &���e�ܾ�`E@�����9��9���\��Q]
��k�j�a%]VY���}l���Vg�O�d��wjEw+��H�km�x�,�m��kD�$��b��
}\DP�u����^���<�_9n���<[�/_ѹ�t�+	�8혙�V��+���=,C�a�`mc�|J�������"�_�%��.P'\J��c7��9qA9a�t-���t"�ɋ�γx�'v '+�֮��뢛W%��Y�͢opH�4"҉m�@S��p0TI�����t�r���W^[S��p;{�t� ��BJX�9��ۤ<93=����|
���]�=Bw��'
�����܊/>�Rϛ�l�y����駟�����~|��}�QTV�I�q����F�i�+��;t�}�8G�Kad����0�1�!��u2j��I���A�*�}�Z���+�׌���\���!�͜�H�3���0FDl��W�'?��� �7
��R_���F#}��k�����5�X��ה���Z����X]:;t>;69�4����$����3��ڷs���?gB7%�Z�����ik�7ȶט�@@O_���NU���QK�B��뎢��]�M��<���mo���sc�u��ؽ�Yr]Y��Ԅ�9~a�H��H�]0.���*�S�#��cC�ZA�J�M��M/.���m�k7��ܠ�D�0����]�#�PcJ՝��;���"k4�a�@�nE�W��k�DO��W�!�N"����&�7��Ƶ?��t��'�=[��_��� ��\�ܼg΄�=�ص+�\�9��n��%��064���n$D2�07?���]�݄� ��&)wm�o�2�
�c<�;��b��@4�'����6r��(Ր�����C���R2���G@T�⃊'�����!��]�uc}uQ�-���1��jnm��e0;�^(��
vc�zL�Lvܝ3Ry��&�����������&f'>C�`E(w��`B��CԵ��"�A.�C:�ݛoad��L
�l�[똞���e	ˢ��mmMr|�E����]s�K`E4F�v��q���p֔��֦fW�,�>}���+Iϯ�?��Hf~f��x܈�G0viHf��H]���m�������\T��\۔��d��崦,X���5ux��&P�����j�,N��`2�V�;�8?���_�s�@�:\0{*��:��	�"*��A�T�
��x9���5��w/p_B}C�{�8W��P_��������cڕ�2	X̜�S����E$ҟ����A��W�����>P2x��r�钦���ؐ���Z�`O�&�Ħ�W�<���}uuukJDp�X���P�c!Ʉ���	�]��cqq	��Jy���s�Xo��|g}+��a˅Q�})�����w*���&]��R�f�@%&:���hX&*�L2����iu������2B�8�z{��f� V���w]�/T$� kL�H���$��{FKk;&^Oa��D��^A�]eJMy�����wڅ�!ր����F����V�@j-ba�����bhhD��:�"�9'�1���K����qtUa9?�}y���c��@���t�_AK���,G�$ç� hU�dB��=DP�hF�������x��Xg�&g���ƄNЩ�'%�"�Z��➘S&&&v||�Z3z}U}���,�c~~V��c~&Fv����l?z�P������z��vz~ܼySy~��� ~��_��r��5�F�XX^�����Q���C�ܭ�(�*�m��|�iD�%j�7
��	�F�朰���`�ËdQĪ�܇l<���V�U1?7��l�{�Oʣ����I ��7e܎��(��g�E��IY�:d����ۃS)6�NS6�(?GUePxv5��%�Z;���QSQ���w�%�sx���B�$�.�j	ǻAt��E��ge��q�P^�C��)a6�5���-��q�xT�ˣ���ݺ��v��w賅�������'/�7���;P��V�G��Ã�?�������"����1N��89�������چ��zQ�٩���֡�kn�y�B�D&H	���|��ν���!�O:��A��pT�����3�/~���֌L&���l��(�p�������ӱ�8���PeU��t��A�ߣ������������K�i�vadv�o���0��Ԡ1��Q&�����?���hke��p~���+R�<R&.��#Դt#AhV��$n^����&��];�����Ҳ�g�u��=�v��h?t"̞����S�x�V�Sժt�	�P�3��*�D����]�@��� �S3���{*b^O͊�1`Y�K� [W���ƚ:46թS�&t,���L��D���� }q��� 1V�L
Q�*P�{+�x$&���HB�S�ē��:��_>�͛��p�a�V)�׷(�{,v�\�1���:+TŚ�]Qq�dm��q9�F�ޭ�'M�����<�N�~�n1���e���B2��M_o��;\�8P�5���������	�,v�I���.r؁�EH�yA������d�9��ʊj������H���O�&������ޟ:��~��	�h�ōeq[�n�����<&��C'ʝ	��@u�����w���/�(f3�{�=��H3�3Bh�'A<	��s<t=�i���H���z�|���U\װ�d��̎�_k6z:���j�ϯ�o -m���#Q!�R�q�O�`!�ǉ��9��{�!p���Ǣa]�vEw��.�4�������wf����cwN<8��a{�'g1��\6�����_�@,|�	M�`���m}h�B��l���1n_AM�Rr�sˋ�2�3`�pe�u�@sd�DC�ƺqq	�����əy������jQ��Lpo�ݦ!D��Ґƭ���^�v��?8�������h�d�>�k�Y�i����)_&���v��ǧz��0���\˾�M��ܱ?{�#����ǫ�,����0���a���X�|g>�L*��`'m�	�-�Љݰ�v���f������[\�R�(!���e.Z�QH�P]Y��@yV_y%�1��K�x%m9`�i�C�@���"�99�#�9�b�,G&���25+����io1��t��X���3Db4_���;p;5��P7�z�v���wp����j����O�r��_���K�������|~�p��cr�e.��$�p �f�0�7�y�v	}�Pp����_��������{��[ܹ2�:�����oQUQ��C<5%u8rO�Br�"`kt�_�=�
�n��f�E��������I����W㰍���f�Iiӝ��;��r?:��PUШ�ų(����/�ĵk7$�q��#�\n� ܏��������^.���PU]�gϟ��<d��0WT��׿�L4&���1%TJc�d|rr���V���cfqV������:�_~���6\����e2#k��C6�#Aκ׋�Ewo�Pp�>��r`y}/'����(�2G�g�0vtu��u�2}�Z��(
�uSV�,�)���&�u��,���ꊞ}4���W�084�`e5��W�R8]>�] ���ȧ`��jF�����u��������pzx�N���B��?P�N`em]��<�N�ZL
n����&�--���J�>6���5�?�5,yr�i��T��=tum�J�.&�L�o^w��cu���k�W��tc�p���7����v��٩
��&2�lCyyN�w`3�Qp���յ5hk�����_��Ȑ���_=ƍ[�d?�Z��,���S�\9ԗ{�u��d�󱓻}t,���!N�=WI��tV����5���p��%��g?Z��Q"r	
�|�*�V簱�.4
z�/b����Z�d�J�;t*�\�E� ��3)=Yd�|�C�R�ZX^�"�!?�;7F�ӓ�졲����X\Y���~/���h��v4G4mY#�َ��h´��_��q���u�6�&��H�G��&xn�	e^:���6�H���,J�jk��Ѧ�J����ɴ��������{4�"ː�����Bop{+4�'�q}y
��?��]i"����־�s�%� �}�����N��t`~eI|}���Q�ﵷ�GkbU8��~;�L����$���֮�W�8M�����(��K,�_u\%�=}�W�]�������e<�q0�W"�9>��GK}k+qr|��S���I�ziyg���8�`q��SG�x(,:2�0v����j�Q(Cye�wN�a�N$���_���ԡ�r��Y������{�y�5^�H�&Je�
�wѝ�ݫ�WJ\{�}h�� 2q2!�����/?�mݨ����܂&Z����^��I�ye������l6����.�J���A��{\QR�V@�l�]m���H|)"�WV����ޝ{��vU�&~��*���F\����uu��j���O�ⱷo Ss��?��E{{a�μ��gG��$mq�R�lp����|���?��H���ء
������[:���)��Ǫ�roz�������F��bfaV����ɒ�����>T��:�|�T�Z������>�&�ƇD��|1�Ƥ���A�%G%��&��
R3#��nG+G��Uh��j<���)l�������z���̺�F����Y$�����Ȥ@ʊ���9X&>/�!9m`gD�qr-����䠖H	��Ѡs}�G�k�R:;9E}}޾�v�ӯT�W���2��W��I�2}1[��y1v���l�PB�֞)��ի����*�n�?������{�@Y��z�t!#�f P%�W*SP�`g�J�[�`���9)�t�">���:�=~�����[��g�����@�<G$���v��jy��u�˨&e�cc{C*N|Vm�����+�S"-�Ѽf����o:�-�?����!ɛ�I��ǿ��Z}��*ʽB��>4��<U���O5�+�=r��L��`    IDAT�y��6��!ܽ{C��{;�fG��j���,��+ ����^��b���!C ��!g����dɥ��ڀ��^ѷ�n&'�0��L�n]�$D���1~�{G���O?��%U�L���9�8=����>�u�S% ���Q�ł�����Sp`�$�D�Q69���׏%)K�"���Z)ʍO�cm}�UJ�k���X|[.��Ή���������焋I<{����e�K>�j�$�̜���9��I�����p�؏\�3,�V�V2�&8�ד'O�"8��O�5�qtN�u��Ra�;��N�#K�]�*xZZ����k,,.
'Apw��]�|�G'� T�,�����Cq� bKQ���LN������:��Ql��be�:t��Z��������>^��$.u���Ј�.U���j�5\^zg��v��QB�1��ɂ���i�Lgҹt;\8=�+�U�ѽ�mt�����-M��,����3���F�����<�@���$y��N%�J�MuUڟ;��To{gO��0iB�b��p�!g����]���b����8�,��v,�p4��Ʌ�4�)��}��n�d����P�ԋ��C'�cns>�룽�ּ�[B�`��鹦t4�8���
��j��nQ#��Ӈ�PXL���d��(A��Z�ʥ6J�'���}<��Y[��?����1&��Q0��A
��dB��2�\j�4Y]]�@0��P���klIQ�:'��������9�Ml	�#���w��,%`�k��u�����Xa����
�n��E]�|5�?�v�?�m#w&�������|�o�f������ۗ/���QG����\�؉D<��㐺6&t�����
dzf�;�y�6��,/S�N�c!9Y��KU����e���-���҂�nT\�������mo�pV�T�潷1�� A���A<|�5ַw�l��GLtE�H
:�Kƣp��.�/&�/Sg%*�ݩ�G0��������AP�'�������3��y%Ѓ�e�L�G�t�9��$�Kw>2:; �wr&ܺ<��2x�n��^MO����[B�JS=����_!�9�s�7��\�����Ѭ��<ķ��a��U�'�%�/�+�ooI����44����~� ��QQؘ��f�z6�BSc-z��qzr�U����\G	Jщ�v!�#Q)����P�߽Y��7��p�#Cڧz.�+�Lgp5t���s�C�x��/�$tr�١��^WB�@G�Í�E�o_U��.���ر�w(iQvpN�M�r�:�(ڽ�4���v7�9�{sZ
�lk ��ʁ��u,,�kZ�N��m�[7o����h��g[�p������D�����i8I�u�1:|��	��PW�B���,0#ј{(��������2��{���q�0�����+2���C�yI�ZB�R���wm�W�V���)z;�p�Ұ&1�e������K�}������SB�H?y�>��T�d�G������09�L��d��u���Iʃ���ݾv�:>����8�z�&�����l�d&vĤ^�����63<v�bYe�BgSP�4�	����?Dd+%�ϙ酢9ˠ3���ص11ݺ~k��x�zNc�B>���i��c��ؙ$�D��M4	lt����ՋKTM#%)�C�4Î�.�ѹV��#H��hR���V�6p���b.�U�0��]���N^``��2��r����������AyU��[4�D���㜢g�q��V�#gRQ�����m9�QpgucS46�����lkGks���~�\q�SP�;N+�����)bh8:�Y�D8�͚�Ǟ�����y�n$��0Y�H�lh칤���B���$z[jpilG�(L67��U�8W6\��6գ��
���0[��`x�A�v.̯ r3D�� G` ��n%�H3-/('ut�css]��77�195HZV���iA��|�}=�
S�:�	�H=�y�βT��u�Bg8��]����	�ۜr�2\QQ�B�9�<�#1 9�aX@0�����Y\���� N�Yj�a��{�K�4K�\�ox���>+�uM��i�F����F�EBH ���V#v��E찳��e5�0m����EfDf�ｷ7��ιY���N�U��Y�7��~��<�9&�+J����h�'�����:�\����w��w���e�h�9�	ԕ�����bquE�]�#�<�!��2�T}=����9����A�=������֡�~;��漢j��|-��?���:`R���X�e^WU���V8,F�NN��ģa�����3M��PT�_~�:^wA�.o��w6�&�����Ǒ��Q�C���%JK���֮�K���ř�;"�.���� D�Q\_�d�i���-N�n,`g�"WG*��H����������Bu�Mf����DY�uM���{'���f���y1��e����w�P�Jm%U�y��py�xH���cG�ˁ��w���Ɋz���w�q�on�������f�uN��'��kc��")e[Y!		Q'G���n��TH#K/on���U���m(Ю�;Ӊ�y�ae+���dws_��`Z&.,蝃wP�ЅX<[� s��}�9c���;���	�P\R���b��H"lo������OiM
$��/�\:�Հʲ�w4�<�;?�����[�����`w���3�b�z��>?LN/�`"�<�4�zZ�v�_]�t�,n�{��/_����}�N�O�.��[qQ)�[[dx��%��6��*��"����|1�3�2! ���{�qsq�VM��tB�Eo��P�{wǐJ��(�������d���6���I��x�J;qNP�%rRxpE��e�:uYq��NcmJ�,X\X���;�O\m=��g'Ǹ8?Ɲ�����Α�8I��E-C��R��$Fq��no�P�?n^��9���D4�$C���&���M���7o'��'&y*��w�����ڎPA!�����W0�oK�A�2�y���v�S�&7�b����]�"�N	A#�O$[>�@S��������hD��F"bN�3 ���U�ch���7���͉C1::����h��Biu������
z2�O�'���*-t���Q6����N�{p���R24>��ق��s�܉$i����/�"t��=���?0���,,-��ԋh�;KS�X��)A�+�`��}��&��э˛��,�ў&t��#K��g��Dvl�&	��d߭.}���I�,�(�zniuv�3���ae(�ͬ��k:���"}r�RX����
��v�wt|��yY5�q��:������D8*++pvq!�KH���Bm]�N}"����BwFH�k�zV�Yﱼ7
�(�D��p�B��<?����+q�l3�H���|Aw�M�)p��x觿�
���M������S3b4��q"�G!C(��<1�fBkG��2��fț����'��)=1z�:=�����SF���ī��hm�>����kr8�IG4�����[���'�{�ۅ�*퀩�f���·V{5uu��;@cSv�����kJ�n�����r����=X���̗���UD�Ņ%�6[�;0=5��O؉.J��yi	5��iRcZJ/�hLl�x,���bDS���pX]8�_��ҳaA~�C�շ �L�Q��x04���*����Z��N�=��}L%�/����M�oj��ck{Or/e,3#E"�Y��T"��*Â��
4�V���/_�@>x� ނ"��_���(W7��
G�t�(s�bny]����h���Wr-��ܙ��7�V����"k��΢E�MO^�y#�,v��b:G�@��[Bf���b��qXLY�Џw�D����+2�]����*��ئ�i6�޽!���"\n4bvf����Bf4�����ݸ36���3Lͼ���)�%�r�3Z��gA���hQV���$ч�߇��9\�
+�r�����_��#���$�Q����]m(pZ�`aNghhi��ѡ&��.��\��I2��$J��U+�2�ǣ�t����`~�w���e�Jf���&6��`����M����̈́�\����S���/��a��+�4����I\��VV���8:�G�ֵ��Dbi�)X�r$�(!s{�^dS9��}�Ņ9]�z{�QVR���q������H��٣�4�BWe�
]6t�6�w�U4����
�|W*:�hg��MA���	�r7΂_UU�����7Ǆ��W�X��A�~��v曫�X��
�TV#�,09�00��Ս��3�����C���S "����0:�:q��]����ʪ�*j�Dt��ڒW��Mg5d��4���	Օ��E��>������РI��種�GCs3&�����Z1֌fΆ�N�U�E(.t���{;ۺר���?F[G��ة���&w��Yȿ�&:���U�`U�>��:�ֶNlퟫ�W�~[��'�-�\a��N�w����� �B��?g!<�DE�[�y ,�W�7������Q"G��ww��%�>>8<���B+�j�1�2���Ռʊr�x���lW��y,�l��t}��"�bbz�,�C5W2�WA�!���ؓυgvF����!���2�LB7���GH�������;ʮ�ܹ#9*�>!cT�8\x7��S�vTT�!!³��ܹ������;�J=�����~����_�w����S�a�hr�K8��*dVwZ���m()�G�C���J��z��PV\��ʗ��_�Q=$��!��+J$��c�:Ė׷`�ڑ5�O�Df��@KM���	u�wF�PY����V���M�32D����H��n��=����#��߃۷_En�U��m1�dmu]yԍ�b�r�D0lx��R��O"�^͠�i��_�%R��9��h�Mpy���������{y�͋�ǿ���VD�U������~4���a5!����؛��j��>�ß�����ކ��N�bi1��ַ�Qք4�ڌ�tXEIrg������B!h�k�K���U�XEUGn�؅��d*'�)
���:w�#�b���iY=%e�ܶ76QR\���Zu�쮝n� �g�^��ʂN)/SN����0=5�dάx��	��f��n���_��'�Wt��\��{$���.g�>���&�����E4��� ,v+l��3�T����9;N�����	��%�$iٕw�2202
o �߻��Q�r�~�^�s�hk��G=����.�p��L���FCװ���픾��
	�3K8��@U]-��w02<,�;'\�C�Y��/J���ǂ����h��׿z��ivY�-�P�	�`{�&��ؕRA��I����{�B����7�~��G�-������E}C�3zzS��O�{�FE�L�q0q�̀��VTp�g2���ہ�������"�	�����tubz�%�:�p�`r~����Q�ܡ�Ԕ�pzx�d<����6��ˋ���V������ryto��v�����y���5.bVgI5��F�`�2w���K����lv+�7&�����
�k���dY�owub���TJS!����y��D�Hd�&Ҙ��i�� ��_��PN]4��U�"f�|9*���.a67Vp����e%�x������N�?4���m�l� k�#�e�k�F$�ME��R���j!�V{޼hmm;;��r����UQ����=��	S������
�B:(_���#@~�pZRX�|�����y�$�9d�n�5����?��^(�|�K�x��i�R����oqqu�?�L�\0��n~qYJM�d�g�W�"��	`&����(o�\Q^��3r�|�W8�?P�mkiEUu�={���A8

�pĒI$35��8όH�M5U�:l��,�y!:D��/ѹ*+,FmM��x��2Hf+�&�Z�2���WV��b�B<��[��0[ͨ�*E$r��U�;)�d���PRZ.䓵���h����?����ׇ����7���0���9�
�!���;�4��h���hl�B<����E.�&���z����n����	B��|19�
M�uhikU�CHvb���l%r:�67�F�p�c�<�WaA'��h�T8,�*F������K*lL��nO��:a�PLX�jBkC-�������ٹyi�	�TU֩��%�f�m0����u�μ�LYf���E�2gx��g�}���8ژ�+����?ByC�
:#,�.���B{m��Hlno�p�#'��B�"��_�L�����c�V7w�m&��ds	>��GS�o�md�&��hml���lV#�7����K!w<���%,����2�%�S�UȐ��Q��Xt��T�iI�-t~���K�J����ӫ��5I_Js�_7j0���2���GT�#��4�e�N�/Lbe��_)����T�Ñ�v'��@UYѷ}jrJ�+>�XŐ��`$����.g**�Ꮕ��ӗ8&@1Z�\z�hy�����dTA`� !��.�M������B6���mx�z˛��Z�H��fG��9�ΆJD�W�/�-~y����6vw�b����s!���NA+>��W��1#���NK����*����Z~��A,���P�{ku;k3�#C&�mAo�/�;'t1o�����d���a���>��_���5�������XY]�o��gjL8q���������Nk�<�EC��:�ۛ��� 3>F�^^^��������q��������S�*�dȇ��b��W8����&Z�Ӌ��.|��k�X	C�B%Dt���[�����i<������H���n�����єA{w�͌��̾�̈�,~S��}
wq%b�����@K3Fo��@�)��kz��%��|K+�095�}�Ï>���5����Ꮢ?rU�\�a��uF�KϢt��0s9����ť9!��=����/��Ս��+��Yd�뮥� �y�.3���L�z�U��l����O�_h7^\Z�&�u�g�faCD��+ף$cR�ƒHbLV����XЗ�^`q�9�Ƅ�}�,��rִ��~�K:r� �3q�����*��i��s���?8
ϲ̓ ���o�wi����g��Xa��'�N�!���ꠅw�� ���~�+�o�h�`�v�l�Wd.��ֆ/�=�M$��Ά����)���m���y�=��6���5ee�O&����{\W�5��D	Y��J��S���)����!N�/`��PX�ٔ���	�K ����tc��.W�)�ԗy_��ÿ񽞦_�C_K��?����I$���F��sQ8��pL��SVa*�`6�8�������B(�(yN.���%��?v�l'���\׀��6��aM^s���;>G�d���v9���k6�r����1f�Gce9��.d�B=���*�-��܃,wN���!ɤ��CP���)��zqy}�چl��i�ojiEyY���`X����:M�[[��2Ȕ����1Y�|	�\��E�n��#'"�y�,=G��X;t�UȂ�Xp��o����H~I�����@?����t��)�[YV�!͈@&X����6y;���;XZ�A6�&2�݌�"�i4�3�Ο���ou���
A@d;��of�a��Dϟ:u���Dp���TǌUo�p��(|��;�{�:=a���������+�dx�gD�
9����;^T�-JڸǦ��l�Ƅ���'��������,蕍]�����c�V;*K
`��b���"�&j]�N}$��_`hhՕ5��ɘ]^���%�f�|d�C��\Z^$�|�:��cFvmyZ��T_���Қ�/�A�
�&�L��9��`�O	r��t2����{E�������G2� �s�3�����D4�D0��Y����'{���!_X��P"��Ek�r8�\����S*���gR]SW~B�]��j8�3wgtPg.��}B�4�m)	cr'��MY'}�m$�X013��� ±�̜`�E%w���%7+
*cV�=��8��Li��LDă�d����$sD�y�T6��?O�+񢻽]���(t��GX��5!O6;��)<?���Y���x�c6��$�L    IDAT_��a||R{�¢2��FE�ҹ��`+��	�鳓�bv������U\���]M��--��"���/羼�V_~@㬒
LL� ��6�^��J��ʤg�Ϣd�f��	��`�U�q���G�'���5����Y2���[��x5���)�I��*�Cq�]�DbIF��b�P:�� ���<�q�P�b���M�����xW��^T7t�w���aw ���"�?���<V߽�=E.�PAwz+`/�����]d,�|�$�hHa���-����TK�k��ݠ�o5��҇�����$���%���g���V���5@9�IQ��V���Y�%�lP���4���3zW�������˯��u(���V����9xm6:ir$�hL�U0�ƭ��ZrLYC�q�5�j�ěI��<w�n�w��,��h8,N�
/.b�[�ܕ���n�n&9 4@˿YH���_|� ��Lf�-��:_�p��?�M����P��/��?�N��H:g��bM���DP�p�!�ā�{��������2hn�E}u̖��������y�@�.�wR����s�tu���\d%�m`k�T����!��D �لL:�d�6zf� *E,S\!]�jʐ�����Bqf	[�B��Q�I{^�uiZ�����7�������;�y�S��}$;���7�Py�S�Z]U!���H49;����\%��dw��/��9����	9{n�#�J��N&�E���AKc2�
�v��|��?Q�6��B��z��hn��Q��v��1���D�j��:Lr�ӡ=:�wZ���v�4V_Y���Z�����{�z;��ڟK�A�<�S�+Mq����<?V��i��'I̽!'�f|�7Jsh�v>��Y���ҲMk'�`dL<�E<�x܅үfA.��0���2j�L���ފ��9O���{�<F�'��L��e���C��h�]�?��!��CV�ff��1�r�� OPbl�)��4M�b#0k�!��JA�P��H�֜r���q����X�`u��ĩ͐����
�F��f8��c�}�S�ң��I��}'d��|�L�ca|�1���TUV&�����ǧzv,�cY�)�aocN^�v]S0ZJ��� ����cr��E�����+?�1!��^M(d�f��EҖ��W�Ø�	��6vO���<©�T�Ny����l�H��w�p%��d�Si��ބ��C9C�K�(�o�fd�*=S.����T���9�������N���?�Gye���X��n�}~}���MM�,R��prW�cy)F�d�sus���s�܅"��}9;����$�ק2���]P��;(�i�iVdL&0�܎[-�
�af��ɹ����5�r\Z��X���Qc~����U�F��I(T(XF��b��x\L��e��3��b}u�������ߗ�}ffQ�P6Go3�gA�GCmU�n�i>��k�R�<E%�}Q:Iu %�t�$�M�+6�l&y�Q��������9�NO姐��etq �+o�67g�6�m0XPPՊ'���4�$�Q��u�p��եH%R��Z�9�[������W����T��W/^#�ex��J�8����n�j��ݻ(��������E��u�qpx����n�b���H\lr�7rY�>u���� k�,�Lw?QA�\_��$�!L��FI9fT�7�
`�`_(�ֵ$:Z�BcK����eznF���x�(+� ���d���Ǹ�����t�g_|�D2�J�������oԡ��W���O����߹�&��h^�UlNF�RI���RN<�&s��"��d]m�0���d�a?�{�ed�BHvz�-����\�X*,����k�b�2��3f�(Qp1!�t&�pد���eC6AqQ!ƆF�N|�f7���fH��@UE2+�.���g���-�=�|Ado��G���Z�Q���ڸ����
B��k������acgW��T�ڌ6�o/b�%��c8��5����uc����YR+V/s�Kى������h ���x5��xw<D*�T$i8����H������H"[��^�D����/5�A�.�B�4/8~���)	����U�p`u}�W~���X��&#��J�_�����)�NUu5�f��ܷQ��Їd"���z�i��Nkbb��ڨ���j���)ȇD���+l���塃[�t{��X�{�,sI�rA/o�A���8>}xG N�|!_�|)D��;*&<S�@�^Nʩ���L����6�n��1͍��̒��>����$�V{̠'�����pL2/^ �'��'��[�bQx�.X���ޛS��䮨���Ξ�Mܝ*4U� /�H<�g����*��t�wq�4�'V��>U�uʜ_Z��e�.p�j�Ja��0	k6 ᛂ�����/M�$�1g3h�*�cC�aqb#d8==�x`z��!kiy�� �F�����]!��O_��)�M4)�@޺�{�$��w�q����^�W�btt�d9�Y�z�L�l�6���#~|����m�X[�DUe�R~�˟a`pPꔵ�u�.�|����AR=���$���|n�U������3.�-�+��$�6�2�T^D㲰�ST�mAOЛ�Y2���vv��ec�W{��������cJ�"{�q��'&�>>�3(�f$������� v�N;♄�Q�g�@��(��G	a2�̸=2����3�����P3�����JC�J�-���˚�n���1�Z���8�p{03;�����-�y� ����5�Q�ˉ���9+�a��[ĥ8=��	$��sal,����S8��Φ�Jf��VZۉ{}�卸�a��P�ވ��"$)���y�F��'�b���u����!������5"��B������*�A�	��
�Y��ˈ����d�TYU��;w���Vw�a��%9���j4�M��޻�յ�nf�Y�{'����B�˂�C���Q�Z��o{[�P�j��ҹ'B�Ŋ�2���ain�W()�G$���9ql��	A�Y����@E}��������!�*�k�{���î�]��#p��5}��o���g7Y�[7�����"��hL�"$�q'��މO!.�o`��$+p��܀��Z��Ti���ߓl�:���m�e�E��{���rtv���w���
�n`~iSz�"��$x��`H3:π�FT�V� �}������S8,�����82f��y�4ʊ�Q����p_ݥ��=N���/��RR@�QB��!,̗�ݳ9!�˜P����"ᐬ�:{�t���	�cA1bj�+��#vs��.�,���·?VA���9�n��Mg:�GOC�2uO�/���0$s�ڜ�G�*��ݒ��RQyyo\���6FҔ`�8~�N��PS���R�9���齅��H��8>:@yY�.m���Fԁp;/cBDT�,-Fks=��6�Cm(ճ����B6:�MY���TI]�D
��hok���b��G�(/.Aeu���^OO�#\[�4*-lyf�D��Ɣ}3��/�v�dx8ҏ���AxΈ�Bxtw�}^�U1��^���YWY*�9�� ϯ��dw�F�sfA
�DC�T���ݽ]y3�l��B� ��L�I~|ֹ���p"��Nx�ܒl"�Φ*�v�(�������T�<�:��Y<wlJ)�����L���-���.6 7>5f��Kd��}���5����������R�aA�IFů�F�h�(��ۃ�H��K5Y�̼�����x-�[\��أ���
�|��L�.��&��ъt����DcR����f�� �K�%Y~�V�:��a�ٰp��9��v�JDi7+����^��Ŕ��*�aqy�������ںB^��wBH��m���g3�\_��~y~*������,��%�8����>��^#pu�<lp�'���&����؆��.5Q��ή�f�-�EUE���Y���N)S��H�~_�dƹ?��S+H��gԐ����i�l"���EQM`Dk{k+z��`���h���>�旵�"��Ƅ��wSq�Kde�Ƒ���VQ]���r��ۏPRZ&�`�o�ٻ�og��7�����X.��k�6;��cB��'�4�.cJ�ZSGSfT6��w���/����6��#�hk�F.�VA�>��:�Ϗ+/6#\�LM��.)�d�M4�Wogq�HV(9�r �%���Z�ۆH��[���U�ags[���}���zj{�H�P�oR��x�B�]N�Te�����,f�e�`ay�K+�R_73�CXZ_C�?7-�9�U׈���nA9��p9�2Ժ�>�������װ����5Դ����Itwv������������QG��_[�箢5�����e-�6��De���2�q{p�Ņ�������'*�4IG#�~��4��n	����k04<���R&le��y��5UhiiB(z���R,�ncfq�f\g�v����/O��ڊ��6M�ggp8��6��!���>�R�"ނb���
�l��hF�҇'��������E��%�LM���B����p'�d���LF~Ȝf�)��8��1~���QdR�X�r)�u���g_�Õ��/�@�Y�	��4˅�t�f�hB�-,���*�/��>�&�~��`_=}���^�גQn��+[r�cA�lm`�u�P ���Rш���$9��;[8<>G�H������HpS�A:���*�7���Ņ^��*����"D�â��%��s�ʳ���ц�B�d#�H�K�zQ����҉7��!
z0`����Y��1��h��|��7���6��I���c��G/?/���y86*	
w�,��'�`�����Y��n�~����SX���� hp�!��u@�,V�O�������P]���3.��m0���3;�B�=����٨�n����0[�HX\_W�Hqq�H7�b#�)T3E&>5��~�$eϿ�J	d�Т���:{��}$NC:����ake�\P=�H������7I&�Y�[_^���*��8������@/*+J��FKѹ�e\^�����n,n�aneW�y,0l�l��9=ȓj6�� �pv|�U	^ޢrԷ�(����
6�K4!w���l��mݝmj�7vPYQ�tֈ}�"6ج�K�j-�\l�4�"I�bn��qIvw�=DN�y����I_��>H%���Z���x�XF�����9��>yPzsG~�����_����[<FMU�Ѹ>:���4�I���G1�nQr^��8|C(��a2�k�)�ٲH�B�I1Y��L(r�02|[ϛ�����G:��&�'YЍ��F��a2�tkG�d�Kk(𖡩�E�g秸=2*� ��>>o��TW�j���Vv�V�6��P'��&ȝ}}�H ����"����7u����PTR�\2��m�.�����p����Wو��7��*����Y}?�ap][�j���d�ԏ3�����{u"\���c7���8��ш¨���[^�����,Tl�e���h��;?C*rq����J���O�ܿ����v�����%�F>Cr6x}��@DY #_��Ȼ2��,T�4�:�*˼(*����˟c�� ��B��Y�U;��©�����Fz��ڂ����������Y���L����>�� m��b��1Y�(������ڵZrY������^��虩Y�1�SX��?�ׯ_���Y�l�^/�7������]zG#�����Û��Ļ�Y�Y,
��)pKz��ddCW���.rS��F��i�ɴ�P�0�z�L�\GG;
�^,/,jo.+���&I�dHr��!��$��88�Ӂ�^$	I�SYݠc ���3d�8�Y���+�w$[S�0���=�,��Д�c�Vn�jC:�;���l���?��Hfo��3굯�O�_�4�&Y�OUг6����ca��~�S(&�ɜ�`��GyA=z�ٹ%�Xb�!�I��ewI? ^"�N�A���П=v�.(��}7��EJ�m��ID��(��R|-Me�����ỾP6��`DK[*k�brR�]2=ˋ\�����*����Ņ�#>EA}�9�0�"���Z<�7�g�Ɖ2�_-�/^��gCEI�sy0>����3m]��C�!lY]V�,��w���Y�ݑ'�P�	u�D��ל9Ϻ����a��d����3!>�C�(��×/^ F�n�(ɗ�`�.op:���������d.�|X��k�$S�������ڤ�Z����^"��itS��G��PAg�9�Ae�?E*�w��C݋W�E]u�
���*Nή�ɓ`EV���ъ��3�
�%=d3�F�r)�dS,t)���]���.��hkk�_X�Q~��-�)�#m�g$\�02ҋp�&#�D/N��sk/''a�K���g����jR��Z���]�ln �L(����'O�`�� ��{:7�_���N��T8o�c��YX���������K�0��)�;�����rxgD��SY����huł�P�`��u �k�R�x\B����� �OJjWU]��Ϋ�3�/-���
�eUR�d%#� �`gJ�X�V#
�v5C�秚�;{�U4��Oa��UXXY��^�-n��d�0�{��A���DEi��wN��u���S#ɂn1�TЗg�Þ�����=kr����=��֋ k��#����0e�����Ɇ���@i�K�["O_�����Uk_�� ����[@�h ��4���ߜ�9U��A�J.%��G)	��HEE9��$���iB��!�v�u�e�=؇H0�������� �mY�ݹ� &���Gy���G4?
j����ޜ�;F��` Í�C��P�q���
�E.8]&�o,`qc	F[##�����6eE�߹=HR��-�/O|���Gʙ~/���Տu�B_{;gf�"˝u_W?��A�\�Djc�xWK�+������9�mlhV1�x�?���yB�\6��8�/�mvϐ���H�½zsS�X��X��U�yK�ѱl��� �G���ί(�F�h�Gm���c~��*����.���;��qzt,�8�|dr�.�*a(~)�&�;Z��ޖ���)M���ё�`���_o�&ty�����9ބːo8��e��3��q�<8�YT�ᓏh�m�E�4?�x.-��\<���T����d�J�CmV������	�;tzC�;��o��;(�8�p��@|i���6k�!���x6>�ˋ�It��Â�b�׭�S7\��i?TY� ��p��Bi��ߒ_��IQ�dJ��s�g(p��/g�M�015��!�Mpٲx���p��@�Ml��������162�hJ��=����u��iJ��R/'&124��86&߭bq�LE�盐{2r���'��@������wu��n�V�~�p4!��YYe^�I����,V�%N�$�y�M[d"B������&�\��ݱB��4!�f�x���I���
�eH2�b�w@V0	M�x�L/*���č��cl.��xwY�,��df[�
�7:�%�C�݆�~x�dX����!f߽�,m79a�Ntai'�����C�9��t�?}�
���ǥ�Ѕ��m�M�߿�u�i��s��.-Bks366�ffF�)r^x�q�J��b� x�ft���3Y��� M��`amS)���Ɍm}��"ٞ2�f�zZ[1�敞�!�����nx��.�@6���,O}��Ց�_0X���� �o
:��κ&�D"�����L����nk](?o&��j�>6L#����;��]�/C���d���K^4��Î�V��������d~�G���Y�M��!tHM)��������:1��P�!��n"B3���zJ�@"�J�*I�0ӦI��nSSS���H�(/�@cK+��δZ���7��1��sM�`�#��[;�;p����di6�O�����!kjc���.z��S��bl2?���-tz�Sqp�ë�wj��L��a~n���&"��ţ�$���G~���l����v���I�nR�(,� ��V���~�tuau{K�WU.=    IDAT�J�#g���Z�������$#�t������L2%'˭�C�p�TS�xsu�ã-Dc7p�3 I�F�S�ȉ,ʋf�s����QO����_��4����;l0�n$�1��)��5����7�TH�7���ƭ�~	��������!�gO�H&����@oe��g_��b�*��[X��CJ��v�$�D �FC]���pzr(����Cu��$+�C8:9��~"i��ʺ�_Bd�rB7��M��!0�YD�z�I�aZ^�,�<4lF�j�Х��#�p5ٌ���zRG�$PK>��z���E\���dn#b����[���+���gz:�������)�V�;˂n`A������GiI��@ڈ��	�H�]�t���B��bg}�&�����X^[���>��cD�A�l~���斖��{����h�jBbD#t۽��X`6Q瞖��id<���{�d���ĝT:OR�r8�b{\6tBƱHDY�΂��Z�Âb���<���[u��t*F~Gz4AH߂\"�͈6\җ��)K(��ݑ�5��X��sD}E~7h��01�/�L�Bu@>驥��G��矫 ��G���Ҽ�ݽ����a��=���-,J����Râ��n�J��0�u��b�C� �ݮ�N��Օ/O�2���������C����A���A����8�𡤼
�PRDT���AA�+s��Cwڌ�����[�%��cZAk���}()����&ycc�z:�T[-(�l�)Z������0e�S�?���7�L5��3@*�Ю�}��<D6���Ңv��~i�S^��{t�����e�L~�W�����������Btw6���+��h�oBG{/��(��aw�ecLĀ�l2��4C��,��<y|g�'ZϱI()*��gD�Y,.o�g21���=�?��g�`����>J�)�FP][\��c�aL'$-��;���<>�?&u	׀��f"��;÷��R�c��?��S�J�csG�y?���f����//-h�c��I؎�����-�m��3�E9�*<�5%�����VS}��}�-��'����UFk>G�����T'dR��1*�]��PT������m��ckg[Dh�9��w/���+�,��a"���DY]����)�����=�l�]�h�.A�	�o߭���L�2tN�dpB����� �f2m���%f�W%f�9��9ݓ��M��Y�$�:Z�T��hHŔ�86C��w��q$�h�Ld���HE��lnD{s�.�0>�VFi�X'�pY�q��0WClB��TE�b`�A�5���:$ѐ��J<}9���ϝr��:3&`2g������d�v�2����	��`�{���mM�~B�s����'2��L�T�,��܊��fA|d�'�I�Y$��]�T��!i�RWQ)����	Vu�������J �_x����JjFh̆��}�l��E�!-܉Qo[W[���B̼���=a`E�"��3&W���S/3���f�Vb����=��l�id)��W:�̔�ݢ���W>T�p��f1v��;{݂����<]ZOWKNqys�O(2ؤg�[WA��E�DR�����0z*U��gL'�r������ R� ��qrq���bL�����5�2�����5��am�s+[*��c�`�R�_e�S�ƑM�q��~.��iY]^���>��GQPR������p�;���^j�4�A?*J��O���]<��,8��.;"A:Ĺa5Y�Wgb?'/6|��'�� �`�9`a@Ky�]n�<ʚ�����Y��W�7=k+|_�[5�s푉G`�$Q_S�{wie����[q/>����0�W���x��C���(Ҏ�ɋ7�X�9��Q(�!��\6|��c�~���as���X���:M��uOL�A �PA����.��:&2F�����{,Y�ɄN��mNx�K$9:��7��=���]��OF2]�_K%�٨�� �-�5�+��� �W7�!��݀p�ǻ��Xz��)�y��Զ����b��+�F�Ubh��T;{ۊm��hEe�W��|7|��"<���x19+�T�&0���\���C}=���/�����nGkS=f�g16�H��S�3�%/�2�l&�Z�u���Ŀ TI��S���!��x��K���D7RZI1����Yg��`�ZѰ�T���"XZ��?g4�q���w�D:~#5A,����mAg'�e�6'>z�P�1凌�i�?zxW�3���^�y�"�`l�LB<�s_ogVJ�i�ͮ)����������X��Ӫ�Nx����!�4�x0����k50����O.��|b�IrSz����cw�ȹlko&�fʩ"����g�9�FZN$� ���_
�1[4}��� ��+8:9V�y"z���g�]�D�ӄD(��N�{us߷�����
�,�Z*�PY$r,����k�?<£;#J�㚆k����*�5�j�sF.|�ZXD,�����.�l@ecJ������CN�ee�"L����iwɆ9ǘҜ	6�#l���	5��__YV�
5���h���f��6����Ҋʼ�i&%~Umu5:ۛ��̈́�D�VGg�ӅǏ?�����~N�݂�c���QT����^�L#ER��q�XM�.r���������m��B�OWO��?��x�J�(g��cd¨�xQQT"�i��@���X{��b�q/@!�B_w'z���n����K�x5��DD����1E�h���Ļ�5l� ��K/x�h�A���i��̔$'�|z�{E`��pau�<�VT����������"��ry�B4@.����c;�d�_Qw~y-#�p("�4��h$�n��̔{�dVSY�����WW�ņ|��c��`��U3�%ǂq�o/�hm���9h�A��W)��@�\�g�Rw˼o#/�,B;��11��g�x��>���ׁk�������!���|an}��{�yJp�
"e�'<D8p�wo&�Gf~gw��z���\�RCA?����lm��1�}.�c7h���.ۈ(���kB�kj�e�Nf��]���2���b�~�o�L�� w�����5���D�����]�I��d)��c�`m~{k�ȥb�H�c8�н�Q\�$�����͌H�Z)^==�������:��չ�{�G���ۉ��5�vO�v�sk�0ڼڡ[mF8�����}B0(:;?�w>�Օe�};#s6�>��c<{�\�r����P �a���=V]�� �N��H�S������2����	��b���$�*�e6�Uu���_a���ee� �P�
ק���z���jD6mD�X���OQ�ܭ����
<<zp�������ꊠ�[-HD#�Z�X\^�?Q��ݘ'GE3�����f�
�ኋv���5>��L�f�g��ю��MzTL�55���$,6F����O�F�Y��i����*�
�ـh�e�N\]�*��ns��*,����E�K��;�We)P�e6
IˤS���P^Z�PЏH0���Z�o�ʘ�:<r=c�m��qv��噯�����F*m��U��{���QZ`��M'�dF��dj!�k���Қ��I���_�b4�Ƿ
���'2x�b
�Ta�`��GbJ�jolF'�/1<<���"����?��@����5������_�x���Uc�¢��HP���p��BH���#��CGC&<��ǈ��� m/����ܨ���ى�c6O�F���>�sO%c�$o����8ؘ�۔֐�����)���6�+��焞���р{����O�jc�[��b����}O����32��j��U���{��_ے�.�l⸶ Ɍ�R�|���P�ӣ�����'����߯�]� !�R*(�T!3������
�|�L���'j�y�����-�1�(����nyUP�ƵEoO':Z[0?7+�^��8�p5x�V�
:w�M(,���k��|d�W!��x��Ɍ�Ŧ������¹����=㿡��6��?���: �0�3�y�ʫe~q0,�#;���.ܻ}�`���bѐ�#Z�q���T"���6x��x�f�f0|{Tv��XnW�V���O�t�,��X�In�Z_UAoh�S'\R^�t&��m����&���s�n�"g���;��؜ڧ�� $�BCk�����M��}�yH+�k4��L^�������_wd���<����
�>Z`:���I<�]������m��:�I����#�(����I��e2��iǝ�~���N�ɇ�n0*u���/_>GGS��%��l�����T�<�]��>�7W�x;�奅�Y-:�.�G������PV^���g����$!w���oK�c�������.�L*O�K�qvr*?�Al���"S�ϊ����Ԡ777���H�26t����R�?��M��l�efLy�o�>?!ȝ��g��cO����/D�� �!�h�F�XyUe��b�a���#Ol�D����ނ��:e�^���Q &{�j�l�hP��镊_�[�0�B��uX^YÛ�y��~�_��ȁ{G��<L�3e���6#��
%[��HJ�2�.,"g���r��Gڝ����D���Φ�@$3}�䉌e������>�@o/&^Ob���No1����-r"`�y�yc6,�0�k�;�h�RA�͞3��yrQtu��od7�9��v����aܡ[���]�A��!�Fc��L���D��5!f�j]#�F���8���u�h�3:��]N�{�[�dM>��w�6������Vw��Q\D`H�k.�#�;
`��qxt�K�w�Jzn#�:�1�/��]�i�J���҄��S�ל^�K�PS׈��=%3r��N�p�C��K�/�W�ѕ�͂����K<��($�H�����u
o:>����<F�{	�U<_���1��l�$*��r6��A�0ک��Y�������!�d�ÂJB0��WW"s�!���&,B�00`(+} �q8,4���D*�E�\N���k���3N��t�1��h�æ��2 �Y��d3\��ק�}wuJ:�\"�,��MnT5�B�Q�5����&ǥ���}�:/���n�j�����ß��Wo)u�RAg���U���c�����Wԣse���Itwr�ⲉ��N��y�=|�����U���T�6�u� f���A$���SÕ�%�(������'����
�N�l*e�M����'�*��B R�QC����ݝ}�V8�V��bcs�U%&�x>9�$Yt�p"�����n������6���''n��0�ɚhkz���DR���DMuj+ԡ�5Us��J�-�TJ�������[=�pZ��s��	�����j�P	1��[VAO�?���w�yz��T�� H�`&�sw����43����k�=���$�?��`����gd˲d�Y�	����9'� I�*Tλ���b�����4�$
U��}�p����7�q���R)c������V?��&�'��Ԅ����מ��;�-ڙP� M�"ꌵ��!�^>��tqCA��ӗ�_j'v�u�n���\���Y&7�Μ*������}�H��3h��PH�ӫS�����Wf���\�bm�F��?�hװ�t`i$\�'�3/��d�K�fA���'?�@���Jr�n^�j�v찭[6��0���dB�{2Wb��γ�O���=���Ѡ?vTz#���ҳ�����п����+״�c������662�DR�m_�`�k�j`o:z��{zev��"P>�
W5���m[���Cv��!;���8��#���]c�����yO>�n!o�).U��mv�Y��[ݠ��+�y�YҎ�3������S��L�P�o2~܇�����~�@�v��={��D�d�;=�O>8eS/�.3U��{���H5����v��Kb5S<}�:����Y:�n�Dס��6��GG{�����;}g�����0B�Eb*,Y�@��Z��|����,�ûw�đ�KAƓ�v
u7_�2(:v�,��N	}i��U�o5C�����z��WJ�A�$�Ǌ�u�h����4����C���ǂ��E��y��P�?<��N!W����Ɯ��el5ۺ�[jp�/_�r�l�pD��nCv��m��,-��ǟ}��IT����U���ŖG���)X,�C��]�M��L�@�x�@��DA�9����+*ș��C�L3	�{�|����ﷅ�{�j��.�����7l��c{��Hq�ku��Z6��S�X������[!~��+Y����w����]X�W��o�u��8����wX$��{F$x��r����[2_�Z�ge�0-jk�����%V/��ymǞ�����H�,��f-�9~BB&S�o�V	ZGQ !���mV��9V�z�u$ԗ����@FN��HBD�"���E��b��w���n��ȘM�\��XȚϲv���J��=t����!�	gn��X���3�����Aw<���<Z��:��ʍ�r�۽u��^����Yu����t��h�`�>���%&_<�SǏ[6�V�=�����k��>�1�� 5(�Vk��T%1ˎSq�����B9�j���@ݒ��^�H�0م���'�wu$�7/4��F�`&���	U%Z�b���E������̪��xQ�F;[�Z�}~�������ܡ�������?������~��T�$�����'�"�n<l�,��)|�W���ƂD��=/������u��mld����:++K�Og��?k_7�=�Wof�jq�j����!S�H����5��ܽþ<���{�V^�G���w�1�z�,��(@�� ��^'�F�A�����&v2�p$(�����Z�Y�--/*�3˦���:>T蚨 ��N�x��*������_�e���M=�m�o���񞺶���k�[O��3� �a���=Q����&��vH����&����svd����:҈�o�O�˙��Q��]��\�N���675!�m�P�WW�R��+�ڕ�'�;t�=�����5n�FrE�U4��epPb���b�;����@�Q��*ǶmWe��7B&�u���?W����`�N{��h�d�W׭��[6�?yj������u{����73��C�v��Ϭ�w�ֲe��%�/�O����Y,����c�}����4,���o���c�wt��H0�^�mX��<�O����}~�#%t����.۾�b���Z�q;wndD���~h�.~#�='��!HH��KYV��E'(���8,I�K׮����:�Q���ոg`pP������Y��o�<���H(h=���a`ӝ=z6�y$H�U�[x��߽bar�Z'9���A�$t�A�V��`�
Ļ��ߦ�^��#�m�Рy$��S1�h��O��^�*U�ٹK7,�sJ~�@�R�+�o�6Iz~��/�9iI$l��ذ�����e�
s�B�b����>o�T
�*	{����6:�٦�L��浹�w6�jF�Ό�p�c�
��Ω��#�[Ż������ߛ{����_�Hz�qe�ޢ-�~l�n��jnE
��Z�"m�6.��1Kc+M��� ����:��������1�������Z��=6d�t�"-����aw����\�ʞ�Eba���"n���W�����;|���w�����~r���E	�$�0H�s�Ob	Lmfۉ֨�f[�9����m��k)doQ��!纷�Gn{�Ss��٣]k����+I��Һ-,0�+�C�
v��W���MqF@vP����=����;	j}e���c�n���wD:���*������+7�����ǶZ��h���_�˷��Ԋ-�S&��o�ɓ��έ�zjR��}z����O��;0(��;����5�9D*(|�Қ/@�`V� �Yg��D9ףVv.||������a�����5��ĺi�VS��8�G
����Vf�kv��m[�f�
���⾚u��}~l��~z��oN����֟��/��J���l�.U��N���;g?��@�ӻ����lcͪ�}a+1.����"
Q����U1^�;�e�I��\p���B��kwڛ�y�+3K�Aeg���}��n����
"�n��g��e[^^�pږn    IDAT����\� &:��*}�TZ�*V<�+�O����j�3yaᝠv>#p����ڔ�Ixt�@�n
���*�k�9{��%�}�: s�o�o��_Z=�,��^�4_k����-��o�"��q�����'��^�0u[b�>���:<hu_ծ~s�N>h݉v�Ƒ���았�OP,+t�?��c{��M>{$	ݶ�xC{<nkkI���3S�yd?���K�}�ּX�b�I�Wc���0
��B�}��&ɜ`�}J��n���XĶm���zr��-8���!���?'�`�Xʧ,dE���'���y"��,ڹ��O��h��<r�bF�#az�B��C�)[<��xĆ�6��yx��m�l��b�S+���G�bz�|�v�m��w��{gmvj�&��Pw�+�mdtH�N�Kk637�����;t`�]�􍭬�$!Y�F��a�c�]Y��۟"�����6�6�f��̔���1'� <@ÿ��j�k?95e�m-Z�۹cLɒ����c6��,l�3��F<��<g3�Omq���rKٻ�k$�M���*|��W��2X��p�_z��;w��;-D�W��Ru#�UB��r���re�x�$`=���rz}���a��v�����?|Xֹ$����O��6�`�0Z:��Ŧ�e��b��g��θvI�'�h0j7��uk��,A�Z�J�$�6H���x��_H{�5M��Ǐ����Xk��9v��l��C{|�y�)I��D;�؞#X��v�(ŷ��dۊ�?r���E�\�ث׳*��ݦ��t� ��+�^Z	ϊ�F![]y'?����Ą��(Rqr$���|w��V�`��P�HҘ�V���߇�k��ﷷ�sJJ4	 ��mdۘ��(�I2����S��翶8+����2ļ�7�k�|��1i�?z��֒i�T��G+�%Z��׾���;Jq�zX�{��NB�aٶΈ�o����?fO�cϞة����!�W�]�"E�C��$r
�ljn�n=~a5�O�zp(n��vwڍ�����Il��j̰7]]Y�����a{=7gV��I	��D��g2"<b���f�d6;?oAܡ���QO��3-/���
��;\N��$BEl��b�>�B�l=]]�D$*6?��Ba�m�r�+�ݘV\&���<�)�����?�������3����p�/����T+���{<跷`��X!��f��-��Ν{mǶ]���嗅�q�t@�"���p1r9�$���d�pc#c'O���R.�"�ƕ[,�O�/�*��N���^�ЁD���b�d=�����VmWg�}��Y�p劼ms5�==bs�uuK��^�n�D}�/e��z�n.��D9 �|��O�Ee
��CFBg���T�XU�${�r/���]����[ZSB�I+��S��C��J� ���AR��G0qMJ[K�����P$d�K��ُ�'�2YA�����U��Kp ~��Y{3��ݽ)q��*y��Nמ��:�CY`�`P�Rx�=����-�I������)[Y[�=�C
��
��#�� �F	,[upؿ���d�|I���zR�=mO)mw�}m/�_��7(A��x׈�9���;��P�oኌ0������Ke\���-T��#b����^��=;ml��=%���G/���9�Y�����v��1�ս�Lѩ�7�˖��mv��پ��鬽]^����X��ծ߼��xG��K&x.
r�-=2���&��'�@�^����?�Y{��YK[�:���ӂ�򙴂}'t��޽u�	�*<�������}�ĞܻjQoN�m�<ҹ��Џ���V�b8�]oV�+��aGU܏0֑=���S��΄ݺu��RI;}��I�+�]���R���w�%ٹst�z;�v��E�k:R����>{���$��������v��M+U}�Ε5G ����槬�1��n������wf�/�o,&ȝ���)�*�g�;v�RB'qFe:��T7W(�mzvA�;��J�^?�c/\�zi]]n��׹�y��m�eI�'�{g��a����a�g���v���3���r�kl�:���ثX�o�M�����lnC�<��`�l�O�Z�����]�Ĉ�d:���w˶��l�=���+��X�Yr0,	�
I)��α�Z����Q������kieu�iSHv��Sfgg԰�l����5>z�\�JUki����c�]��M=�i���f�t��{��(�3C�P2�H�^�LrͶ�w۾��,������;-:+̵��pY瞄������y��*g�@((2/�&��̼�A��f�Q��Hf��]���f-�.����z��i �7������[c�1������1���%yu�R��l��T*E�zdA�߯��;��P_.Ś�@�Ċ�OY���h=4��nڒh�l�-���=���]��	��~q����j?N�JԹr+k6��Q���+�w챁�!���)�
4��i�z]ںRȪV�cW,�Q�E�1it������n�o޳��_(�KԄrO���+���KU�;zBU��Ĥ<r���t����+u��y��*�����ޟ?h?b�L�޼��lљaط��b���� �GŅ���I��{n����jRUWG���r��0`a����D��^=��Ǘ�
+��;��]2m;�ۑ�O	}=���9Z�0K�1qp�li��p9�N(W%�����Û�T�p�П���*II3��V�N)����O;���Ҳ<�}5�VX6o��MCv��-�CFbm�L�������c��S*��[7��ˊ-�38h_]8/�H��t���Q@ù���^����S�Q��C]�Z�+���C���j�.���ա��y��[{���cY(��re��APc�)�`��Wp�#�[U��M=>O�����u��4�x�f�5�yH�[����}�����G?��=|t�&_<����������W���?������y�����8Ε�����3�Y_��������7n_��*x~�����1����m"~�_�܁��ٽ��ݽyC���-��(��[^c��g�@UZ�o����(�e�^B�w�'J�t�� ��5�ǀ�ynA��B�⁠�=f����7��A�Sǭ^�P!��-	�L窖+2�X�[���6�=��._:�:���=!ao_��|�L���n����]�v͢-�{-��:/�̆�c~��o�|1p��\�u;����꘻��U0@�D$��]&�f�g9��1�H����n9i�mQ}�On؋�ߨCW!YXK���QH��ڐ�CȦ���G�S4�o���^شɺ�z%����aw�H�mp�{>��.�zf�
r�}<ⷣ��J������y$�k|��
��.!he��	Gbv���pCB���
ҹ�Ժ��A<�&w��c��?S"ޱs�����[������B��~	A5@B) �e�4E&���w��������A<�u� w:�8�Y@ٞ!�������[c��=���cD�E��{��mG�1�
dnrf����S#�~)|J���.�˗O���d-�� ��>8�����'r��>&-�Id����>�/eJ��������7��h��OB'G|i�C(39����9����P���F�1���~�����[N'�sS�-&Wm��ak�E-��,V���4�\�fE��nB�o?���?���G/�ք��~�������{^��oۮNpN���7�ض�c�b��y;��B��yA˳o��Y��%�Q�R6/����NAe@�����MC����;v��3E�Z[aV	Y��f_�VG	C{qqI�7CCC��X���;z����+�,�\�I���<;/��nfV�`�UM�>x,+�O?�D75*-	������{���N�:%���I���!uf�\�$�L�d�3����V�.[�ϊM��2yk��b����T�R�5�qAcW�S$�dv"�X����L���ul��V���餽���"��x�өs��7agN��׿�Ut�?9+��H���Ç����߳��5����[z��&�0A�W�ƽ`T�E�ɳ�{��Y�C""���٠ b�����`!#,�rⅠO��U^^KK�T������m��c)�A`��m����>�Hǀe
u�Hx>DfpE+)ز��Q�PI��/$+qQk��� �{�g_�����.4�����E	�N|�}�v������ػ��_�d�ָ�ݻwŭ��0�y�-b@��}�V��@O�*���S*I�s�o��tI�?
�V�g��D������|d���eS)��g��˗�b`Gc�v�+�^���.���#{��k��-���wؾc?���q[$�|�}/W��E���N7J^$fB:�a�&W-�g)�mtt�>��+�R�N�����������0�Tx�����=������۳o�`{�ko��x�\�����x����uX��S�k�=��G��k��6]��E¬{����[B��|�:pP�o�޽*� |�lf>J��1��8#X.w�I�I�r=oOn������$�R6Z{Fml�	�۲��A+I�@�O"�e\��w��{�������3��?���OQY|�z�~��em�@�Bx	&���;�=��W��^�X�ڑ�8�?�؇��=��b�bWoܑ�H�|
��{�h�K��ƀׂ�bjJ�>q���W�~�ײ��m��z��t��֌��	�C`"q��_S�T���`W/������tR	R	��Dﰄp�!�a�B�юQP�l�tF(ީc�lh�_1��y��%k�F���1�ϣј��gW�?�b�.R��)k M��drնoiHv��9��ƍ���<y:�.%��ϧ>N�vlӸ����a5C���oX����x d��}B �Z�[�ƺ�B���ݽ�����Ƕ�ڰ(hA֭V�U���bm:i{v���ڒ]�z�|���I�@H���z������'����	�Ͽ�=��|�'�@�A���&������J�wd�@6?�l]����rCC����{�8���k�#]U>�� ��k�u3]�zM��$
�؇���y�����D�s�����҅�ldt�m�aw�=�Q=֔�h�*/*u
�b6m��e�2�'b]|~~Y���Q������qP�s���K���|�_��mݲ����a��J�����ƽ����WK�^Y���Ƕ��U`2#%�ۻL��#v��ߵ`�˒ɒ�|n7���:F(�
"*�D'Ұr��!	�k�H��7�)�6�9�V0�	JX�n�V���ON[!���/���>�D9_�_��K1�Y�{p���Ƭ���Ç Al������/.�:�aٌ����M:��,��ג� �g��p��Ʉ�I�~`�f��Dm!� ��]9���z��@Udò,ֻ��?k�ĀD��V��_��T��#�5������D�o��T�j��V���w�����֘���[�l�62*H5��;i���w�L���?��z�x�m���)��*E7F>OUs�<ҭ敻 D< ®�v�=aM�R�(iS�ۺ�я\e��u����cIu2�o��d[Gv����] u���g�l���S"3*����g6�m���"b�|e���%�k�)����6-AĂx�I
�r��fKtu
5�p񊽘��(!"��;|p\F<w�ޒ�6�����:pp��ܾ/і#�NJ����$�%�)D�JŬu����@��^8�t�[��������ol��]����$�p4jV��nyI[�h\�8Ik�(!�f6r�bj������mٍE���k���Y��`�BV���?���{G-��X8��+��\��s.[�\V�]���V@��6�)h���=��~�β|�z]�.<����vٝ�7�RK��p��}��|�A�R?~����鹷�ZX�lh�D*u��uĢr�{��P�\� )�*��.�[<�0��Z�a�d��󉩆���Rk����S|�'�)$Z_(f�|M�^��rnMkkSOnY�S��;g)_���A;x�c��٬�LC@D~*����YG�3��3�� �޹yK���n*� �-��onܒ,�K["!��4��}��0.�;��#�^f����FL=6��o�)��h��Q����)0Z� �����1�|�Z�W��u�۵֗�钿:v���	��miv޺�:��>��R�?v\��ք�Z�]m6<��b�]�q�n�O��	�Y\߬j�Gg�������_\������W�W.��2o�c[�{�n3=����ߚU��k�^�����e�F:miqU��
=0�Y� �zCV��6��kqh�gp��gT���]Z[��90P�ZQ����H`�
R_Y^t�,V������;v�w�v��ck��t1���!�Wn�[��E
d��%uJt>�m]63���ݑ�kn�2��bPI�C�x��I�n�%����-���mǮ=�yl�=��K|YkT�Z�f_<���W�����L;sE�ٺ�N~�9e�����JƵ����9FVw�\t�#V�H|h-g�k���Z�7�)��&X�%�������3��d�:G���97;/�ۃ��������&�s���)���~��0�jOX������s��~�0�+�H8װ��[vm}�<�c?���I;��z��_N^���-���w3v�ү-�4k~/���#�3d>��ź��@�ÈBB�.i�̿�����u�H�ͤ�_7I٢��%�1�����c�a�ݻ�[<�7�����[�_n����X4�f_^8�y9�|����S����shS���1���!]	B_�!듏?����k���}2!�|1��Q'F�K!���o.��ꚍl�m��=���k[]]6?+~����m��M��G���D�?�=�r�U��=>+ϫ[w�ѦR��~�9����Z.��
�Š�ok��l}u�Z[�3s���ƶٱ���g?���!g�~hk+n��"���۶sǸv�����ȅ��q�CF����;��y�ضQ1��EI&�`����a4F���1��5�Ξnmk>|D���'Omx`P�axTw$z���+{6�Vz ���-O?����[��t&3����m���[k�6��VdBD���sͪ:{��+n������d-���x��6=����y��f�xEtuu*����?�{����/�������?�϶o�ۼy�֮���mc;����Q(hy�dH嫕���Mʈ�L^$��[XZ��o�g?�L���ד��4d�N�򑰸��!�����%؃� DLt�Y��܈x�_��׿������WҬ+�|�o�F�m��3��Զ
�I��ͼ �SPI��b���:��m��_�+�\$���E�b+������;w���B��&�sF��0C'7 D�����Y���/�;P;*v�6��u�I�ؖ�~	B�]NZ�Z��7��nuUh��w����6�S�6��N�0��0N���i�5�/_.歕x��,����n%����9;r��]�}G3�\ݑ�bL��=��O�����~c�NB�W���?/Gc���́��#)��c��m���A[^I��"���|�u+xV	�9'I���"��tsJ�* R������JTw>�E�א��GGF�{g�j݀)����������0׈�Y��TΘG���S���Y	�����:���唼�a-3{�]�o�]W��ss"���c`P�sK$jW.�Κ`�vuÞ��q� ������7����s�+e���h5W���=v�ӟZ��d�`>4��s%��х (�;Og�e���Z�6:�.���X=+C�z�'�  D~�҉�X���u߷[�k�k"Q�<pH=��O�<�Ì�b���Zb �]�%&�r`_J:�n�tZ]J2�;��LeܑhSgI`���D7��,�R)g;wm����'���[�X��
p)$���b�o���'w��A��8�E;6ۑ3?��ޭ��ʺD���|5;r���RQ����,�3J���t�3����nz����Q2�"���lk+�6�uئ�mfa��V��Ȅ�p�
�E�������;����I+4L}���YX�|y���Q�ZC @�}eqE�N�O    IDATOO��Ŵ.���=;��b�{z�oeiݦ�ް��;���rYV}����Ϭ�n[�W���kS�QC����exj�s@��o��f�C�O�.G.3A�|��\�Y`�	��#���.ك{���|��q%a�~�c*&�OL��mh�Ke�Vȣjw���.F�-��?
�&��g2i���Z���,:'H�3��3���ʥo,���Pӳ�O$����?���u{6� m����{���������o��~�k���C�$���!	rӼ8��g�TB��#Oq�xX7$��x*�g�_��~s}x�s���"����3u�g�|��j���B�K~p�V�sv����5E`H@ӕ\���%B��L�2����lr�T��j�Yo��ݕ���]^�#�r<�\���)!-+�IKgKv��I;� f6QjŔ=�yަ_ܱVE$F�7h%Yϖ=�}���v���J�G�ӰZ�����Bs�⚑F]�
x2]m�T�Ȥ�S~�/��^�d��]����1;v숄d0Rڷ#��]FXft��k׮KY�&�ޣG�5�549M��A?�`�Fm��A�j�|����-�g�֝�����Z�㷇WoZ[$��52��n>�o�K"�&b1�j��d�Q�@��WJ����r��
��M����{��uu�Y�W�t�*�\�Z�T�z{���c{���&���؟~��Y��?A�	Y�z:o�JE�/0���#��[[{��}�jܒ�i���
�ЩN��c��D�j�N����O�A��6HW,�#̋N2��ʒy�u�hkw��D�F�l}�뷚$��J�٧[�/�bc-� ~>�?���9���V���1,��T�(Xn$Sg`d�Vf�M�fV���l׎���~���V�md��j4�aʶ%���5l��-L>��wΙ����X�J�n����'?����={�t��	��Y���D��9��TJ��P'�Q�!���V�W�Nn�6|~�JUKgVe����C�F�B`@�ؙ�D�:��[���?�0L�iP�a3SS"��&���u.+a��#[}�s����H� 3��	��������=$Q�gS�v�#�Q2Bʾ��olcqڼ��!�Y81`'���Z{��~�#�f���\g���5�%�
<M7@�@=�'D��-�>g���O6��gg$����:]���0����jv���\j�.)�_��pv�{:D&�"�
G-[b}�[��C}R#����.1�X�H��E���N��lx� �g�Zq^p	r�E�|v��X���o�t�⭽J�=Cc���db��Vt��D
�KrE	iyS�_�nt��Z(�H�FRxJ�BB��*i*�uH`[G�u�={js���KGF�ivK�r����oW���K_ni��:��~�r�)i6�a��=y��6�l�ޮn�ta�c���]X�7������G����f��>o��v��I��𱌍�m�nx��=��s����/d�|{�4�i��d6�D���ֵ�VP>��4�Q� K\:m\�(J�� >�� BҸc�t�"��8yL��믿�j׮"��V���ж��/�8g���P�F�� E૊�T�f�|Q�O�����KSx�Y5e�<`Q �3f�������ʜ�w�?�+�ҿw�c�������ˌ�B��3oe�ݺ`�/�Y{��f辠�<a��m�{�Y�s��,�#�5���{�Sqe&͉��<(4:6>��b��sJ����uu�ؒ����0;#�͝������W�R�4`�.]�Z�W�����u�w��b�S��ְطۊ�m�d�U+�=��լ6���-�6�e���ڮxGs���%s	Rm�j�7�ؓ�����F���R2i/'�-����Oa_�&_>�dj�*����:��XX��C��g����	�O�������?��c:ra���!$�QJٲ%ڻ�[��b��X�*���-P#��p�$ғV�� �N�Tw��V+P#�c���
�y��٥U�Y_��Y<�&����]P�:�����s`�#�G�ɗ�qIA^R�`��"�����S'_5��x���r��d�\�b'�����U� ��\Ƽq�P�W�Tm��6�,��e�V��L6�d�c�#{�ȇ?��'�LP�0��0K�C$������U�y�ur�+�����zdA��^���2�J��5H�(q/I<0T�@�R{�E]H[%\�|n���Q�������Z[(Ңy�濎���mu����$w9��o���Y�԰�D��.�$$��d�ʆݽ~ޖg^��k����X�f;y��r[[\ˈAM�$��F�vݺ�cl���>��`G��H�߈����Qg.Z�|ra��Y'��̰�q�%�Zn�,��z*� ��$ߪ�ѕ�+b�?`2&!@Q �[�?3����E�Dk���ZZJPx��C7��6.to��S��V�[^�g�Rް7/nٛ�w�B�!�Q���&;p쬘��H�[m�)���q�������%��R�� ��#�a�Ҹ�2�!a��Jz�$�94�{_���<�U�\_���i���Z��]�՚*`r�ሊ ��4%Wj��ttuة'�s''&dR#e�|^g��8�}�ydr���sK����O>�d1e7�=����qR��_<��g��[H�@	�?ڽ�v��b]���u"+Kx�{�>�-��#�I���A��Ļ�Y""�H�EEg�Y���2R�ه�	'e|�n!tw����`��xa�بݸ~����6�o��E';Z�J-�Y:���o@fK�hT]���9{����1j�C}�Gk�ć��y���4��m���i���k:w�:�m۱ۮ\�-�VK�I�w��"�uE<��K){�ֽe�Fv�x�Ti �1B������ t�)�q� �ɵ�\�F�n_)�^�,hLW-���=JK,g���჻����-vĶ�w�����'657c���=����ֽ�W�P�V�-��zgw�-�lX��C������Gl�첁�.�9���o,�������N��7n��R�v����m���v��s[]IiO�<��e��1�T��۵U�ƢV�b����f�]�����G��ā�L����Ww�٥��b�����X+����v%t`$����e3��"���IIB!f����qӊ9���JE�R���G���*���	�$~^�x���X�����ϮA�p:�і�<~��Y_�眊?���Ҫ���D2�k����dk�D�������d��!�֨9Xt�T��v�Px�mҥ�Չ`I)�dS�o���C��W��[o����w���߷b��=�g�zu�� �^4X��p$$r!
d ��;~ 	��� ���|/U>�,�Sz��R����� �|V�$xَ/��%#V�WK�Gت2g���d%qM"�����F(R���4bH���q�.H���H0cymE;��ת��]���VL/����_֚��#v�Zk�� �|)��o�`A��o�['l~�/Ȇ.ӑrFkV'q�����D~�*0�Z�d�ؠ֊*���� �@J����r��.$�)�j���T�A��aղy��v]ٓ�3�������=��!ӿAk@R�~W�U�Y�J�^=�aӯY�^��D6U���Ͷ��YkI��h$t�An
���)�q=(����!	_�a�C���gձt�ｂ���V���)p8�2$(;���9��:�O
w�	Q��U��so�*A�����p2�⿫�ӖW����]Ϲn�{0���g(l=�ݶ����
�KF|s��Vc��d�;���[6q�%�H�%��v��#�-��o����,��;7�u�������H�*.��5T��E�ی�b���y��	�&*���޽{tAI�f�5nܸns�o-�y2"-
�<s:ی�2iI4;rD���S��B+��Ɨ�ѩ���m��sw�ص�r?L�����%9rvzF�ꃏ���ݾ�P�v4e'e����f�ݲΘ,Bx$�gx�F���. w�Cs)��rș�2+MK�B����ae{噐5��"�x���y����J���q��^�|A�0$W<G��p�� q�[I���>_���#���ׅuIv�9���ۻeNC��D��Tq<�XĖ�I��c���}dľ��լ�U�W.ڛ������r�ޠ	������]v������Ö����K߈垫U�Pżu��3����5����k�~����ա{�f��l��e�s�淕BŶlUy�fNу���͛)v%[���`��\W锜�?)�����7�U2���B�<����%*Vw��V���7�dt�<dT������� >�ZK	��K�Z�Z������Z[���f>�CW7�iV��y�TxT)GQ�#�cLz,_r���#ު2�v�_��Y�(� A�u`d�8��m�k�`g�Ae5�K�/A
�n'1���u=�����]��
���ê�3O�W�&b�|Z{̬G!`@�&�������W\��:�9a
gr9�"'$��16�N	�`��/JVH5�G���Ƞ#eF�������L�sE%,PTڬ^c��ol��ͳ���J��|d�X�.�9�sqG�".���I$�f�����k��b����dW�T�>�0���;������@ixG7;Z�jR�Y*��񸂌�-����W�p4$�P�@@��9I��T���g���p^Xs���+Ho��ع�Jڞ?�f��^��Z��*YO�f�{����{-_!<6k�8��k~�Sp�ŃQ�itU��:��a�P䋳�s��v��xV�{F��0��utu˾MP�M:�����ۛ��g���y����BN�#H��^EZc���.�d���ԩAH�2@rb�$�*���l��={p��Z��t���Z�����G�~!��f-�q�ȱ��)P*�$�g�/�?�Y|�9�}�=Vȁbl�� +XO]F#�>B:�[]%'��FH�D��<�I>wg"��Ami��d�"1�{@�r������*��.DӇrhI�g$z��A#����Q�ڰ�7�r�m�P��t���uo�g�����\ en����\>ڂr�1b�r��˚
A6}
p� I�qE(O�7���S�E6}�zJ���<`w|��W�6_8f%��~Lc@9+b�3}�m�o�q�%�	@b�]��z�Zm������!�8T�b֦ly}Eg�����)W-�����͕�v��	�����+@b��c[���/�̙��X�x� �|�ۄ�����٣{����-��Kww��_��_Tc�3�jj>��>��ݾv�������w�h��.:������܉]��l�1�!�8��O�h�و�Mx�D�̜u!:fV/�a���dy�I�]�n��a�N��b�u%��x�E�
� (3��!h���C���r]']9A��`F$p �3tJi��
$����g&��8i_UePR�@?O`��B6��=�}��՜#Xy�T��?������TF�"<��8H0t��yŢ�@�E��� YP��T���� G)(��$)�?;�l�u���
=~��62N��ș�qz��F����U⇹ˋ�P������\@#I�e�4�Ӟ/�m��Ԭ�<�� ��������%��xlӓOE�*�X{װ��:de_T^���6'��}Tm@��hUd5:r����[��C��HƑB�3y!y�gt��h���pPA�����2'e����Y;�t��)9G�tR�˖�( ꇈ�<͕�V/u�p���y��,1#a#���<�ݼ%{���--LJu/��[r-o�݃���	���-����(�5��;�N�I*��s��[��p�K�9�"W��(�,Y��QT�z��Q�`��(�^wm6�5֪��s�+5Gg�s��/�y8�޼'%�㚨���g��

I�=7���gr���o(�꾀m�a�X�R�^=�c���6��[�k�Ə~h�N���QD:!�/�<Q��J#ߜ�K����"��V�� �q�#���1��o	��u��M��dr]gÍ�ܸ���^vr#��(��rQ$I~Q��E��� zJ���<ʹ��)�U`���^�|��A� yx4$zf��
G�5���WOo���(oX?�`�r�un�k;����4́egAЍ�3W�XI��%t]����jm�T�Pp������&�Sn�V� �v:!niۭ��K�	������L�-�w��9V��<��F
��h��{�����ݽ/���{�d-�-�Wl��]�Vm��K�{�������A�3h��zZ"�=}�X����c��u����+���n����Z��{�������'��IB��k������C{������x�~����v���p���.�?����fJ�S/�;�b�uy(�1	� �y��m�i�q�����2����̤��Á  Qa�48`��[��"�ù�:�%صUcd_%T���
��y* p��hǘ9 �^���L#�*J*TX��Y�p�@�k,��E�
b���@�ɋ�΢V��}�j�C�3��~�j1g��K�t�T�T(X�R�#�'�xG�t�Y���HQ��:����<�BE���kE_�x��T.W7�g��A�n�IГ�9I�% �mSO���~��Xު�g����"I��}�og`��!�+v$�fB�1Ԗ���0���"�QP1;�j�V�lqvJ�4�3�a+[���[���2��E %H*���`���K(R'��q��V��߹Y�KD��Xm#��E����'�4���Y��/R9(�E���cp�8+�l�.���f�o����q�A����p��<��e����V8��ձ`�n�O���C�mm�˔��ۖ�����k�״�KQ@�(f�

D��y!1�2t��3�5V��%\A���k�&��g�Y��:��W�e�Aϼ_�����L��z��4BP��a��?!�t'(�u��R�g��J�K� ΦS�o�n*g�iأL�Nt8ޢ�0��d=mQ[�����[K�c��U�����c{%7����4+��J�t��"i��>��-�BԔ��;&4>*��4�W��6W`�Y��4ߗ�nHQ�d���g�jL��'$^P!^��EE�\��и������w6���
#V��#��;Uܘ��� �#��ꀘ��ޭ+����Ik����Z����v�w���vh�"0a�焆�c�=�(�t��n@����ƞ^�3�)ৡ*
A��#v�Fȹ^±�Yvk��ɜ�A`��j��h@(,�;�:��%�#�Zu1O���O;��W�8d�Y���|��u�^������D�W���!5�G�צ���}y�+��ZY��B�B���m�zqb߶?�O��oL�?;k��z�ߤj��^_H�<j����ɷ^�Y$����w�R�A9�+ѡ�Ԇ����禭R��^�y7�	��P������)�-�{�2�p���ڙ����+~@����t^5�q{�<�h^���^��А�q�aEA�#�Pw�����	�u-���%T^�o7����X���F�y�Hb�RY���Hw�k�F$Ѝ��`w$5?��ϣ@����1#&9I��q�P�c�����A���F�XP@�{�k��tSHG������L<z?���\j���|\�g��]{^���	X�&����g1� }��T�J���ԪD;���Hf����-ot�-P �1BK��\bo&G��]�rp$��%`1Éx��W���5�ytיĥ3��oZ�t$<^G��yc�պ���f�Cwݾ-2\g��>�7�F�{�ܴ���Z?.u������j��S�l}m�j��3]a���K��o`�Z�;l�n����oS_�3^Z�g!�>I�8o��\���Z���I��F!���&�еFB&p��I�|5�Nps�L�ٹ�\�.�Y��h�u]=���X�"��v����}�qY{V�[p��T3��)��ȋ���Ogk�f&�H����O(���Ͷu�n���D._���7`�H�6�i[O%�D)&@�=6-Β���.h�����{\W�&bp��M^�3�~:�ɚ�fǎ��~2刂*�"�4�׷�^�����pK�m0���L�j    IDAT�ȹBl��/���[���T� �Z�(>Ƣ^�ԭ8ﳂ�y��&ݴ�DL{V*�N�ݺ����@�]BL����"�LX��b�F�L�&W���ؑ/�>��t#ɴ�,�H��\q�U�ʕ�$�A��G$}��;E@6���c]<�OH[3vw(���q#B��Ӻ�:��@��
c�X� י�HȨ3ni��{2��_u#�PH6�Ľ��eiK�3�B�Vj�	������m��zyj��?�'����� ������.^���\�7^�y>���H�u��ݎg.����QLZ0���LLb��9����&�{dG��Tr�2�5%�J�*)O��b�6:�~��|A	�R�3�/��O��.�x7(��`j�H���uh��C�yU�ό��`����Ы��w3%w��!�Cř��,�x�"��5,c5�s�!����A���/�l2�3���u��A��^���`�6G�� q}���o��~>$��n'ש0d)�Hf��� #@ܿC�	�.��5n@V�"�����~?6����ܟ7�������8�GA� ��<h�"�k��_���-t�/�ZInX�=!ȏ@��
���u��t�}�4�l4�η�Ģ�i��Pr��n�cC�zJ�Ƒ��Ї&D�g�뫸@�H�0��uc�ʹ&�4�mw�V5��D7�;�0�VwIn���R�d�P�3�	�-�p������I�rD��	jU
���H��D�Eb,�\��ܔ@��Q(��v�`R��\S�"΍}�_�9g����`~7 }��?��3!mè�n�@�{]w	/�zM�k�&��i�m�6;��*��?c5 ^SH֧�n��QB'ȋ��;_(`ɕE+�׭V*
���[w?��V�kD���ѩN4����Rǈ�u�XĹ��@<!.Ppp�xv�s�	���L����،��+)#��3"ɿO%3:G��N��q�!��ăl�pR�;�V��+���F5'�5Vג���j〢��X�x[v���Z�����|��~3�nx���f&����Sԋ��,m�l�o��>غ�꾀$VY%���0��ڠ�����3onMP�qO�ŗ�*%�=�MQr+q��GCLw"Ly[��h<��2k��5V��$9���K�#�]G^"B��d4�Y�=�q1��8��9�ܯL6��K�AR$Q|Pp�3�b�ys�&���]���׭��Ǌ�G�E�W��
�K6��1qr���?}x�ߘ�������+�v�Z;�l�K���Xh��1C�д�F�ă���భ��d�x���ү}�z�6֗��´�-/X���Z�`�|^�_%f>���\P����\v�0j��}>�;v5�z��D�$@Dȡ�Y��{�g%~����:QK�K@bMВ��z}�V5����tz5�2CJz�������vX2�M��n\�h5O�Ba��ba) ��b�YP![T�!DA	��	k�ஓ"3�(
t������ۗm&�M���U�^K��1��1��zb7`���F������]�a
q�qm�]�[W���� F��XAQA����5�.P::�;�� K���(��$a����&��4�p������`#E�C�67:`�) i�][V�R��v�Yɼ�աm����	�4g�U������g�}�Yp�5�8����J��g��W��-��������TwO��<+�2��N�V�G�r[yur�ו�B�e�Ba9�3��\]����v+nߞ�oё�X��>Ss��|^����l�k���{4v�5����O���"v��F���zX�Q�<���&
�b�G��P��(�_6�(�%DVd��[��`�����	� D�[
K;q5�ݍ'$���;�I�˿3�it��q��9l� ����A�����p��E����������Z�+��l�>di���b�|*U����?�ow4b2Ex(&�z��p�p�Qpd�f��s��e��s�*]vc�����Yz�Z�b�hk�<M`�&ڶS�2H�O��t���Uk2����w��Ů&ٚB��^YA˫F@ES��ɖ� �.���jR<+0dO5H:K:��1��郕�x7�.6�z[�x�B�:�:�#�s�����$D^ժ��KZ��Xʬ�����`�3��*f$��$t����k�z�F{�'v������ɿ��	�g�/������w�*�R\MZ@�����
�]ɉN�c�J&-��!���#R�joiׇ�y���|v]��>8�-f6żf ��H���#���ܤZ�ܤ�ˋ��^�Ե-Ń�$K��`�}ǥ�x�G���y:y:A Di�7�f��w�y�����V-�t;�kvm.h��J� �Y8�%�H&x���i���x�]���¡>�{ȁ�8�.S���U�}������R�3;��f�v���?s�����ё��5�v?�������� �=����.��	8�����p�R�rc�|!+	LV���L�	Pt�ε��UЀ�8Y]KY[�Ӳ���é�n�4ߦ�f�h���q�[~���C����1��	jE���l�=�����u��$�f�*[��S6g�B��~��	��kp8��9!�VX�t�'��MHc��r�����X�^��0k��Uk9�l��[A��G0 ��C�,x��/�54�0�$�~��$�
_��7�f�ߎ�P{�N4��w��{$��M:
{:����P]#��y;.|G�kB�
�c���w�3�;}�E�.�����:{�>1"�sbT�X�����qs{:A����S$�s�����Q�f'ݼn��^�"�?�t3#	y43E}�f"wl���{�;�u������ �t�l�~�,�+6YdK��J�ZTi���m#3�3_�dEm�ԴU1�JK[B�7��0֡�ú4W*[(�.a�<�˓K[�i�ꌵ��8��Hºu`�r� t��"W���T֢�p�Io;��;�]�yf��#��tS1O\��		��)	�s���r��+�6�t�=�*͇D�N��1uWX`��c	��yV�nB�>״Y�j��5��z�V5+y��Db!�[zg��V˲��s.~->�m}���wl����3'��7&������7�u%�W��-���@��!=�$�/|G`���H3B}��F��ɉy�����aH��y�64�	a1��&c�V�
{j��gk¢���0M�f�XM"���5D<a�¡13o<�Tg��5�O͙$sxUau�d#�H�$4��	y��?��z���\�%!Gd����tzC��P�]����ąz�L${���s�@)�A� %b�Ԡ��<��	Zt((�Ԇtgcf�$e5+P)J5D`���<�)x��G3�@��Lpl̄yx�g��+���${���̈{*���F��!��ϗ,!�;BA�]lZ.�<to��V
%�-Y_�����{��u_�߭�{�V�����f�b�(1(P�
�my䠱Ɠ��gv������؀x�9H�9X��I���&�9T��M��ί��ofV��#�fW��;�|��%%�����]�5�����b4�!{u'��w濋1�Q;��<t��pcʽ����V�H�&y�\��Xx�k�A�n�[g�,$���s�#n@�7�i��\�D%%�=5�f�/��(��JM�"Yj��yU�q*f!�� �Rf��xD�D̢�%�(E�Bu��)]�i��4�j��G;���m,�	������x��$��O��0C5��#�Y%Uk'N�\��U��jD��G�z�a�]7�H��BA'E�d.#�D4��iHT3�s�g1VEX52l�ȉ��븜�Y�s+ͷX2���c�E��Nt?�j�U_�u���3�H~|LA�J��qc���F��a�������,&<W�@LTUv�ʔ�{��i#)�Q��H�JC�7� $Ş{tFas���� �z�Bo2�d�05-G=j5�ͥs�ڞ�N�qʎ#H�iPV�f�u�M�5e#��o���D�[���������;Bm�\#�!�C����ue��K�#���$�3�+ �h�*��F��r�+�@�8��@VT�)��0� �|/z������b��Ѡt�J���\<�=��J��o�;,���)mp�a�pc�֐�h,�Wv�[���aA��^���w�~�K��Z.��*�3�
A��a�b���⯆���X��]�	%03W��b�,��ܷ���u�|�MsRP�hv����߂.��6�"��N���l��m]��u��:�1< �hEk�;9�g�J*�ٓ�t��/�4�H���r$�ΰ��S�;�:m������cx���2*�Zjw,F��@
z���بQX��4*6!��⽽bh@'0qi�B,R��.Y��]=8��]%_YC�0���8�s�kց��.�[���*��]�?7ˤ������b�G1/[�X�s�*	ݽ^��v'1)��k!/G��+\� BP$�I	� �'N��Ɍ�JaQV;��K��<<�\�Ȋ�t7
9���H�6UЅ]߹��&�б||Yw��JB�g8�	]��yp���:�~(62�T�<6{]�?������V�p���P�i�P�PV�4��Ǎ�l>����!�Ø��.^gj�i��5����Y���C�F"�:@R(M`�,=�����A����̃C���]��Fb$�vz i^;HP����O�<D�h�<s�w�:�pJ�ۼVt\TM�,�d��琇nWsMވz?䙑)]�2������_w&��z��;���E6�����k`l��������pջF�.� 0Tqj6j���5�=��YD��q �5Q�������q�$"#v՚x��r�攩
��w�a���P��B�m�� �X�i�U��Nҙ�|N}N�$�NB�s��~^��*D�z�~q�����l��̴#1,���]���6PZ,�R(�@�5-Io<��{!S]ۮ!aF��jb2��\6/�Ar#�q���=�wz*��Ud�s�s�u�c����b�s]C䉰YU��W�k���b�T�6dU!�J2ؠ��t��+�.V�y���ђl6aE�媄�Fu5�3V|t�*x��J%�A��t�+�	��k���~��������K�%c�N5ch��´����k��n{�ߝп��ۻ}��-#����������l/ٵ+�T��@:݃5k����p���fJ�8ECJ�ڞM�����%��@N���S�o�CUԴ,T�������$�I��Hu�*�O:P=�7�tVM��"Х�C葢ہ����7��^�q�TU7H�MK|���]�+V�%L��D�#��Z�Le
��eXL���)84ka(A�C,�C$�A8���1�ڗB�e��!����;�!G�����ݦP��IFM��ӗ�z�h	E�3�K� �F��1;�^��O��*"R�;��.\χW&��'ۇ������+�N/���	^>[��E�	��Hu�b K� as8/�^�bYv�=�Abx���-l�x�8���zl��ݴ���n�麢}\p���b�H��n_�������V(��|�cR��N���j�!�\7�ߝ����3.S�"�u�A�}�3(Nc����N�:���#���X��=�I�^_���F��w��5З�U�Mn��#�+ӄ){��t�׌^]Y)E)F|o�!QUVQ�jX5w���U��-rG~��S�iK�0\+(�)�vȳ(�S��U:+awlC�,��}�?�&YU��'�;|ɐP07o���ul���5�Rг)&�]E6��hXN�Б�,�az\81qxe2c��{W>����g@��^[ `�M�5g�X�SSyg��=Ө����6���I�#���"��\oM1�iL"�-�Z9\v�I^G������F���A2��U�xBB�$�3ϑ��s��xZj��N"�O��/���Y�>m�B�ct,�@��p	�G5��h�����3Q�6d�w͈�S W�_�H���MT82��^,�<�e�����цn������y}���$��Ib�O&���U6p]<��J
�Ra��A�B�x�A�1S�0�1Nes�0#Z�U��4J���s�bA��|�8���`vnK��D��:w�l�RI|/|�H�Fz��^��;��������{����xz��jKb��D竦�������ɚ���-�"����+��UT� S~(��G5T�p9�ƣ(����ų�cIW>��&drY�g�[W�|;22B�9:;F>�\yip�z�{B�����n��4d``P��Ƞ'|�l��b�O6�L��>�'KWΉ[Z�9����By^�!�v��W�Сt�<o0˵@��M��x�V�W�K���`&�h'�p��P6��_H+��rs�I�h�˰��&e JO���~��,�<l;��l*x]�	����!��Qp	����Yζ�H�B�T��k��!��ah�*Tɠ����&CMKD%��x-�L¢�N�	�:� : �<h�V"m,(i���d�� j(�'�2+&�<�<T��$�0Z�%�J�����}�#_��DvE<��]�
�Z#�<��1B�������,�;D5e~L�����G�##"��:�4��`&�O-T����<,�H��}����P[������Ga����G+YcH���"RTx��lR���=*\T5[<�b��fmZ���F�j�T�c��㲓�Oҝ�\$��"OT��������HH�(�D��IW�H�I�J؝Ո"����D�L��]�C��+�"C�<]yj[�����ĝ6'��DNһ������7��;�`��p<"H���·��f��c"�Ь��p!�q-B����@kj��<;4) �EYD�@2����rxD� ��P�/:����p77�A���:�!�8���=��.�%�=�.Ӣ�gGK�J����ϱ-Z�t�)uث��G�Sk%���	Y��$��3خz0hy�,&ņUC��:fG"E䟉�* $�\X-��Y��u�z�2�׋3h�ș)�,��r�:>�%����G�O�;�ߞlF�dZ�Z�����2���ćÒ��߃�c�%�@I��q��rg~o��8������3m0�ۇ\(�<TEvݾ�w«P%i��<o,�T+�M��Òz�Ƃ
�l�W�@��+�%EM0>yn;��H,���I��"�m܄U˖��D+��@?
�
&�'Qj4�&�Hl���E��7?�w݆�������OO�������xj}�I�-֬���Pޜ��~eA�����۰Tv�Tl�Q���h�I�UaGFY(1~�<�jYf��0F1��*�H��s�{t8���g+��	�R�@/uq�"ە�ז-vO�bQ�EchhD�v�La�	+�&��bAW0�b�+)�2^ac��;0��b]��Tj���d�dFl�� UJ^W�C{�D��u�L^��6�7���mBb,%��M6�p����%� �%j�Je���j��}�ɭ3Mr¦��x�p�����q	ip��>�/�F�@��Yh���ʕE2�W���.]���H�T��<X������� _
G�И�VόκI^#�S}�f5���n"��C*�UM�%6��	i�*=��A�4�Zqh[�3y�~��̢иG�pN6�H�A�kI�>=9)Nff"#��,�'�+��jM���*\�!�^&�m�K�{!ex�G��{��E5a�#�b���T���A��ݔɶ�w�f,�_'�N�D��O~x���ʡ�	����7`XN�'I/"ӺG`���d��ۨW���%�-�{�f ���fF,tH����.yaPr�\5�"--��a>�ɞ&�OR���4�vU
(zZqYN�N��*�0�]���(���&���Z�|��2�ӴIr���=��vM�v�!�
Y��#�F62��d��DBM�h�.�4�%/>f�9�Q)�˵�V�D���@"�Ed#kq��~K��ڈ:�#�FT<0��H<']�K�y#��J�I�����<P.�N8)������޶�v���{˗P�����+�j3�Rh��r^BA�*�?/�Q�|�� �q�	�a)~�*����ڒ��.=��2
��¬�H3�yv�s�%�V    IDAT�R^$�Y@��"ҤCSdXϏ*�p��(n�F[	���d���'IL�	]/e��)�:� ��ߎ�VPV�V�0�kX-3��>
�5�Zr��{ϵ��ɤ���i2��EA��!��J�2O���Gʜ��0	�⩞�4�lؽvf<��(�2He�[�}�y~� �T�p]ڑ�֚�D���8k��	��XЍ�������}O�>���Ll�X�AN���3!!��(�q1�ú�n�鳓p�(,��:.B��^&�N.:!)�"\�thԤ��.�����V��#�M�~T&���L����јLq��Y���ҁ'�ÝZxB�p���
QP.d\����M%&$�,a�
ՎZQ�U'��u�pu1�Po�Ѱ�C�N?�͊kTH#Y�C��=�/�ON��F�XZ����s��6��^�@���'�ٹ�U����2�f�&PX�'�X �d*3�RJ���ґ�H���|qM���8��IT*��)�+�2ePRM&�38��i�i�0����Â��x%�3������sÓ���$��5�Qi̘A��^�(6�	]|�u�d�������d4�ũ�(�3!.|�t�Dj.W!�q%�N8m	��b@�RFii-ۖ�%O�ucA�_��
Ẅ,pfzLݻ�!�Tk1 RҸ��>��1�����h�����=N��k�Bi!�����c��2�I<:xE�r�H����qNQ2^I�Q`+�o���rSc���č�π�lRG�4�VcA%�Z	�h��~����� ����u��I�R�k��v�&Sv��Г�!��
C��f6Ł�3)��T� est�yP*i���|���gYu(k6`���m�	�T�~,"OB��l(��j !d�0�N�h��
�KC�6��mQwn5eMCu��b==0SYqd�fc"k">���Sh#��1-��G�Q��Hez��t�{��󎼕�?�Y��xXl�jMP<�u�T�n����\s.;db���>.�C@�,mF[�<�!f*г���]D��=�ۂ����E�O�:"������#����R,;��Y��y��5dؒ���/�;������bՂ]�A�,�
���ͫ'R���34��<�����';"@t�=>�Q�B�R���;&E�P�}מX��]7E�.��Z��Mr�fsM� �S�޼>$3s�)Ƞ*�a��r�9�k2J�x���wV�b��)�j ��>A�k�Ed��t$���=]Lz�=���ͣ�j �0�f�2�9s�⤘c�Sg��m<���i���G�H���NA��߷v�w�v@&�9��,y`��?=�����}�CW7��,�-G�?.���8����#�z���4��!1�f��h$�a»�@���&�.L���(��p�Љ�-��4�Jk��.H��3�z�����"��JM ��;э�<�ԉ!��Ts�C{?�ы�����BTWӻ�Z}�$�Ea7]DC,�,��:f :�^;Ws2E���Z�ޔ��RZD_����oa��Ii ����� F�oB���CB����/& �RK��D�B�^��x��l�<��rx8�;H�?t�x����2Sd���������X�������;<(�!��n�c���xZN(,�F�g��s,J3���Ӊ�gH����L���&���/�+��H8��r�ӥ9�I��ra
��!0U2;�P�U�P1�FW2G'*28��JE,-,��=�T�� A,�v/^"&���d�~��l�X�*��'��^�;����7q�����6#N�	�R�nC�oZ\�����I��<Q��43"��dy��pZ*S��ی%���`�l2"0�����l��i�A>Aa~���p�P��IY��Z�,(r�<A�TC��OC�XԊ%�BI�I�v2�dT��p2���a�&�я�I��.X�#qV$#��r��V$�z�$"�A�fz�H�Pop�F�)���YP2�Ò� �C�ø��t��x�fHP��Z��z�,�;��ɰ�"<t笲D-c�1��,q����8����*C���0��lpRW7!�uI��b���(�捹�:�e��+�� R"[$S��E��Ƅ�d2^-YY�]D��i�Mҗ��o~�w��4��QȐ�-��6Z��p�K^���@֍�p|D�%N��&��g��l��P�Pi�dl��޲)���1��i~Q��k��(���4 �;�� ���<�h d(�4����d�澜&b��P���z�ӜE��p����od')Q8+�=Q��F߇�kh5h�TցH4��ŉ�h�jI1J3B���;�(ᐐ���C�����5K�n�D�Z�j��-��]u׋H<�������ڂ�p��'"W�A<J�rI�\� j����3��C֌`e�wb����y�]�������^�p�{���Z�۲��ot�!18� ��ظy'
� M'�H4%Yǒ	N'��F�S��XNJA�ًNqfR.����	%҈�i!�����Y�w�.2�����M�u& E���xg�J� s�;v��af�� �5�k�ad��	V��D�uL=*0��n��W��b�9>��_�����_i���+�hB�z��ۯ��.��=����z�߲��[����@�B[e�dCh�)�����N�dB���'$�����@9QZdzR�B�Ң��� -���T&$}�ŢM�7Q*-I  �!#��Չ��H��2ڕI@-N��tQ�$'��e�E��BO�W9-A�)�b�&�����0o���
��}񐏋��Eq�:��(���]�Xf�]9N~�Ω��BG*�CcaaI�9����$�I���V��Z
��Cl�J�D�F>8�<)��g4�á<�������ks�[�l�i�x.��-b�z�К�g���8�ɗ�}8WJ�#��	zK��p<���:W7�[��ڸz�8Ν8ϩ�T3HFzK���E�o���P'�&�Ωdwl�h/Z-U��1�LI��/!�	�T��Ii�b3�RBWbh:���IT;,lJ�x&�8�{ڭ��e1�0���`�8�'�1"�Jf%�}H�Y��o䵓LB�ˮ,�?_�y~�����q�b��.�	Q.1L��ؔk6�	Ss�K�P�Gq~RM�tzK���$;�Xm��آ^��a�L�:�ӱP��U����T&�d:��B>֝5�J�S�8�m��(�;>7䣰���<&���ɥ���=�@�gTl�T�Z	���1uI�S������@:Y6�mى)��c�����9S�x�j��8���{D�96l1��☹t��)�R9,�]	AD4D�A���Y
|��d�P�M���lO^<��,v��W�d���"ڥ��հ!dT���Z,��b��>�Q��I� �D�$�TA�����ފ�U9��#��E� ��B����^�C:׃��^�	�%��p#qx�	|��SdC�o�����m���߅��M�Fu��	ju���UA_ѓ�}ͺx�]�л>�7��������������ڡ��V[^V��I0R�tv��e���,_�~8�K�N�R��`��	�Q��4�[XB����ྏV݆�]�D��fZ(�;���f	�A�*
��9���_�|d�'o�0�j�b>baM z�Kx3Yh=YɭU��rjN|֪М��V�,�z�cˑY[&�H�bG�²8��H$M� g(C��D����]3�+̦�iZ"f@�[��2�~�I\�t
>ٖ��k�c�}����b♒.	|*�sN��H;�V�>���]`3�L*@�;l�F<��Y���@��Q�UzzN<�8}�K�)�ǨX`FQj�� �xj��^���:C�\����"��A��y�,�|q���dP���j"aq!����A�F�:�XW�O�w�F��͏P���dB�}ަ��1�r3�^���X�J�B����	y��A]�^P"�阍t`g�a�)$�*J�`RA��JB����9�:u���}�`r�)P,w�
i������K�kb�'�_&�&LR�h����\rx�eJW�i^���^C:N�u�X� �m���=%��,�!\��={�En��mq�A
c��\�_���%�-U�K6/$�����`�M/��$y����k1��g�R�!�J­39M=C��Z\e��j%��rEY�ru�5�ٗ��庍{WZ%GذR�lFDz�3Q��ux��DV��f1ix39M�tÔf���y�t"A��C4��%$�0e�MD|K���s�1~�B�-��~ۀ�Ȣwx5
UK�sa
tS�-���*0ħ��tJ�Rl�j)�&��aA�I~�%���gҭ��u�XH�O*ֹ�VA�\"���CO�2)�j�&t�o'�P �<�N\2'j���9�h�	]'���])�Xmԥ��Ó\^���I�CLU��鹨y-��P���̹���PI����U�QsL�s��s���I�#��YpQ,W�M��w`�ɷ�K$�
�Ra�.�]#�+
���s�CAR\҈Ȅ��Bt�� �.2Xs|�檨��gS�$�҉�P%��b��]m��,�P3��i(yFoٵ�h~�Ͷ��B=��&g`�䵍�¥X���xD5�bf}H1���CE�s���X�ˎ�_��?.����s�����6m9:/���V��(�=}X�~+��_N~$5y�p2�0r�����[b{׉�4M�4[����"��M!�>���g~��e&���f�rhZ=�ts�8)��%��j ���H�q�4O�+I^6�dR~���E���OQ-�
"�z��{��̤2�'��m	���2�b��͕��a�FiQZ&M�pD��J2�3p��x��'q��	�>v���	|�hŇ�
%d2�*��<@52����&�G q�� ���ۈ�1��1�E�G(q	h��1;qY�-�G�����< <�����Vյ+�h����R����(�N����َ��i$D'_�W�t�=O����d���x�5!LϢʘ���L�-p�p���^Ź:<����ă��ܯ��ū�� ���G�f�^T��q)�b����	����bP��q�E��?�I�/ҥP,X}��9�z��e!Q��-T\N�t���٫IAW6a��C���Ԯ�JC,\J������	贚�@��|�=4sBbԓ��}�0�����"|F��5�I�0 R'ɍ�@F"'S�G���˸�,e��r�0N|a� �����}��ܺE6�-q3FQ�(P��� ����0�U��x�+G:�2��6��`W�#��%�6�G�7@�qL1�}D:&%�F5�@��|��x��I%_�qzZ����� u:�)م&���Z.�Diٛ�b�z&��H�g��" w��e?#	`j6��,N���������=CX{�TZ,���B��QI� B�.r���bA��v����*�DB�7T{�5@h=�M-!]kG��6���qRl{h�+h�kR��j%�N��rʔ';�P�CK8�SIB��ΓZz���ێ��8�
���Ң2K���Dp^ �$N�r�;��=�8�m'�}[Чt&��J��nA;:�����s��%����TH!7���R�*�!��~!��jɮT��OqE��2�#'��B2�Q+@$D�H\oQ*k7Ь�ѨV����hv��jB\0>!gC�K$��G'�;�$dg�Њ�J�~�iar�rڳ��ױa�^�\�z�D��`$yD�����ȫF؃e/��ŏ�$WA�i�B���(������������<����?׽���@�V�	g�Q���)[S�ע�M���'��G$���7���CO&!���S�ҡ�
%ٝTʦr��Fa�a �D�S�������}o=���������3��9�$h8.�����"�jIB槯�q-��#?2��ec�Z.B:%��r�N��^�9�F	Ն���܁=w�/��E��d�jqiW��cf�:��f��780���0<��� l����NʋKbQ�n"������Ƶ'���[.r�c��߂���юS%���G2_rʐ�{"�F&==j
��[m�B��!Kԃ�5q��)�ë¨G*����X�	�Z7���t`�`F]�iBg|�����PX�<�I�}�.�)��g���~J��LX�����]����ʞ���@�rE�@8=����]Sq��uu���p�J�]��m���O�������q��G�f�>,T�Bd breÒeKQ'��*&�=�p
X�Z�HixjU	!Ag�{Ҙ�~�����Ԅ�ǭܼw~�a���Z��B��q��$|BN~b�Av/�*�:<�0e'��U�ϰ9LD|<��`i�<�j 7��}����Ulc��${�+g���RTNd�82�Q)FA8&����k�h�[�P6�˧���ן�Z�A!�F�
��s!��n �[2�ǘf�kT�)-o�
֌ť9b���IX"�(��Q-a��9��%T�����hrEK	GB&*"H�k�e#Ew6�Ӑ��A;M���d�-ty?qn��i�\�m�!{�6����ԥ�U|��u�"m�,B|�H���`JP��PÂnh�x��~�MD�&��ʵ�@�����YX���� ���r��I�;�MS�HFc�1>Ӳ:,m*9�J�[��w�����ȝ���p�D1#���j({g����?�v�+Ji9�/U����	�E�׼�MO5M�yW
�:H�N:�*���J\��qГu)��r�*��r��D�*�ڳ�g �>�T�14�/z��;�s�gaK+������{�,�¤A.��'$	e������Z�x��6�~Kޑt�ɟ�p/~���ٺ�@���[!: � ^��Hz�s󈧔�:��Qb�.\�az��xJ������$9�Uh>l`H�l�*��Od�^���!!ǆc	�D�a�{�rF%�[q`Dl��md�QY#�J7j���~5]�0Iq�	}EOn|����ڽ��}R�?����=65�7|sB�䁰:"�P�̋�I�l��\/�l�_c�Y���za�j��~x�8�^��ĥK@ˁ�J�΀Z�5�c�ƛ�B`&P#S�/���٣x�_
�ji!|����[P*Y0)	�CR�Ϝ:�+��b��i�"��ĒȤQwZX�e�oہ�뷢Ѡ�����r���ړ�i���m�����`faI�,,J�]�����? ���'�&dFa�I4+@:?���U�}�n�=X,�^�H1�Z5|�W�z�pX�S�|�[�e-_�CC��&x�sї���4��g�07��ɫ��e{r�вeHe��c�j��#�M���?�w�z�f�������%l�R��C���a�(�]���U��:��&�����Q��i��!���v����@π�~��Xf��n����{Q������n�\��"N�8�f��YUf<�C��@��r��\���8�|�dE��^~���_QZ�@.c
pρ�qӮ�1]� .D��F�ͦ�	�Di�naffNr-h��������b���h�+H1 ai/?�+��y�g`ۃ_���{Q��>��ˈ�����R�[f��IOB����ylؼ�D
e�þ��v��^���0{�#hN�A<�7������h5,	l�������5Tˋ�_cǮ��X��flڶS�*��9�0ȣiU�a��q{��)C���"�1q�'����0W�&-F4�Q-� ��ieZ�q�i��d1��aza	n8�L������u���מEP��������JdQ�.���Mv�������j�9O,���-B����%lmj��{�iL���}_�3�i� 'K�Ʌ�I�2���LO�����F�ݑR��h�y���ebHG����`��	
��`�������x��.q���S���}��E��\���:H�F�ʔ�XU��&I�3Q���ȇ]E�("����g��B1��
HВ6�d�5���N3��a�hۂaROϵI^$�9���,�->S&*�:am����@�K�E5�]��\���:�)�[��Գ����B��@�f��Ͳ�j7���q    IDAT�~���bfM�����q���BÏ�� �mj�e��PD��|ޘ�h�=iZ*�U���s�L�XJ�s� Z�F�D��`;>J-0�p��4i�E�;M��`�vq"v"�,�j:���ų�
�xE[g�E�)���f9��6��!Y���*��9�c�r,A�(����(j�-�,Д � 6J�#^4�g��1q�����d�}YAP9�r<�Lx$bGCrOW�f��[��;�/��6˽�n���_�'�g���F�At�d�N� �������L#��Ŧ�����aل��������(�������W`իش�&�[.�޵�+8v�CF/��{������M!����p�^��/e���8}�/�^%,_���J	G��+?Bcq���l"*�'M�K�*"�8ʶ�����������P��Ѝ$�aO|�P/-��ֱi�n)�զzA�Fo��,����U��P��ɺe�y(�ģ>[(�ll�m/����0Ri!�tebA��?�0��H�����h� 1@ο([mģa8��� )����Ʃ�6;)�0B�j���K���1�f�lލ�Qu���<o>�$LCGvhv�y/R�A�SiT
:qu�:���fν�c���ˇ1!��X�O�@��݋��Ѥ!L���Za��oP�����{�ǎ�b�{�g��^��Co`b��	ia�ƅ�g�8�=��>lٱ{���%�(=��l<�Ŀ�:{�tT�v��0��sUBk)I�24I4�5}�&q�������ѴB�rL��Zd�WBK�E�m8b�w��ӿ�W��y�[v?���e/ꔦ�d�����ƹ��Q������)d�-�H˂��a���ؽ�.y�\��9聇ן�殜A�^B��2���GN���HM�!���˘;{a3������p���7[�p�*f����>��q/��5'�#������8��k��Uh�+�U��}�{��o�l�j�<�&�Z-�Z��Ν<��kcr�"�''��f����5lRb),[�I��Y��"ߋ�k����UY�ŊMqϧ?K3P�i6�F��4;����(�q��Ey��}ɠ������rtuY��m�f��۟c��IQh�,>��_���IsJ�LT�Dɕ���g����iAN��
�Fz�78�M;v��P
��Q��l�Y�� �8��k�|�]^M��L�ӳ�x�K�F(=�F���:�W<a�W+%$�m�/���%���_zF"��W\�I�\>y��x!C���o#�D;0E6K����hs�	�&��0�x��M����4*rF�WQ�٨@������Z�Ajd7�܃L���ΜRY��Պ�͢�&�>a�\�B7��&B�mDd�K	��n ۶��/~���8�1����m8�зa#G`Ѹ�<)�V<����!D�D~̂)���@�!�F<�DiiW�`q��s�ɚ�0�b-�D
���h�S���1a��+�\��)]6 ��@�"��o"��xKp��tn��b�%��v4.�%�� =.�	#�@�����$zC�����1�
!hհf0�������Il�e+�lۄP4�#�N���uԚ�d��\�=��f���[���QA�������n��[�A�cA�]����4"�z<�F�z��<]dTt�I�\;�������z�ظavܼ�V�ęS'���1[��FR����	w���@�~����8�{����R�����%R=����je�;}�|�DT
"w��hR�n�q����l���E8��-{�­��G*ʨ^��wQ����Eq��}x��_���$���6.�� ����C9T��"�b���dzݰv�4\�^@jl9�|�a����T� �@��[��
g���(Ǥ������F5�C�
D����7����;8��K�F#Ț:�f�$�"���ΥI�իSX�i������n1Ԫb����K��]"=x��#$ B��v�MO��O>	T�ѳ<�8��xF4��DBH�7��J���r�f,۸f.)+n�����=XB!�t������`�XEoO3�q��!̜9���^�u#�ٵ��Y���8wy��2\�^�>l��Al��V!�5=Ob	I�5O��_PgAϐic�]a��{0_�"I���*Ƞ��g��{���8�\������LNa��ی��~
=���j8�}nsZ~V�^��{zk�ߎrKq�QG ��G������$Ϥ)�%�O��X��#c�2�h�!�Z�[n݉�9J8�ï?��'�C$ ���3�w������x���Q���p_V�V���kW������bG��x~�$��-w>���E��A����¥��@�+�������G���JA���ud��z�0}�
N>��+�q���
�,��Ξ�����<"�l�w7FW!bf�x�M,L\���<!�v���m��GE�	�Q��jbi�2&/}���N�]X��`s��"�ZD�@*�u7����[12�����D���G��t�o!�7��|��Di�b@s-8�Y�?q��{Gɱ��PTAN4n��H���|�뷣h9p<���z+�7p��;���+Hj�VS�E��+��W�
-#�F<��7�I����J�"f�0?7#;n�蚗��E���?,��*�X
A؄c�q���8���6n��W�榝hYʁQ������"��J�U�@���#������[V�5�4��O_�S?��Z�������~n����T���Qd���49���l.// ��Dff�)��T�۲��Z6rA/��(M_@��ZX��V��ɿ�R�3���.-$�FSp�U������ȹ����0uA����jsObu\������ן�����}���{@<? ��,���U��j"�)�<�p(��ª����M3�\�M�~���^8��t���E��*�
� ����96׿�$lJ�%�'$Ѹ���2A2@���1��E��x��1:ЃG>�)|x�8B���+���pibR
�	#bh��2�ό߾n�w�v`��m�����_:1;���KAr'k�$��`���N<�������t3<�}�gN��]�у����oɔ02����x����?�E�V���q����,ar��X�7��'�`*ƹSG����DN����K��G�s��	��֫�+E�Rqe!�9�m��_�N˖	mrj��N#ˢPo!��c��� �ӏ���?�P��E�H�{p�C��@���>�{o���SA>�#��ޑ�Z;w���+� Oa劍��Ñ�.��a9!�����Ь6`z�p���)�K��|�k��cB��e�v���q}�M��	I]A���$�v�ۑ��a�X�;����Ea����/|a=��S�����W���0���_��� �^����W���)d{Sȥ]l߸C�4.��(�X�m��P�փ�EK���	ܼo'�VYv�/��'�Pky������q}n�L�=�;�|t������W>� V��1���W_Ǚ+W1]wQm'�N�bq���{�c�w�E��"�:0/��G2�g�1ay��!���.L�I${ۅ4a͞�kO��9�3�Г�Sn$v�-d�)�p-K�&�k���G�͡�Zp�x����X�"p;�2V�r|#���X���c�p䍗�%�F�8�vY�+(�!�F���՛�ۀ�O]"ۧ>�e\��G_>���{W��3�@8����%�L2q/��IL]:�Cy��2�Jw�M�:۷o���<.^G�n�Rn���pa���<��7oG�VA&ŵ��p��K�Zeh!�T�����美�[�c�L/��e�\�po���� ���o���ۓ�h�7�|���M$z�Q$���-�߃�{�B�RG����i����"���l�� n��AX��:j�����`'a8j�͘�Z�%����)O�08<�O>���^4B�L�o>�\?wR����(���O�D��lTù�@cv��ۉGc��5A����|�@�ր��E=0����G�������f3|�}�z�E��l4j�QaA�O��p��t1_�t��l����e:tH���<��I��8BX�n��%��W"��¦M����Ի���~�T�-��{����i'<WG�P�P>�ReW�_���g�4qIHWh�ҋ6z��Mؼs?2��(׹���N� J�8��s(�M�q�=�b����i�U�|� ��®W11~��)c!����`����r��|3V�� V*fZB,��C�z6����Q�:����v�b���ɿ��N�EdϪ��)J7�h��¥�h�r��d$F�ЛMc��e����AͲ�lh K�Wp��gp���<��ȍ���<�T�� �,~Cm���h�fa�q ��g=��l��9q���$��ĵ�'��o�P�v����-�߱�#dT�k!��U��#�A%9���5"�DY��������!ľ5)L�=!h�C܃�?�$&�_���UԚ�8��*�\�Do�}kV������ek��v�~��_>>7����{��%���*T@�)$
Sɗ-_
�ƭ;v�O/��&Ν�񃯠8=������{RH%����;�c�v�z��u�^�[!����8uv�����ݻ��gp��a|�E��9�x��?G��0�'���p��1���p�����a�a;F�!ƥs1�/K��I�>F�n����	�]8�w��
��hil޹w��)k��]|t��غ�v�$���U,_9&�~�AK֪�ؔ���b�D��e�X�}�ф���s��'p��aģ�����<��o��'�I(��bi��{�g�=�o݌���5�B�!�vx�FW,G�Y[@��/a����n�v�L=�C/�V�ȉ��x��� 9��w^}O�8��a�ͫ�K�Hxf'�Ĩg庍�+�p��U�c9�zB��("ɨH���_����H�ӏ}}k�c�\��#Gq���O0aap �O}�N�z�&.��AX�l�ǩ+�X��Qo��&v�u72#�����U��KO�%)�x���!�ۮ
z8C�k��p�����4�ؼJ��+��e�� C�����b��5Ĳ�x��y�[aD����/~m�G}�2�����kh�|l��Q��y7fJM�R	h�I<��"�4&1k��E6Ff��͛q��Y	��Y	/>���
��~��ѕҨ������3�}x��Fv`�=�U��\����C�<��#}�el]��n� ��B�6n���4-"�/>�
R}�(�!������9j.MB���N��p�a�� ���>�����|����p6���I���/`j��������Oc�M�~��1�����
��E�Z\���ßÆ��96�r	/>���?���SX�}�������OѮNa8B*�aê1$�8~��K���E�O`�0�R��ͷb�������<���BDo#�7�_�+h�z�	<��c��^|��=(L^@�����Ә��;!055#�����pu��%���^<�w�7����ȳ�5p�����Ы�G)��J����z�?�N#��������9�#o�3�b$�F�a*ղ���-,�P)5q��b�]�@��	�����{���
o�"��>��ȗpӶ��䦓�V����N]��8=�\�T�4TLsl���5�u�ܼ�v�L"Bݲӄ3?�����%�}ش��?� ��&{�\>��k��;1{邘/������#��4x!"�;��?�y$s}R��pT�8��
��g�=&�!�`�ŪM�a߁o�dE���#��K��a�L���R?���5��$�*�Gh��}`ho���C#�D�fa�?����W���?�)(����[�wp�&&����7�Fia
Vq��{��yQ,�j�iy�ãشs��CH&�X*W�j>҉�]�s?�!�e�Q-���c�ν(p��6��F�䮺�ٙ똟f�}A�.l�7n܈D6��ec���wV����N��HX�l���)Ͼ�;Tk5|����R�{�hL����<��طn�w�~���vA?5�N|��?�ʩ���j�C7
:�\�U|t��[.�Fưn��p\�s$cI��ʫ8���h�
�y�j��%l۶��-ǩ���Z6�'^���~���A�G1����ks03Yl�}+.\8��}Zv�Q#�/��H�3�~����Sb��1��q�.�G:���r�̰�Z�&�ʖ[v�Թ+(�m\/��y�m�����15~~8����?��kW��+/bif_�Ӹ}�f)P�s����/����"RLQ�[ĚU۰��=�ٳ/a�P��[w"K"��������0��	�ڈG��-8�����,�x�^}����C��Y\�pa~NqD���zxl�8`]�x��۸���b�@��%�����I�[�"u��
x�?D6�f>��oY�d��6m���zP�ԐL�`��J/_�����q�S	D�3��)��E����7���<���Ϡ�u��'��{��Л���,®�ɯ�la��;�����ӟ?�sWgq��l�s��������8=���27�t:�j��wq�Nȝ�&�f���O��
nZ�Ǫ�<�/[��?8���A�oߺS�p��q�-��b�/Oc|���_|��#h,���'~��UA��`ӽ�ź�wc�fc��>�L]<���F��/�-cC����,J��%����K�tjh=�����w�b������^{��8w�=!�����'���H���۟�P�3�eM��~��.�<q�����������׿�G���W_����W�a��ز�6AeN�����E����y�ܡ�q�a��{/��@��F����?Aua�ɘ�߷���P�X��<�%�&�L���Yy�̗�e���=*�d�m/>�4�|�|��Al�}��	;���A��jXџ�M�"l$��^(�05W�#�B�$����"n�ħ�a����p��ui�c}˰�O�ff�?:�Ӈ^��������K��JB�{��w��)T��A��ʫ8r�$�d�_��+8�+M�|�g"3�Hx�=G�ފ�D��*��wO��ݍ����ىؙ����MwW�J*y��(zR��H�@z���{w/�p����}��<Kn&f����-�E3�`D߾$�����gZk��D��2k#�">��#���fx��}n98����.�������>&���,ɽ��Mn��l���&w��A_��ӣ���)�.U���~�5s3�XR�df�QF}�y�i�"Ic`yi��/k-��**�7Ҳy���������?"�u��ݱ����Z�f5c��Ǡ��w�y��р��`Q$D#�!�˂� �
�� �[m[w��[��""B�+�B̧�����>t�AU����=��6�F��QID�ܾz���7(�K��<'��� ^��ӭ�N��ݽƒI^u#um{dR�-��5�:�-]���BOzv.o��B�͡3���@o7���'��mz\���%���i����jJ뚨�]#WrQG�$pLq����WHO�e��Ô�]�\8({��O12����8��j�*	z=���`_\�+5���_�JNQ91�X��xc��ܤV����<���o�HzN&�M�\�y���=�#�9�7U��]�������_��<;�?y�k��C���]�	�ž������ �d`+�rd���M}�Z�QQ�1Ƹr�,�c�X�	�R�dg$K%�Z�"�J��D�&��fB�cY�*�����Q�td���5�L�q��Y	nI�(��Wߑ��ٙ!:;�SU�OU^VK
���DWB�߉�|d��ȕA�/z߰���6ZpE\{�ɞ�/�$��K��2Ѵa[v�����7��e�q��V*3(�ˤ��!��L	�	=d���\�*y��Z���YUCEC3� �$�q�+F�< Y���^X��#/��0)hu&�a�Ξ �����W�`5h��czrT�9�:��ދ_xL	�/^���}r6�o��z�6��U���y�_=#o*k>���"��;��<�5u�R,Ilڴ���IV����	�7���R���u+�@���Jl2��w�����MjA/����nݹŽ��)�I%)�dҐ���-���    IDAT?�ƠL���BB z4:�$�jH5��%��݋��m�RҲ�C��ō�o�Ś���rӸi?���Z$�T�q������d�<���	ov�N���������~���/ŜY����'�6B�tv��KԽ�Փߠv�p��]�)kق/�C�p�ˏ)˴��FX][D�EK<$��~���6���&��"�^��䌍Ew��������񭋴߸�V&ɚžw�
�����c�Ϟ�f��2x�I~A.z�!l�&rG74�Ϯ��)/.������d�$�Kf���eҾ��m�o_��}�� ⏲F�;q� �\�`�c;/�0�x�ki����wc�Zj35�l�	�/�pB���gٹ� EUո�v��>���!�Q���݇^frv����Q��#0���uul\��`� 3KN
�J��|f,S�Yt9�^������9<��_�T|��s<��*�!+�/��5��|�&�H���{/��ӧOJ�G\����N4�"{���K𠫏��E�8�������������޺�E��1���7KT�F@t��Z����$:�O�I����N��u-�%�t>��ɘDII�<�g]|��9�*�^~�̂J�Ifݾ��@��cHֳ��7)(Y�����]���PY���'/W|~\$k���u:�xX�;(�oe�ex�C�V��*1��������)������1���h1
3X�D_��� �O��W)HNA_'=��LV9�tG�~�C�lޱO&�E@R��"�����T]��rE���k���n�� Y)PSZ�w�������2՚L����b��i5��)��B�Q6<�*y��҆��z�s�}�7Qj�dd����o�2&�lGoo/��fϖ6��;x�q���A���*)%]RI��0�R�f3�7�0	�x���'���y����Q�f5�xH�܃�ܺp
�"��>Ϯ����[o�4;�͛7�p�
*���'�MԷl��rZC���*�N+:�~�{Q����5�$W��v269I{�"�5�8��E�}CU�_�d�<��礸������䭧6���NU��[�x���4��R\�$ _P��aRӳhln!�>��\=^��Ł�����������IOS(cd�Zd�R��6�$+9EU���tU}�ܹu��I~q����W/ۦ|r��M��m\G�5�ѩ��G��N�?p!�HO6���t���/�a�aQ��2e���g1?;GT�g�]��w����\;�=�T#��4TQS���P�$Ref��t���J%��ڵ�l�S*O��R�l\�G������<��Š���R\��s/��(�z��9~<}��w��뛩*ͧ���[7����-��IҢ��q�=�E�&�}r.�]�B��Ζ�-<�w��7����Z�O���~�ۯ1��I��HOK������~�-f�G�q��g1ݨ.)'����y��ާz]I3���Y�[@c�����^XS��z*R��d[��7�0��.	Gb���K�YP-�*�bzҴ��os��[�%=7O&S�����xH�&��pҴa7��]I�HӉ�v:.��"�H]Y.;���y:8�%�*;���%B����PY�ȓ�)�]��/��O�#�Y��w_������=��\�M&����q���$��2ر���RL&Х�3Ye�d��)��GF5�\�)�tv�s�����R^}�%yC�sI�F�����,��8�-ř&�<�KR�\������rհ(����3��/���<�����XK*ɯ�&35����t߽�J؁F#�;q"�-��P�v;N����N~�	q���:Y�)����Z�b�J|�}
:����e�bIɠ��{N�Ͳ�M�W�����͋gy�id��y�gƝ������\Rq��Kx��!�Kv,9�r
�e1a_rW
k,���GW�L/�ܛ?'//���?���.�X@��7{�%���~D�&º�T���Bu308(s��9QXZ�cҩIOK�����O�?���a�ٮ�_X$3-�ގ�<�q�,óM\�G�V���KL��W��:��i?��
�h�(�鴓��)�۶�iKs�>æ�t��`�F�X�6gr����p��5ܼ�j�%�]��޿!-����1n^�HZ���k�Q*C$$�>'#5G�IQ
����q���� Sv7�k[)��#l���7_�]^$MP�n={_x��?ʍ�g��V���:�� S�C� ���lR,V�;:e����A���iL,/{�{�5�|s���Eɪ\���	��Ԛ8�Z�j#��OP�����McYk��eF�������WV^��
	���,��$�\��	�Kf�r�hl�Liy�:%w����u�o�Up�����k��������u��_����lB�e���ʔ��s?^b�攻t!?Yv�1g����Q�K��4L=}��O?� 0�dv��6YUD�	���8�-�X@�4�J�/~�K�mh��3g�q��-���8#�%#�n5[�&;���TI:;��F�p�#lS�`M7��`��
���)�C�m�]E��Ѷ�ҿ|wϦs�@u$,�Ǉ���8���Lщ7�HTF�EUK-(:"���]�D^��5=��խ��.�'j#��^e��	ue�ڻU���G��ɲ��j����������Ie�f��K}
qSWۻ�߸�ѩ	n\<#o U5u�����`�����y���HyE	9y�tvv�p�inl���U\��@������oIy�����������X���ջ�����\�~��䎤������K���n�rs��V�� W�1N�XH�䜃���Lb)���z�rѬ��v�3>�4 Bvq=�^�Ψ���<9Ѹz�{8��,�����yRRS��͒�s��W{=df�J>����6l%�4��~�EPkd��tܽJ��sr��[��˯�����ˏ�Ʒ@KC9��8����f1'���Go�H���T+bJ��.IPJ�+����������7�O��o%a.��W�~���JN�<��`7�5%�5W26҇V�D��L�Y�R0�#>9ʷd�16>#����k�x��k�C�޶���|�}�.Ω/~��6Fr�
����[к�0s�ii�ܻƓ;Wi�)���P�TD &//G��2�se\#z�J5��=���ޢ�����E�M�m�r�Z����� ~_�u��Ӱaa��مY��������O3��W�03����A�j�����L�^%ȥ<������q��#<|JjV�����}��+gI;1��}o�
�?H�tq?�~��wY$3ҭRO)��.D)�dlL����W�b\��?�2=��[�cQh�����A#8�^����¬޲����FR4f�^<I�>�΍Ͳs���1�����z���ܜ�7Dc�:�����5f.���_J�_�A��H����������[̎�� ��-&ų�nVa)N��N�2�F'nξ8�`���tY��9ݜ�v���մ�n���y������`b��?���+��RSĎ�2�l[�>�����^������S(��"��d[`nq���z�>y�)���zv:���E����4��WIW���D�b�*e���%nȐ;�$\:�G��a�W瑚�aζ _��yK��4
!r�-#C#c����(��?6�|�Mm[�s�"�O��p������^y��Y�&?EICu!i))f�b��pbRf"@B�RU�q���9�x�.aU�*B�6�~�5A��@,N�V^z�]:{���e��q��/�ejr���Ȱ�I*�k�N��"!,�5O�?>%ء�!7�e�^\
��fh\���'��*�W��Ѳ�5\A��V�Y� 87����4��?^`rjV��Z��%R��23��2Q����y�iھ���k�����<}�@��b����*���N:�^Ǽd���ҝ�����q`JJb���dr��M�;�%tivΎ��f�Fj�o�� ���۲ae�1���Gߢ��I�<E�{��M��Ҩ�,��W�135�����%���/㏁'�S��Ũ\����V��
	F�:�1	:�]Cq��	˳��@4.��"X)R�± ������4�ZW�?۽�B ��g#�nW��_>���.F�k�/d��52mD,a%��D왭L�b�0���]F��&�7!Qݸ}�2��)�uj�{�e2,��"բ��x�|���cHJ�G'h^��Iw�Αi�7n����g�'�wQZ^��W_!ɒ���8����T3UuE���1蓘��� ?���t�%4�z�Ƅ�iڰ��Z����og�i7���#Ks���n�ͦ�����ύ$�Ӻ�����TW���}	��()������Q���?~�KFN��͝�Ӊ2� ��,C��s��'L<F����G�*n��kﳒ�.iSa�<�?�G�S�4V�Ѳ����֨HI�`�$������)Ib�D�H�����<h�n��[Z�y̙��Qv��m{�}�It�������;G]i.�9�����1$i1[�"1B@��)���� �5M`H�k��r8���۰/��~������4��Ȯ�/��'_0;��K�w��zN�������cIR2?;,�WƤ�$�<<Ӵ~#7�'y4:O���T6���e�S_�#~�,f��^�l���-�w'�$[�u���n֬���<���b�^�Q�s+**$��`N�oٶe;A_���z�|���9/�زs/����Cԡn����{iܸ�1���1	�Y�����4�:v��w[$ow�4(j|A�Kn�{�/����ڭ�L���U���ܺq���.aV]@2���%S
g����t���Q�>��� ��O�ɐ0 
4������+k�wr��SZ=;v��M03:��߃J����:c��(h�Eh%	�ZǽK�	���۟����`ttXNl�IB�SH��.�K�p���Bfm�?q�eo����#$���X�F�Z��~5G^{���a2�z�J�	L=aqj@�C3�J!����)j��1�fvlQf^�Ks��(���������u�m����g��j'���W�ޣ������=����(���uD�QT$�f�q10����,!J��L��ʌ�'�b�_B۶�x�LOn^����Q�|��h�PZ
����I�,&��`P�p��W��Q_���S�ٰi�K2023�D|n��q:�ٴy+ɩ��y���R���#TԷp��K\;w��7.KI�H����_�K�r��y� %��+Y"������l�}�nu��2e��N��G]dV7r��QV�.N~�)�S>g�[6q�ţ<�igb��K3ȳ&�r�$$LE�T�e��F`���$�M���f��"#���-;ɮi��tc��9����N?�ӐPLG��m��zD��u�(�#}(�6*s,d�'�q��m�`2�O� �d����IɤXt�����P���ƶVɎ�y�K���2̼幗� ��3�s������ܿ~E��V�Q�'�YY���-�F:�>x�̂����ֶ��c����=�DCr
[�%'O�r��7���tx7���������K�oD}��i�:n=���0esJZfy�l���4�@���j4Q:�o�8��!���/I ��(p����b�j�3?ϒ4�ZS�o~�o����a.i����^�;�����?������$kb���5Q_ш]��E$�_��
��"jW5ʃ�d4b_X����,̣��y��(�����+2�R�J&(�NQ�O!��{X�~�xQ����;7�{�<����y������@� g��J�7��Y]Ozj���	�`uy���ɷ�Χ=d�S��ߊ��ʌ;��U�;�}�������<ȺM;�-:�v��3�l]�H�EGUy�#�赂٬'+%�J<����$�2hn݆����>��7XQ�Qi%���O�H�Z��]����~�yK:l�8{B�{V�QQ�+�C�}2p�b�J��� ��e���iIGo�忟��֚���[����� )V;�º;p�]ܺr����lY�H��5�&s��C����`�5/;��s�BYa%uS6׺���杻�����W��ߋ�og��/Q���G폸w�"m�k8��fƆ��?-�Hn�	����T�N������NNiC~T�s�M�F!�L���������,D��wҲ��LǛ��<�zA��74�b]c9W���q�c��U��MM�����̼��-/.=Cuj�����g�]���Jp��%�J0�۶�y�f4f���O~����$����t߻)o&Ii98}�CoMB&��*�A�j����	]�#�WӶa׮�f���D��R��޷��5��kW䨽(�̫G�Q^��ן~$w��? �ڢ>$�]=O�ij^#Ii�:{h�"��������L�s��		$�rϷQ���k��� �У^Q�~�<)1;�64K����$��6$���㔕����-�e������%����'g��#��$�͇�LA4�����_&
����tm������^��Sk���P���A�e�g%��ә[^�L�Gc�-y�?p�������Va�9}��8�!Ν������13�}���5r"�0�cJ�̟�<�``h���r���m��Q��B�ƭ#�`&O�^���eL1��Ȅ�/ސ��w�
�Q��-8f�xr�,�Z�-Ie��1����rt¤#��������ts���X�
�T��r�Q�eu:t��np��w�e���;�Aa0q��MB��W��黯>�jb�Q�t�-�QE���>��5Zs�����"�ݕ�������%�uv�e�^��ƻ4žu�lX]˕K�eCB�$Ӭ�$��13� W,�P���ZF��?�GmL�e�.�kq��_"��/~�w�[�o�k����[x�3����4���/�z���	{�)�$3?Q_�ɩ9�IIK���38���<)E%lص���.|���;$Ȫ�~-������ܩ4U��}M����O��a%	axc�+T�q���K�9u�2��<���Ϧ�Ǩm�c~�1_|���A�:#���GUM��F�S�m�g���`򋞹`�����dUC3�./O����dlz�?���m�ʚ[�E�](�#t?�C�c��[���A��piQ�t�<�$�Ք���{�]����Ǔ�����X�D��J��q���P�	X��+�ψ>b+��"`�zm_P��b��܋��tK�@uI����X����h�GOw'�D���,��~�~���y'�e����q�K_.G�����ٿA������Ξ�$��,��9�W�J�rO�V�3[�i�cht���"*���dS�j�D�?�;�G	��X�e/m��K}���<i�OEa6р����27=��>Os}-^�Sr��-��&S:���T�nc��c`\�`D�O��O}��@'uw("�ï�����̬\��d-G��j��)�I�)ș�qj�*��ɑ�b� E�<>Y�ٿw/a��a�M�������x�ִm��r��q|�1~����ڝ�	�>}B�n
��Y^v;5��l
r�X�w���@�z�Siٰ���Ǚ�?��^"���=��{�����_QY��/�63����m��e��[�`�kuFTIh�2�
opTI��<=����Oqx�$'k�ࣿ�t
=J�����l�������������S��B}E��Erok2���̐#+��+�e��#�"+`_\���OW�{�(i�_~�������hٶ�������~�?��*DE���kWu,�Q��7�֜�Ơ��sc2���U�+y��G��(m;�����������U2-I,�ü��GfA�/_dij���t�2-���Aݿ���YY,,.I`�ťff�u�^�?u���y����(((@��˗OA\��:�W] ��{����0���7���g��3S���"��t+)&�\�%,�`hx�E����J��(C�S8�!�����i���3
��T�Zǎ�^fz~�ʒ<67W����)��2r�p�R���lN<�I��#%#���]Ե�`����=}�;�/c�0F����5q��s�}Ky~*;�V�0�Kv����B�]��=5=��j��w�r��X� YWt�dt�U��Y�as�v23R�uQ�)J?ѐ�e*K>G���DU���4>��Kgh��a��&|�9�?�u]~�0����@��z��PVUC릝��|��9:��)�Y͡Çyt���    IDAT�7.���s�Fǋ���PB��+i�)e�*��#7��NM�&#��}r�	�H�(�oh�΁q��f�����+|��	��C+�o���M[�w�1��67ɬ���.�*ʤ���pRVR,w�?^��%5����y�;J�ج��<�<��|���:%�D}⑴*bzj�mg����W�����,��׿|�ɡnzK���w�S�I�X�/��;ĪCIN^��78A��4+:ۏ����s�|���{RPSR^�����$������J�&JO�MҬ�X�z�5Ue|~�-V�i���Ѻ}���˒+F۞#���ej��|��2��lͤe�K�U6���!�M�$+�-�|��x15�*s*��f|j���y>�IPV�Ď��I�J/��Qz:�r�I
��Ԉ���@H��j���7� ��ān1���*��_��q�O���r>����u.�Y`EiT	ǅ�����{�@C\�U(��!� %������!xXZ��ε+2<P[V(���ZV��;��%��&��Y�7�dz�Òp� @濧f�UX$�Oo\������LD�Z��&9���۝t�ߧ��m�5d�)�˓�H���l"�R]]-�Ss6٫=tQO۶��%���<���Hۚ�MԷncׁ�.vr�gN��i�/Ǩ�¼4)�_Z�Ǣ�SQ[M��9#,s��s���z�6Y�Z�d�Nv�o��	�C���Qr�)o��7�Ǎ�`Y+�>�˕_������4��S�y�dXS��N������Ԭ����#8�
q#w::�8P���?���k6�u�!�	a�
��g�gۆ��߳[ڎB��D?�üm��y���x�$���bp����ַm�>;��/>���@L���<��|#���>�bT���g[kM�p�f��k���@�V�1f\ѱ�Ya�����F�k��U����9N}�{���E��R�n�<З���i`ŵ�7�{�
�)�H��0���I^F�|�.--ɀ�9Ŋ�㡬�L��22����qi�hX�	�2�7���c��ϪM�hݺS>\E���sL�=�.���U����FW�c�C"�v㈄�\�R�2ʸq����~�=;�{s��'����eA�L��o��m[����?�=��$�Lz�E�����f�e�=��H�x�\>&f�q�"�5���E�TbJD������~Q�$����}�m2��W���^�{��a��U�i\ENfC��=���B�е*�sU�)���%w�i�]���x�k�S�Hv|:3��ʹ�>���'I�"�%)<KA����n��SR���g{jbe<���jfYt��y�_^��o�����w���ف�j�I���7�:�n\Ż<�[/�&=	�'�$�L@���[-x�QIe�y�{(���{>Oai9s�Kd�'����\¢���^��2�~�� �2	E0 C��9F��V�X��f�ɗnZp!�	�����e7�u,���{�L.y�*�e��-ܹ|����tF�v=��������U��8튟�w���L��Ċ�5-#��=�2\[�����X���^9���KD�K����]�R�ٴ��v��I�kʳX�藓���l�6�D�J�Fì�!(U2a��p��C����LiY���Ip�����viU��LԷ�e�+8�!I�` }���5u�<�GJ����RVa�г�/,+e"��_X��]��08�(�;��@Mm9�N~A���h\���G��a�I�����L�#���%r�733�ŘD�%E��*(%5��������L�)iXϾ�;�Mur���\�V�b��c�d13>.[(���T���I����μ�,�_\"�P��[������Ꮢ]Ŕ^$�4 �EB���u_�����p,�B��Z���]�r�9VC������j����@�^����?��3����Ơ�k|��8�c"'���@�hqC����2�O;Z����]�޿'?l�dZ�H�c5iI�)��"٤������fzGf���}E�h�p�Z,Y�rg�{�&W��L����#Ǩ߼���e�)��`��ŹbLh�R���:��)<���z:�R�$��W��LAq��W{'�}�w�m��bZ��c��Ä���etp�s'�C���xaa&EY��'Mj#öEF�m���hZ�Β*�v~����D�8����h�1<�0y��y��$��,9^PKؽ̉���>�*�;v�c��87+�Ci�,,��s�!�I�Wʝ�#���o���z����_b2�I�.��_����q�?�0=���{%l!�Z����k���/,�_PA�!��2�Ǹ���b�9,�@3S�>�=Ks3R��q�*j[0Z��y�+g��~U%+� �%e��f�!�]��(�����L��{�=�apf��?OE��
�@H2��Stx��$aLLw�-S*u�@�}���R��*�3���1?9L]i;��ʗ��bᐤM�]N����q�fX^^�c�I����t&��tq��/�/���z(_�����[���[u:>�o��mͼ�ws�}T�� �Vt������Mfv�#�O0�us��W	%�X��8�8�3t�����s���a�2����lU�gɪc�ICc]��;8].z���]��)qㄢj7lB��N8�']�fnb�O}�:�Cs�U
;��M�^&�~��V�~���@�6AQN6�W���'H�k��JgqnkZ�之���N�܌�̳��#T��efb�[�N�]tp��nl��k?g��亠9�f��\�ލ��?�/s
�Q�A����5a[��;2ƜÎ���\�@/�N|���8N�eR*����a�d22<�ݛi,���M�f�<r��8���df%%�j�+���y�{��E��ūo���xD�F������^$i�%��:c�� �|�=�,�����~�/�Fba�lʈ a����=���F�B�#Fݦ�"�$n<�g�梩m�֬���3<�}Y}D�m�4�k�ҥ���	��ވ}~T��E(��\&+'w@8�b8=KR	[Z\σ{��}<�&���C/���̉��:	{C�my�m;�1�m������-=�|�ZL��.��l�s�d#��(�oF+1��މzFg�5���O�-DC!,�8��?X퐗���H��]���"�@�^�q��Aq����>�jKQ��b:!�Leiم/�/�´���d�@��ɖ����͵���|W����}/280F��`�6F:oS�c�p��Q+��T����1E����O8{���<�i�s�~�7���s�}z�S�|�"�Ü�Ǯ�� %����Nvmj�3׃&$#+Sf\��2%�^L��$5%%�E��Ԍ&<y���װ���]�K���Ƿ��ߣ0�iT��u�gji1EU����|3�bx�Z]��_��z�O��������D_�)��DHPឡ_�U�"(!t��D��̼J**뤎N�O�sX�ù�L���\��V)w�j�'�QR�Cey۶o�xF_X����)�TvL��0Өd��m.}�������{�-���-b���rD6��%�eE�dX��"3SH��C����BJʫ(���,�H$�Q���+G�ͻ�v�N\���d�Ozx��o�nj�������,ؙ�yyC��+��a(+����R��\��1DWd'���/x(S��p�ܪF����\JR2󈅽h�q��Ƹ|��z5):-��r��l0�t�$B0 ���(�KK,�<4��@��-�Wnժ�y�ۗΐ�l"�3��O�ǜ*��a�>��g,�Γa5�eRȷ��t�r��F�d^f��f|��2%�/���FX<,C����"���-{PײY�'D7������<���@Z�2L&L�5�l�Ԃ�b�U��'�|��i�j^G�V1>��fRq�8��GئG1'��Mp�7�9�=��c�4����!N|�y���ZMT���i_�����E���5j��M��U3<<�̒��D�G��0'O|���8�H����l�E|�H���dl#���c})��F^�xANN�*�����T�Ƨ������T�Ӳy���&�!��C�?��Ќ�덟�]R�mn^�)�c~bmL��B�m�f��mx|n�?|�ݮn��m_TIm}��kY�	ǂd�TL��p��q4	?�[Bzbq5��_���03��&�D���vƞtȟW�)IB�B�e��ҩ,+�63'�9b<9������c�+��^�����7_�<3��=�5��a�Q"J5sK��w�GY ?UK^zz����Yrre�]���a-�c3�茌�͑��z��o�CL*^c���^���;ƴ^��_��U �n�/�eb�!���� �p�{�.�{I5�h�������+-{��O��3�`��c���or��2B��Kt�>�I��q�CW�sy�Ϳ M�d�{E��ecr���u���r ��"��������!�(��Fo�d��܍$�Z��!73��;�d�S���ky��Ȍ�Z5Քa��dW[X�D��X@g0�>}B���
y{�4Lϸ�c��y�v�o^��t7�N}I@@UBq�6`��#����]�li�47���\N�P�$��0��ݸ՚&U��#3ؼ1��tNPմ�֭��*�Ģ��?|�,N<��0IT������ /��D���^
3R$�ܤ���I�s/J��&L�,P߸���R���|�����.��)�m��:�����Ǭ(�4�Yώ/�����bk[���ɞ�y�CR�)�Z)�ءP�M�v`����嫌�;������;��i�g�HI�F�����oP��F��Ԗd��,��a�o{�Ӂ�d�0���

�$��~uws��[�լn�e�N<��v��+<zp]R�	a�r��AK�8��5����*VD��{]u��lϖ;z�>�(�o��g��J�.H�1�H��#a4+�5,4"])t�����"�����hyF�3�	<�>���k��B���V���Kj֯���K���ҽ~�_K<��� �f���=���35!z���>�%�Ҿc��p���IOg#�=x��R@ R�^��5�9���\Z�l�`J�j:��� ��I.��D���qk�표w���23 ��i�{����!I�Z-E%e��X���T�"�,+B�'��Z��`},���_1:��*�;$������5�x*��J*_g'p�8=�����M�b4Q��-ӧ�&\��x�ߏ��nmcM�f�#�b�	C�̌�>cFIv�Ř��ќD�픙��9�}l CR���,fgg��-Ҡ$��Ѩ�?Fq]#u�Z�,.���T�u$�?�_��<�WPH[��G�*D(u%Ϝ��.�JCq^q��Y�k/�@AQ!�X��O���a�Ϭo^ˬm^�t�4�����}~rDu�Һ�{c�����Nzr�����8!��L%'3]��n�BX���zQ^~>e�e$��ݠ�@&Ȳj���?0>1DB�����{_��@Q�4��rG��~�AC}u9W/��>3+�5"=�5%��
xMZ��6�[Q�'��2d��M�xsX�����_�0�Ȫ�X(W�����V"^�۵���v��Wǿ�4��㪺��ԯ&�� �J�$�$���S�W�(�.��װq�K4�~�1GXn�0٢��÷��M��J6�����uT�
����ǽ�<!��j8���>z��{�J��ǿ�'~�q5�[�R�~;��
��v���*a���>�V2�����2"Ms;���a����g�>�k���d[����k����h6I����o`�-!�b_��I�-<�9�RH1��֋I���=�����%��W��?P�~m[��h1�W'�϶p��q:��%ͤ��a�F�����K�Ɯg�(�^�_=IMa-M�d�g����ё!*J�X^Z��q�(��ev�íGOXp�QݴF���/��A<���EB���oH�/��0a��)̠(;����dNԣ�gf���SR]ΊB����{���y���}�(i��xG9���x�Y�$�ް�}�_&���c�?{������n
r�Y���ϕx����������_�ǽ�a�*���)�Exc1�;N�*8�����#���W׶��{_e��b�K+�\_I�ZVKժf\f���y�����c�r�K����Ǜw21�f���(���D�K�}��P7*���uml�{�pLɽ[7�M7QW��oi��j�Vk�J�^�xUb	��L��,{#L-��_����������ç�C��2f����S������D=4��{(o�i�zfg�%�J|�,�@��Vq�v;c�N�jٺ�����0f�I��;�]F��c�F�B��c�gV������n����'뫊���[������D�?|u�?�b��B)VIRX<�\�1��X<N8!�,�QR�˩_�*Gd�@������*��|.O�gjb�F(X#���Դ���|�����!M��⦑��ؓ���2٭�+��w�ǔY S�ꨂ��L�����ׁmvJ��D�B���/X��Cx��.�J�!P����c|.;!����;ٱ� 1� �:�
�J�ky�H8��������	x��!	o�N�B�sD�%�hU0�i%ʵs��~t���FP싷z�`"UR*�
z�K8%I+��c�L��X���qm���F��b&%'���RJ�j�37U��3U����\;y\�xM%z�U�i�Dc14J��� �si��� l�I��N���"<�$+�H���>�?� ,S	i��FB|��?ɟ�H��m�������Q��r���X��e����a�SV�^|� Yy�8!ٛ5��]PƌMt����4̪�\��}�&�b�,�@ �� 			Єd�c�N��Ǝ�N�o?}�t��77�?ם���v�xvlk� ��$H!�y�*��ԙ��w�oo(+���y���ꜽ��}�����n���:�"��s�����訴���0߸kn�gL;		�y�z4�hV�ĭ컀��0
��:;1Z�i3���&M��k�,ƴ�31�:o�A߹���O���,";��+n�d�Q/�L��V�)E�J�� ��o�������Uޑ\S:�b{	3f�ü��5i
FZ�n41��Gc<���۱��A��0w��W�;U?e���mE��?%�ʬ��
Z�1��õz&�Ĕ�0a�T��l׉!��z������c�ӛ��G9K���w���1u�z�6mx6u�-L(���0�|u��F��W��_��/b��Ś���K[���� ���\�T�Z����Q���Sx��? �M p�5i��/���@�\D�q��8��>�?��(�c�R�����,�O��m�t�]�Q�h�Qo)��C[��[[^F{�xMf|���������b9���>®׷���qt�W�^�k`�5\|�s���H��9�|�$�_~3��MDY��H��r���{�᭝/�T�j9e�g���*\���o�����^T/Ǭqi,�5E�`��o��ٳ�ݍFmgϞG�ՂZ���#'�bʜ����f�ȦR���f~k*�'t�M�Ƣe7��m\8s
�N~�K}瑣�@������.��?q�<>>~�OS�&��+Wc�M7!��}������w�a�����{Qo���:���oc޴n\�p>ҩHj��A|���X0>�����g���/�|�,��{B��*d�M�S!��71t�����&!�kWߧs-T�)������}h+�a�*x�g�>�\���ƒ�׋DCr��o����Sfc��c������ǹc��GV�Y�>��z���㽷��53'�ԫ���#��l+5�>�#�B�,~x#Hc�M�b��K��Y��[��?}m%d;'`��_�C?q�c�}�>�Ok����8u�#塌/K,��w��W#��a��]�����8��P7	�l؄��3Pm�����dZ8��UiOp\k��[��d�
5e��7�L]y����|�o�����N��������$~؂�Ja���k�b	|�Ȇ�Z(wM�+נJ���;���/&���Ud�l+P�D��R����Q��$���ɶ���ƭ�|�����/����X}��6�j���]��9��MC�8��ӞX`6�ZPn���Z����8�2-�    IDAT)aK�1�k���'d��Si,[���-�gE,�҆|��j����3��FrN;��9U�#��J!d�K+���m�3p�5�z�Y|�M��i��k���~-g�&��r�3�(�%��RI���"1�ϟ?��7C�vW'�m(2ke��,�<�R)Lnk��׶�������v��?�J�ƣ�b�Z��,��-��fs ��*�� ���{��9g��͙B6���t�-���<��Ґ����r��y�����g�3HFr�O��&}��G����j��:S5j�D��q�H������~�o"�N�����]������p\�D�)�.M6�c#�8j:��8��Ã�oJ%��i�f͙��Ӧ��K��l����>��٬��v��+�b��w��u�|� &���l:�|N�jk�`xh �ϊx��T���-6~�҉R�ã�<8�A�o!�wv��}O>�.���6���!�=I���JE����/�������I l"e�SQ1��Ub��D*�B���l?�Ҋ���f8ih)����羊��V��n��HC[>���gD��Zؙ��b�uK�`�LJ(��?�қV��7c��T�%�A%mɡ���/1z�l���Y����$\}M�b�g��,�N����ža���I�J�q�8�_��ӧap���WC��1��ǫ?�	N�H�3垉X��G��3.3�(��C���B�?�6.�>��1�\�ُ�a��	�4m��Y��߈��!��&"V�Հ4�Yrp��-����(s�l�'SF�k�����K�a`��|���!'ӕ�*�Z9'�C����3�U�q�*�64<��q���)3p�c���)������
�ڎ�vv.���џi
۵f͘��ǰ��g1p�3�L�|�p��Q�I�@�M��1}��X�lJ�{�{_������Å�Ø{��X�����������w�7k��T�
��Â��g�{xyۛ�
]
*�`�6
����P������S�	E�
V�~/�X?��z#�8t�38��G8��ADn� ]�a��|�$?���p��E����,wŪ�1q�,Ԫ�������S��-�,nX� F��3�9��>:��Ձ�mI�w��kQ��DJ�{�}��u�V��C5�^z=��p�����4>��P�L�4q*����*�z�N�w ١3�7��,���s��ѣG5A��g�C�P¡���Fh�����K�X}�øv�DN^��<��=��5M�tВHe��ه.ݘ�-�I� *���7Ο��ݵ�����_��������_�p�:)�i:?�����B3!:�f�z҄�s�58�͕F`eD��(�J��#���!�����>��p>�}V�A�������>�N�%[�R�E۸	���9��k���o�8�&|�!��mGze���щt,鬈P#������@Xw�u�"3��ŃҠS�����B>��ᣔ/�w�x��iO!��i4�#W�I+��>��|�T���_ߎ��C�Q`1o�b���a4�.4BR�1���f*����>iY3ۤ�n�>j-W�:ۘ8_���`-+�ő����ۑ�ea�KXw���완�zM=ؔK$̙ͱ��"*dryE��炵~�h�C�҉����<��4N��oyY�H��E��d�jp�5g\۩R�i��آ��]M�jUGQ��qqd�b#uT:��� ��	��ĭQe��<���~ �Y\{�J�\s\����}!7��� u��)�"L�V���v�2[��	_�v�ZM�d�2� ]�rh����-��b��Xv�\5���pN&�ёa��D�뿤@���]�g���=�����z
�̀*�s`+`Ǝp��||h?�S)��,ݺy�B�P.��{�{�4*4�l����i�:�Hu#���QǸ22����J�#���/�tXG�	Y��">�{�r�b��4l�Ot)�R_/�錂PN+�Lo}dmm2T�r"'�cg����D��G��9����}��>o�8c6����a�糭��Qd�@�]�������6uN��Q��]=��~ʑ���,G��N���'?±];��n<��_�D*�5S�S!�m�m]���sg�N����!�O�,��3��P����h�LJ��Ԭ�Ж��on��/>�vp�u�x�x�{>��@aFZ�Z�`�ʘ�ꐐ!���n��
rt����?����+V�٫k�$�:{�f����7��W�C�BTX}׃�2g!�lQkӕ����3ػ{N� ��@[��z��}W��0�?���YX}�]�9wj~ Ȗ�x��Y<��DTF���U���Oa��QC=���؋-/=��'>F�&�'@w[�.�i"�����яO�‬�	8�; '�E&g�%�bG���}��QcI��u�c��0�R�>D!r�%��c�>��}o�j2X���YRY��XC���C�0i�UX|�rtO�JR�>"t�<�O����FT����h(Tʈ�:�߽�����\Y�(q��y�J�<�>>����8s�f.�+ׯCy�4}�R>��<���"
���p�����W�m4UB���� �ڴ�n�A����;b�O�;�{�T\��ϼ�:\w�t�LV��O�1ZBƩ�=:�Q
�p=��s�Hɼ�=rR�I����EO1��_����v�F����3s�������8֡ӨD~Yz��}��Œ2֬�����2�*Ԛ
�64�H��C.���ՁZ�*�s�{�A�C��Q�h��P~^+@&��F�1"L�N��f1���L�A�d�ȳK�Nxh�M��0��\͡�"el��c��j��B)�l�N�:P%��[sZh��>�t`��z5^K^3���y�>
� V�ɈUZD2��q\���v�؊#GH��Ѫ���ᎻD�*"p�������[P�a|��8j��L�$�d��0%�<�v�IYȄ>�fSƞ-hd�r�E._F����X�hU�Ii���e���{�L�vr��&�%�-��_Խq�y�~��u:��$�!�1��� -��o�hԆ����X�!�Zf����sp2i�|�v�J�Za�V���� ��knŲe+0a�U�7}�>�/H�5U�2�D�24�5e�$-j��P�r�~b��"��c�U�zH�{1m���:�6<fm�eM|��Hf��1\F��F�YA�����T�BGf�������ή�/�7"�&r�2��"�P���֬��H�2B�8����V����FƦC�~�k�[�01����*Ξ8�W�~B�\6��<;�G�ρ�4��A�2�,.\�G�R����
Zd^�'Ć}�t��.T���d4&������^|j3�C�<W��VI�^F���=a3h��Ô�xA ���gIs��u���4ڵ��;8��-�F�4<��g�l9�t�%��pxȦm��������r�B/&͚�̩E[�� p�(8>N��/?�3�8Rw��l���3��/�.�NF�[�4�Ď��i����'�S1��N6W@Ǹ.uutO�$9S��Y�s��D�ٶ���h��E!n��1c���e�t�J����ܩ�������^,���>c�հ��<w��3��Z�'�����sgTJ��j��4#/ڐ��B�(�~N�	�Q=TJ%H:i�\}��s��Ց�FL�laN�`Hq�P�9��2V޹	����j�t�I���uT
E��ӧq��I��=�̑���#�'g�Ϲv!�͚�B��UD�rG'l�}'>�X�rVl|�>Pm�1������'�^IfϺj֬Y��gN����8~��̾7��=WMA��󃣘�=����3���&V��26��@i�4�2��Ն��q��m�����_�S��ػw/�y�9�<sV�	�5�.j���Ѵ5v'�<ˑ�\�\��{�¯�����}�]� 4�2OY��d�it��)g߾i�������з;;�~�����cc+L�R��i����!!cӶ6����֒1�����R�7�fT�y�y�hdC/T� ��4�c��������"'e�P���ﳡ��E�"�>k�
����6c�j"r��3�%+Вv���6[r<|��f~3FzJN�	���dZ$��-�����\:#�v��1V-6J��yJ�р�QV*ka�:H�QB�.3�R/oy��51Z�b��Ÿ��O:Y�$Z�`���Ѭ�����u밙�"4jJ~������������DB��x���)�vZ6Q�PA�~u�M�9)z��F�(��Hy�+�1K�С���E�\�lAAS&Hi 
>����*`d9z���CG����뻒|�h�J!4�^C(5뽖Q���w�I�����P(TtH�4�h�8~�
ۅ�YA���Ȩ�Ữ4���B�	1r�Bk��<<<1h a&�B�����(��2�]�v){$�wΜYH�|i*0�d�ƣ�l�2��'X��
eS#�ύ٠���B��	^e��}�u���~%�]h
K1�#�N�G�Y����0�~ �aq�[&�R��w��́ˎ��)��/���^���*C�*�4���=�<XJqp0�j��J%2�����,eW���9�Y�dOxr-���,����"/�� �e#��˔�����\KC��\����b�F�VY� NBT�HӜ�^�r�3Zk�#d�3��I\bF����!p�9!�4��+����9�O�ˏ��<�:etM��~Q��Ȗ
BEx�I���Z�c2� Ҝ5/����U*�/^7	��:=�w��o��Ӡ��]_�#�̘��&d�{#5%l&A�4n��u�9��|�H+�"*Y�"������3��!`��7o��@�Y�^���ti�|NH��pkJ=�lR��0�WhgPkE�p�=��EZ�_G�kh8����P.���X��~L�v5Z�,��<C�-������)��QP�_�N��Ӊ���H)PK�ղ`�s
�r��m?�>N����������Rü/��Z#�,g4�B�Ν>��gOi�iڻ'b�܅�8a.�(ww��e��m[��3O	��tOƊ�?�r�x>��R!:�i\꿀�K��=k.�q���5tL����˚nZu-Y��5��+#Ŗ4�6�G6����_D0ҫR����=�L�����T�>@W����쾛�O��m\��7f�[�����=�������T=��k��-����ޘm0��}+Z~��ޕ�6mZ�Xnӆ�a���#�Q-��8��=�а�?o�C�]�ƭj(���!��M�j��p2�J��+(�	k�Id"��7dOn����0C#c�"�1X$�^�X�s�y��:�7l(c��!��J8/Gr�(���2 �,�thÊX�M��+<��t��es�"v�ى�;^��j51{�<<��g�F��x�ti�-8�Y/k��.�!i�>�Ç�a#\Ӛ�*3�<���p���ؚ!g�ё����&3;*�,8>̴���9�1�Z�>�QX�Т�t�ju#JS'��d@���C��
i�-n^޼c��(�FH��1�jZ2~�ff�t�.���DZ\��@�N#�,����Ͽ����`p����q�t�8hj�\9�Qf�Hg��R2� $+���^K�ά�P(�'Y�j_���3�u�**QD)���R�ÈF�Yg�^@�c�(�J��Eԩ����զ6
Nn}TF�HI*� J���Y���Xl)�BG|��2���b@�`�Z-�V����s���q��;*x�������bɦ;��|�˰�.�AZ�JGhxM!(�J=F��L��7��)�ɛ����!i��pM���2�	f5�i4\N���jC�����%�,�4�u��ATܚ��@�y��R�):[]!P�l8�,��0�[2M��u�a
�zK�$t4J&�,����/����G�!���p��,qx��R���#��ғ�@&�=�Po�0n�l���s�K]h��ϒ�)�U�
�6������mlD��1�s��	�Z-�Y����A�j`�:�l�4ؕ ]TwE%W t�`��0
]��\���$9M�Lz�f*{��@%4�O�}���Is�`���:��c��8�@�(Z�(�S����!�/W��}�A�bȦ�~i����	�tV��X��A�X����6��W�4P�/��'�ٺ?�Т�nN�IU�^WٗsM���	O-����Yt�j�����4ʕ6�ý��P�ܶ"TJE�wD�hC�-�.U�����s�0R�!�1=�������~Ee�ոa�"4�r��?�����)�jT�l6p��yi?��9ƻ[��\����%ڈIYȀ���Y��R9��מ�C�N���z�ٖ��9k,�Җu�ѸRz���3��[�������O��K�}�T�@�ܬ��E���k��s&F�y;;������`�̫��9c����B�Ԫ:�Ɋ����s��!F$c1�d�
���@Dk��N3��I9$�e�l���P0�1�C:;����v3Yr�����][�(�;#w�&!�G+���Y��4Ƅb2��)��cVC�DGaA�� �//�a�0Є9+L#f`E-˺2Gβ����� �h �<�$���P�FG�>��`@D�?���Orבھt*2�^�����3��"��[4fd���BBo��7����ҽ�K��10q�,<PDhv*z¬-��(���p�^��\�A�w5����u�^N�� ���frR��R��1A^�~iHd ^'�
;���&���f�S�ry�ۏ���O��3f��5kq�Ï�s0i��E���D^�Z�#�/c�@���b^�d6^�)�F}>#�2f�i���f3D�ߧF3[p�:��D��(SL��7��Ty�R����"���(�'jeq���r�!��T�����|&�
^5�:���&�A@�9�.݆��h �b	��U:
V�a\8�?�s؜:֐.e8Y<�� �L�e�صЂ�3C"Zn���:�t^��x�z
�,��}_�.��Y����r��ܺ�1C4Z�L^@����(�PȧE$e�@h����&�ȤLi�F��k��Ut<�=��2%4��g�f��;�)�A�,�}��"Z9�4� ^]��\S:u�4is39������yL,l�u-����O����U�'�5k�������b�� �����T^��zr���J	�}�'%kT\�.�w4��r�
��ut�;u�1��������%:*�σ�m̒�[c��5Q�]�1yg	��5U�p�u���Z�,x�	��3Z��I[�{"gr<��|e�$pr@:���.���wq��h'����!�Z��F��F� �6�F���D!S�Ic���i��0��B�΢>���t���4��2R�|�}���zhԫ�� ,�7-�BWG��E����<h�`|W'�v�CR$����������Xi�ܥ��2�GA��{b�,Q��F�|A�Ą� ��O��Ј�/��i2$ێ�L�_�j�ٶ��z9ǵ0�s",!�f��A����6z�S����������on[;zt��~��7.��m�ȱ�V���W縺�;�w�#_ر|ō[��L�0qܤ��r�?04�u���#��n��Mv6�Æz^0��qf˔D"ec$RQ��F)������`T���]���	1�{�[|EYH�T�u�pQ�X��Úߛ���|39S��(�C(��z�HCC�)q�c�9 tFn����ZL�����.�R6�0�
z��-���
ZR�X�m���_>�={�T-ī�ش�^\wU��6�,�5�(j��`ZB��nK}�^�7�� ��b�F��aV`��V��/��D'K¥KH���D��vd�ȌW�&K�[�4�3B��	��IK�Wg3�����ėUVɺ)�7���An2���p#_��t����.n숅z;��x$�#�F'?\��?��Kh�����^�>��G�kʑ�a9��fB^R4��4U~�����9q�(x!��C.�E�YQ['k5�s�3]DAS� ���ѐs6qVh�L���dnK��ʐ� pi�j��3����3t֡�2Wv�|='�0|
"gY�X    IDAT,O�ɝc��7e*1��-Rw�,���=3Y֦G���G�A5��rG�l�<���8�����?��Y���
�n`�5�x.hy��8T.�z.q�"P-���"��ҵp_x>�,�2�S�9�>s^;k�%X۫K4�+�ȒM*�G#E�@
m���-�M�W?l����FD�iة,l�� jG��'�E2�� �N
�2U�Åz�I��m����V[b�N�Qk��Tp�셸��Mh�ܧ�!����k�YN�#���X�x���&:�B	�zݠ���H�@{9��'�A�o�����,��~e�m�$,S�g�/�e�H�P�9w|��ly�|�n����	aI����<�fz�I`�s��Gt�)rYTG�����n��	Q,WԮ�Nr�
�+X�ƍ~���2t�X��S�������+0u�0E�SJ�_�9�D����v~?����t���f��T,W
���(�TQ�u�\,rpRhUt�����2˪�g�^wqi�g�Mϯ�h�4�����2�c��V�y��6�1a @俆�F��ua���&d�Q,bx��g��2��k<�����C�z���{��B1ˮ��ۍR�cX�ArT՜|'�K����]��^9o����[��F�����������e���Y�ʩ�mG��h��뿵��[�.�r�3X�(ʾ���~���|
���0��ך<plac(z2�g��h��
���2
"��`m�J�VY7��^���}�0�j�)e�R�1�f�Gj?��0e���6S�b�ô<d�k�G��ś�䟸�L}CH!�,�3p���Y��I��D__
�6p2����OLX>�z����/~�QZ~6�������h��Ẹ��	� �L����f�;3G<:+!$:R��N�BN��.4���1�sHjk�g�A���cX��#t��Ӏp���~R9���h�2~�@+����9�d����@T�'���x��ױ��*�tv2Si�w�K�0a�A/��P.�c��7ABD~@C�]��k����|Aм���!���1��=��d�)W�p!,>�x�0P\O�b�p�1���{e��Qk����ڛܷ�Ĉ�ߓ�Œ���c��Ek�r�1lEUjI��B�!�uX�5��0/�B_�����z��,�X.#���{����Ъ�����Ð5��{-nZf��dˑ�����qO�煾�cPq^$��=�<�Ð���	�Uf�J��H���#�;L홐�yS�J>ߴP�ܓ�d@ɚKg��&?����4��7��?$�i}��,1?��^���oV�4ti@��y��/�#�yT��d[���VY��!��l���̮HZ��zP�Jg��0GM�	;Mt��ܙ]��A>�Y�=-��PuH�K'E�g�"M�>���Xw�T`�P(Ă���h���3�w�><�!׏�����ۜ�˶�%�x��x�k*m%��]l����0�f�b����_C�4);/�B�����bN�l�Tά�Μ9#��؆�u��7 �:����/`6+R5�7�K�5Z>'�RIMA>	��AzM���F�'g����:�VӖ�\2Q��s���y���Ʋ�L��=��P%"#1[6�	5r*���)g��dE?q�ܵC��*)KƧrN�Ør��MԨ=��&u��~�������F��¾}K���o�7�,�TO-�v迾�yu�M�w-l�:��7H�E���旯;_Z�J�Z�n�aupcn�-o�ƒNw��9�z����	�Ԯe�M��@{	��l,a؃�CKz�y�r,&�נ�J��Η���h�)��Z��˛�$Cj�{~�IN��{�Mg�>n�sk�)��:���r��QF�<��d�9�9�h�=�K�ɗ����$rk6�B�]M>C�9�cge�7�}�ӧ��T�>v��L%/S�YG�A�x�s��in3� h�cڜ�"G������;j�c��٩�A]x��xx�
T��6J���ƭ��r�y�Q�d\�8 H�3�Ԛ�Y���ǎ;02lڛ��w�uf͘���Ƈ�����ԶB8"%d��P����M�J�92�cP�^l��5F��6���O� ���!����Q�!Ο��CG�k�4U�c���؞)������:d�h OZ�9�dؒ�G�l�w�MYA���8��{��������S�9��$s޽a#��Y �_dUǆ�
�FF�}�Q�p_����'�]N�g��o�l�16�o�k03����Y��>���H�D!�:��&���g�l(H��g`J%ɟ�Y����d\���[�9G����������5;u�~���y2�����H(�[ך�MU�HϘ��!��$�ҩS�I��7���<f{�a �mV�1*��˵����1�����@��D��~&��ٵ�]�I����:r��j�"&9�V��4����&�J�ۋ�g�g����y�Q�3{��󵗱uۋ(W��_�p	��aX( ���0q���� ����W�=�O�ЍϠ�M�+	�\9�)��u]|r⤂Ζ�Z�;p��$`Qp��D��6O!W4���/hkdI>v��$��,���,�_�q�<6B6Ͻe㵲t��n[�]3%��m|�ё&'"�"�Q�GX�,��\*I��g:��;���{�_���u�C��+o�|��7�����pr�
{W.��_���/lk���|�S�������oz���_kx��Z�%�Z�8r��EV���K�1m�n�ԙ��8�X���q������HpcFkx��:tnf�rאR���ѩ�[d�S��u}2ԯ8t^�7G�(����G�q����J�7�7k%�9~Fr��ߎ�.eo4��!nX�L";�a�R�����h��l�����꒣�c�Z����0���3z���8;�������0�mk�Ra� ����>[��8iv+�8�����u1���t�q�E)`�p���;h��$�uc(A���Hlj�69r�|����֐��)?;��Ƞ�K`;l�@mdX΁�H�NH�����6e��S�1'�@C��;��ΟF�Ւ��1CWT�{�y0��CT�eܝA��=JG���2�4��,� �,���Ҡ���j�1�h6Z��1!�8���N�G�>VĔ)SP�p��k0窹���U��H���$?�h
�?���	z��N�>�Y����q�"}��B��y֞[h/�+�3E��pXҊ�+�ob�$%�'i+�=���x����\3�g����A�HF4�6FY�Ʊcǰy�f���v,��;��ҥK�f��̓,XJ�>Y�7�	�r:}�4icD>3A�ʁ�C�5p�g��'��,9C��Và�Bø�`��8���i�(��;�>�W�3Ƹr�&a��"G�{S�{c#��e�L� ȼg�e6�ַUZqO=�8>��}T*E��u������؛Z���-{Ӕ
�������֯��7�ĸ$j����ɡb0��a���lDԖݜ[��p�Y;����4$Hh"�b@�gA���Yz#��u�,i����\��&�x�s��$��ÔTx�u�R)���|QD�ju��Y9x����j��������T�����&�e+
`�M�ʥ����%���ɟ�}ǡ+����I����nٵ�o='�@�{t�K����]�n�����?�Fc��u灅�����zc�P�U�fV�-8"^`F_!U�:q����Þ���Y͇ǚ*.��D_f[�HQ\���Q��_e�+d����k�_|�y�@E�	�}�j��B���A&�3�"�I	Ɂ5�]b4蘮�17�p>�w�yG��$��e�V%&/��:Q���Al��m2B�rT$�b�C�VS
�c�ڵ��_۹SF��P&P��&�k�΀`�+FQ�vqФ��a�
ATĐ��N偏��\�i��$za�=�1�A����q�1c���p8.�r�Eb�3&F�4��l^���vٲe"�����R��$��IƦ̊�}�����{�Kk��y��i�lf6�C��M���A�!�'�o�ˁ�؟c����/;W�R���K�O*;t�/y?�9C�!�A�n�`֬p1;�s����!D�ρ�CV$Q��Ae ���Sf�Rj���seL��{M#,�6���x-l�b���2�7�<�y����I_V�_6�sl�z.:�Ke\��!��:$��
��z�wR&��Ñ�B}~���혀;qҚ�(�)��a	5�:C�{� ���!����w�U��u��Ӿ�wy���:�|ou�С��Tj��+���:�,	��K.�!�@��KOL2dpN�$���<6�%���� 3n�7qw�L�%���`�|�'�{Rrк��K�݌�,��\��"=��0"^��%ɓܻ������я~��Lm�%�]��>L�4�5C#�̀�����?rS�ަE޽b�.G�W�J���A�q�q@q��� E7(N��h��,$dXS�	�ǒ�}d83v����]d�Y���:�}���NA*�Mָ��.w!�alm$N�;9`�B�B1:�©E���d�u���94h]����;r��}n�úu��u���lX�P!/��>�dDwb9�{ŢY_���{�����п���wn߽�oj�?���ΌU�~����z�u�X8{�G��������ۿ��o��cg�����A:��]g���^��+n��S'���W�+ʍ���Z�J�<�P�p$g��yP����+�[o���s/<���gd�@��j�j���Cg'���X���𵹭�O���֮Łw�Q�2{�%p��.Ae2d��`�@��Yo�C�a"47��r�FOal�x�n�u�Ѷm�����}��7w��Y�:]I�~�ؒk��2-d���yD���-[�j�2d��+��<ˤ���Z}h�9�a��L,�R1̘2w�y'�}�!��xU��%=c}��5a�u��Տ�R �d�Re�ZX����&�!��Q�
��ZdF����+Ūs�n�S&�t�}�q�>�dbg>֩�g����=��$b�����˦E�mf"+��[�NA�������
w����z����1��X����B9B8�A� �d��N��ٳ-0	�������5�	�(7߃��r�ls�x�r�^8tPY�H��
���j�ç��2���2��_�b��^�&k�1�j���	x}b�sK�	Kq�}�Bۑ��=ɢ<'I�MG� K��1gG�3�}&���K�3� ��}p��x�d�S�O�swb-frD��6m�l��)�N�X,+�R�0����y�wX� %��АYsTT����q�鰑�qp����"r:Tլ+[�>�,c� �Ac�m���.��6(��ˏ����������O�P�Ω��u�l<���$�uN�0�]�l&/m����^I�c�B�Vq��2�3�cK���3���*=�b�O��# eB%�!�̙��:yo���C�I�QMgP����Ʀ�g $�ƾ�FK��+�c�����S�� ���i�4�i��$zR���ԱR�Y�.��}��{6~}֬���e"�7��y�]˶����rפ�#A��$2�	x�P�z�+�7�.]��/�r��O���G�����{卽S��[��B�oݲk���׬��I��������FQd������;����([��R{K�Fv�z�	0���W���'����f�89�d�	4�L�N�7��*R��d񬍭�i��}�Dj`�$��f��:1(�%�[�xw��{�4�U����s�)s|�����;��>+7{B>�fqضEp&%�nnrgc���2s\n�8f;����6l��Nm�g�#U�JIE������7�Y�A'56���o-�!=��#r���/]�$N�K$#��qF�sBL� ZWr��Y��� M7|j�>�m;^5jSq	&y&ӓ��Aa�z�]�'�l8n�8�9s���6'�<=�8*��G����b�?���UY���#�����Of��Φ����lb���Y�y��֋F�g�5�g1Ǡ�V���$;3�(��s��``��ɧ��A�Lb߬�30���kx��;���{�~-� u�{sO3&R�#��ϘL��� c����@��Μf5Xh/Wp��M8w����2Ae�Dqh�[�M&�!'b�Cמ���K9T�E(��Չ����y�g$QJT������$�q���3O���8��]�`�,Y�ݻw+2�:/�l\�Y|õ1��q�ϯ���ղEG���Bc��-�9�?��ҥ sxpo��W�Yc�I4e���,��VO2k��C��k�Dc�!DkE����z]ˁ���s��fn$��%�z��]2���H��0i�DL�6MhY/��9��!ʚ =	Դ�,�>2I���f�;sV2�n���,��O	�tR����3�Mť��8{�<r����ffg[n>W����J}~z�P�WDnMl����[�|��::T>$�Ab2-!e�}>c;�,=�f`j8O�\"D-�ːa;qZ	�h�.d��6h�rL4G�k�%�D��mZ��rN�5�q�k�������=+W��5�+� ���s���;�,}u����R�_]��JT"��B�j5gt�_�g���i���h_v��ym��Ͽ����Z�����ԭ�����]����Ee����������W��.���/7�ft)X#��ZufL��U7�$�N��*�Y+T}E}xW2��W����&�7��H4
�I�q�]w+�~�3��V02IAbA��2�kLE0�Ɠ@$��lŲ�qݵ����Cؽo�T�Q��z)��@}{���H�s��םZ�f#�	P�h�����*��zCm1��{��7?nZN�ܜ52���cG�Dډ!LH���Zj���:]���x��gUwN^�cG�Z\��� 9m������c���I�����qj��胣xu�����8�-/
�6���L�Fmΰ�y����U�
�6Ϥ��t/3��|�ITGɟ ��F���Ds>�'��ϻ��B.bL�Fg�(aч~X��Ϳ�~�F�N�N��S��/�	��a�;��j|@$'�8��/Ǎ7.��8t�}����Ψ\���R���s+'�jz��)�Ct�c����r	�?ŃjOˡ\,⡇�0�W_}ϕ�Qf��fc�]��ӆ�ab>�]�L(�:���勒ŭ�c�*�<�ܳ�FZ<ۼcN�"�cr����5˸�N\lxr&�o�J{.ĭ�ުkg�ِ͠�t9�O�o��|,��{TE�#U$Q#x�}��ԫ��3s6�_���x晧�%aF��kE֓ӎ���+C�D����^>;�O=����Jd��Q%%�V�`�H�*@�Г3w��:���˗.�«���ȡ��r'���A2/�~�w�� S��H��M��6h�~�������&������ٳؾc�h��cʱIr����= ݇8N)�8W�� �Y���ŋ�y�޻GϜ��;g��6��{��;Y���hZ��šI�!h<�$����ٍ������8}�e!���5${IC���Qq�9�o�����:���R�xp����\2��o�~x��[�=q����l��A)�Tơ$z��i��Э����9��|��/;���ު�/o�f��`f{���_��V����	քڿ͝���������=���I�WY�9�_��9WM�M7.�C߹s��fi�b�/���y�M@����f�!�#]{�-�;{�� o��¸qg�pr�h�����X/[hG��j��/��+��o�=���ʺ)�"Con��x-dM2� ��xj��P[)2��x��+����=���$����OK|%��d�t������'��>#6�t
4X��|�AL완-[��໇t�c�(��|8��cF��ڴАT(�ϖ:���G1u�lڴ	�[�m��ߧ�z�i������q2TG��K�1�D��z�^����Q$��R��Zv��n�ݟy�aa"%�09W`���r��k��c�"7n�c�%��(�$�*)1�#x���Γ�߬�i+��Nµ�e�X��ܹ�Nl۾o�~�BNuVQ�    IDATY�,��H8����[���8AW�!�x&2��`	��>{����|2�g?��8}�4�}�ye����L��M�(��9$�W����ƙ�Z,{1��u��($�hb\���w�Cڲ�����Jy-�����1ҩ(������t�l�&�J&; ��E�aժUx����uL}U{>����T�O��[��&�D�������0R��{�fL�����ϞS \f��k���k�`f�	Z�pP����5�g|�����c���:?/����3t���A�7ᮓLɶVM{I/.&T)����8�oa��X~�2���.���!K%��ɺ�K�9�+��_L��$Dm��</B>GUJӦ�6E�'�B�«71�����������hP���58��$�]܎'�o|IBe�Ҕ����^^Q�5kVi��<����j�ZC��Ô�T�������.+ ٬���i`��pٽ�Z�O��Uk�(X|���:�l�%�/I!�J#��n�� <5o�����g�.����vwW}Fc����o}=�m�ͯl�������|�DQ��92�d�Կ}`�__7e�����������/��s�B����*�fv���;n�����އ���s����GO?��������&ե�׆��D�pFUk�ӱf��x����ē�p��h>�R�8�M�ńX6ց	�Rk�i��eD}�M+��ٳ{���{���0�5���M��;gi�(�����Y�ˮ]��׬Ʈ7���ݻ��ƨ��m8Jњ�)pk�%�N�|�Lc����137Bv��c�w�	�/�;���߉�Y�:$�7iˋ%hǔg���ԕ˘u1�Y{˭r;v��#G��]����:��Or�bB d-�mw��	��144(G�C�����s��M�bߞ�xy�v�fp��`C|�0p�$obr���v�%,iIb�����A)��C>�kx���{�
Ų������B"��=%���]&/�Y��a����ʯ7�|3�/���^|��J{��3*!%�s&0ֱ'�l|N�K�����2���t�M��[�ҖW���}�hvl��5э��U�}|�4n�����+��2�8{�SF8���u+Cg�������dVHQ&^;��j�̔������a���Y5U���t�AE�<��Ğ{�8�ۏt!'�������|ǌ�o�Ω��4kt7M�e��o7ވ_~o���!w	�K���a1�7��L�bzk�+q�Y�����A�(�LŊ4�󶵷`t����zJ�?�!M�8��Y#��Hދ�2��	s^g^�ҶIR0��g���V>��3zo�t����6�1����қ��xfK�<uL�32�Lܸ|�?r�{W	�\O�or.�=�7	4Na.�"�����O-�`R�C�XF����C�?������6S{$$�ݴ���A�yb���/'Z�{���,G�ȧ���R 5<<��l��t���(
e��zB~��/��(%,�<��q�#�'pJ�d㖧�'�9s�L�v�:���~(�D���$�B-X^ȧ�jت���U��/���/�[|(�бc=O>��o�:�?���S[꧷�.�1����/<�өC���r��������'�>���)���7T_8mܓ�-�����W���vqo�n�_~�1�4ҙb�5������R]c�.�1k�4�]{��.���Gu��>f����FS5#����k�ӑ�F��v|�WذH���NN�!��ܲS�NǞ}��o�ۨ�u�����R��,G5��KB��&ɈF�sт�q�u�a�޷����p	��lA�̾���~��1�\�ț���RI�����*���a��Ix��Oapp[^zAb-�\[M�
y%�JO�j�W �*ք*а��gF&��4�D4Ȧ��f����C2�<�|o�m�ӟ23]F�$U�}(�P��=&?2��_�M�߫��7v���|q�4���V~bxQ���&H �>ד�a��C[��/~�w0:2����~
Nc)�V�3vTW�8Í[̒�@,�����y�ϳY�_w����o��W_ۡ���	=�O�������ʐ�hH����a�D;��wm�����ʔ95LN!�:gR&�aj�I�4�z��J>l IK�JT���h��{<�������O=e�Ŝ�Ƒ�:��������!=c�+��ɢ�Re��DK��p��;q�5����sx��7q���<q��D�Mz���MA�,Ŋ��hYE.�[*��>nX�L����wȡ����d$�doQX�r�G�ߔT��8��#Y2#�@���/�;��6a��3}��S��ꅑ	��u�RѾҠ(�&h�X�1���D��^�)&#o��ƍ�V}���>�+A}$���e4#x��|\O]7b�G��%K�캥x}�x��!Sv����2��(fQƒ���M�V1�"K��xerꔩ-�;#tq������?���xy�V�FFaQ$�L#�Xm-V*T>~@17N?����X٩��Zps�93����/�Ѻ��F"y;�W�D͜S>�K=���i$�Q���,G�̙36l��{��Dr�ދ�0B._P�)�s9�:l��Cw��z���&�k���+m޲c�k�~�W{N��58�����?�v�s��_޺��:������KM�+-�ّ���1���-���%�n�0�v?E��~�G�v8��R�*g�K���l`V��� s��k��^O7ke��.*U_��ɮe����D���Y�;3�1�
�"D��Ą�ݨ1k��p����T)⥗_��#�"��eV6�xW�J8�4|���bV\�W͘%b�Q�᳇�F���^�[�ˉs,(�Ȍt	�2n�S9 ~�X�L���3V��*�-���فO?��ǎ�&)��\C##*)||�88,�p#3jBٺ�DIo�W�V�~�6��3�h����&ty��傕6?�>:v�&W5�C�CgLCD��(��p�����L��6J]�\L�:�������W�K�U�������\_�����g@2�şU(���"~�w�����޵���(������WM��I��2�!Al�4ӥ��.׉Ϟ{k���[�W]u���?���;�n�Г��<[�"�N$�;��e}I���v��xm�xe�v��mhp���_�]��(CG$
�㠒�ΐ���eH�Ɵ�EA�'O⅗^R@�/�55��H�ސ�(����Q\2h1��s��#	=�:��JE\�t����3g��֭"0�s��`�E�����<�}�8T�h>h?�M��V8:R^��7�V�֭�%H� !q�[%L	���p�^�+��M���Xj�+����X��������N�<���1j�(2���:`|I��n)�]�0C�lӳ���+<#/���5�WcѢ�:���
��^P���@&�~�h�qJ\�$B����k:t���0ʹ�,\�U+Wc۫����B��+���q˱C���7yR��?�=NW�_�_T-s1s}L� ����3x��geS���VF-v>3�R���	�]D�b[ʌ��5��eI�(i�]]�ƾ)�I��1@�*KC
���_C"�9�-�J]k(�W�}޼�r贳;w��B�]<���&	�EN������ln�������m�}���o�^E�>��ݯ�=��g��r�x��/<|�n�?i�ou��Ͽ����:v�"`��:�tt���36�tݢ�_>s���^/zE�S��/����7��-V��5��O��`��������3~�L�K�h��'75��#�%ͳ�]����8�M�1e�	�''@q�V�!&$<{�<M�9~�T�����8�$á$�I��5\>ԥ�.����eL�J���c����8�}��4�Dr�Ee�{�P$��R��y�?��/k9$i�9�~�-�2i�4�	��ň�3TD~��)Je��M$q��[���p�$F�5iR�b�/����g���44P��L�S�3�ӌ��ONϲ�a�z��ҏB)�a�ƹ��w�3�hr�cI|cu���=���OJf}�w !O#4=����+���p��p�#}�{�'�	��'�h6g\��d�w��,�P�Ys�tS��I�T��}�?����2��_A�5^�2`���#l��,�7�g�h:I8�`0#{�����m�p�S�9u�d�+k��+���kќd��֧Np	녘<a"��K�gv��	���)iѡ���&[&�N�Ř'g<f_�q�M�S�9�����>tw���ߎ��-F��%e�gΝU	�Ap��o��b��Zk��O_���1����%r�(�i�(Mڏ(m�4J�HU�R��UՏ~�_m�(j�))�j	y R��<j�+$`���ql���~�j�9�>�^l����Q��=��s�^{�5ǚs�1T!;� ��k3�^:��s�Zo���Aq۶�̔�����|P�T��=	��X!�a�/���87�G@��^�������}�#���#�?���9t�v��6��i��%%���5u�F`i�:��R� ��@.��������α��N��xN�#B=�Oz-�B��7�B���w���{����k=�����F9��ʟ�U<����ĊUS�R�ŗ�-��!Yavl�fnۿ������}�t�K,M�
�8=!�b�x?�.C@��A!YNٕ�܂RR��A�{��5ڰa=��/9�n ��އχ��� �dF�z��!��?p�By
e[���)���L�1e2�jl�o��P�k83h���'n���?��[�. ��k�T�ʝw~���~�ׯw�y6o5���磷����׽�e�����}�s��w��ڍ�n;u��:,�3��{���K�_��o/�_��&�o~ ����.��]w��R��nn6fQ�
8��7D�V�]�tG� �u����""&.��$#e&@��՟���k1��`E�9$4� @=
��5�G	�+�eBKQ�=�Z� -i'b��@��;YLr�/LLO�����.p4�A����n<�Њ�ra��d�SsEw(�%fn�.`@���	�2nX�Ȩ@�/\�R�:H+Jm���� ��&%[�;�IXhYF�
VmG��AJ��A���Ĝ}��RaN��!!+;j���Ea���!�&�:z��-8�Ib�|�� ���ŢÕ�H ��R�g���i�
h��k�#O>nN.-�Y{��y�I
�(R��ًKJ�I��7Ͼ�<��ˀQqA�%$̗43׾�}f�����)��1��bD@x��'�3�>o�H�J=��g�Ι��q�L��ѫ+�����1/���Y��������R��H��s	s�V�}��@����0�З��9�li�Z!�^�u�=r��߃K�<��*�����y��Lo�Gn��\���ļcϿz"���6U�P�_� �d����V޳:���� �\ ��បRB�\��|s����=��q�vnN:g`��]6߸�[B2C��U�v){Ŕ���MA�x&�Xo��{]rQ.�B�: T�?�#�Y�u+���"����\t����sT�)�-�l6 z}�?�`�mj����FpP�υjk^3&%Qb�U#�V	����9B'��έ[�-���;��Ǉ�0�j^���/N�4����%�iMLp#���&Wt��ܲ� �#B�,@ȫ�7N�4ӓm�� �� ��h�� �`ά�Z)"��C*s����4���⒉�g��5p"���kXι��frrΤ :��8;�t,�=_SsO_���?��?��ݿj@��������G�fa�mܰ�d��C7_��/~r��_�C�����������f����Bcjr����ܺ��w_y�]n���΍�����a��G�=���p�C������|��M���ߔ��h^#�!x %���H ��b�V��	^"' ˱�QYDB-=�qa��
�EֈA�Vs2\U����d@H9h/��ۣo/�m`��+(@��`0��'�XPy�b���x���3�v�
ΐ�
�s,h[����us��baW�c��D��3�9`;N�M��� ��`'�g��굀����"	G,} ��p"=�4���u;�,��&�~�@�>R��Ϩ�7*	T'�[t	N�V)3��J?�����#� �/-��O�l`k�,$E����s�v�`�4F��_��aFS�&��|�u�?�⸌֗Pc�T������rG����"Vo03�� ��Mٽ���+:�u�"-?���74�q�ff�����J3�t���BV��V��ɕ^+� �.h`��J���fnvƬ;k-���^?�k������!�]����z��^l��N�ڲ���r"����W�_�{� [N ���{�׽�z*�̀�ӌ���������U�]J1t����[d����w�A3@�^��:���
RF�G�C�hX=�.�a/w�X������P\	\�k?8![Ɍ���۴�.wLo�g~���0�����dL�&b�����:K-�P�Px]-�p]F@G):�](�����у�B뀳f��s��7�h��N���0�&�U���ys�w�cN..�e�d��"�.��O�t�%�����86Kfӆ�̇>����͘{�!3���i}�<�m�J[��H(M~Ԗ���]@Y@�P�v��C���N��H�D;�/6��4��ȎMk���?���^�s��JP��ѝ_��<����k�F۴}��uW��§n~��tܹ����G_YZ�����F����V �F�j����?�v����-����]�I�|�Г;�Av��c�.w�����ِڨ��陙�u�y3��^�Х�Zlq`1d�[g�U�Db������S����-i{�O{{�~������7@� ���p�W��x��u�6" e0�a�<� ΅�
-X�F%p�zn�1U��2���Tv��|ƮT/5�iZv��!8�	�E���Eo�Q'q	��H�K��A�*t��e�D�B5��wl��.�YA�&���X��ٖ�T nl�*qa-i^Wp2����q�j����'���Zc�ڳMv8Y�j1Jv�# (���H���Ҽ����+X�(kf	v��Y1���l-S�,L��ǀ��*8f�TPc��Ė�V�uNΥ��Uv���'���f���HK&C8�u���$	�P�#g5��j�A��&�F���i;��h�ˮK$DA��0gAPN�=@���%���;	�"��4|�/��}&!�+%�N�׶:���]c��E��)/+���CWyS�R�0� ��yyl~ޜ�i��u�`Am��e|>}�cI5����UB%Q�)蕠.l�P
�t���/��;K,�@	��fC
�H���0��/�
�J�;ΐ������������ob���2�"`��v��A�ss*8u���f�ٛ	f��9a���f{z�$H 6|�d���4Q��05�)��r���҈�9� ��n6����D��uS�1;�P��?q��!�0,�馩�Fn�&G-�=�0��+�}�y��6?�P���67�t�ym���֮?����Y��0w� ���߸�l�|6����d�n�i��桧~l�k�=v���C˞;t����v��&&��߼�o?sˍ���u��^ye��?����M���E��a��<պ��}��ɇ�^yZ��7t|��y���}�s�޺y��������i5�c��͇Ó�OZ� �P�7�����tVD5�_NMϙ��t�T�����g\�FK�� V[I��&��$m��I�dt%=�x�,�TJ���� љK�ӱ����������6�ա��?*�?L�H�xA$�3�vK�/�1��	æ��U�V\f���M�uK�Krb! ���r7���1������v\��'5X��A�Cg�L^
��H��}��M��K0a��P���)
�<>jz�
Q ����&=��b!(�w�(��V!�>���&u �I&CQ�c���&
� �A4d��'kl�^ VI�h��D�  �IDAT�&�ꇓ���sL�#��ʝ*��9u�b�,�_u����c|ж���<w�B��7�;�F��1�Վ��� ���}��� �`y�����+[UЪʆa�J>A���Pg��լ��q.p�B��-�IP�S�i� �{"���C�^�
�Q5��q`7K9յs�A_<0 ��=�����9�	�;�3Q���9jga�}�r�!5-�+l��6:���m��+�
!8Xt�6H�w`���y#�xF`�����w �9fgX0�� p ��D�\0`��qC@�gBa�sA�DHr���;v�(C�{p/�̆�:'f�֘���F �^O�KO٥��@����·�y�ey�.�B�$Q�;t	�40Ruò;B5^�8!D\4���K s/� �\�lh��;��� d�q��g��q�(��� al��MS	�$�����?Ef-1h/x����v����e[^���K�� �nM����	�S����X�.qs�-�;t��c�b>O���{ʘ��'�x���}�s�{_��~n��x��u�,�8qb����}w?z�/�z���5�n��&Y�޳����{��w��OO��_���=��m��n���ě56���=��#g�sv�\a}Dm�cd3�����0S4#�'��ћ����B@��/�I��Z'���.�*��R ��d���\�B�R�{��$Si���i�G�P }�4cؽ� ��h�tc�=���v�B�e*@�B�m��j�����`e<�u/�m�ާ�j��;�9� jm����*%W�(ִm�UP�u����r��H�9
f�:`�`��h�1��34k�gVL�����P~ER�#�=�wU���u�/l[T�Ӡ�� ����l�Y5Ǫ�\=�0�4؞#��e�$���aw���:#��*����S�}�yDv�D�N�C�RȀ��A���?+Q
+�}8)¬|��Ȝ�B���`�����;v�4�}Bv+�q����%�=V��C�~��W/�`�����<BF,�C�3����\5	��v pW��\@����n�YE&�i0J{�V@>5�U�|"$�Gٍ�~(a0ݯV����B:-V�L�?��OKbt=,A�h�)h���վ�ԉ1��|5�Jm=�I�x���)o"�Z��Łc	WSלp݂PVu�ʵ��|��^]�/}�+s������s��4-Y`#�n�g�5�Մ&E���Y�d�1!=FM���tش�O/<o�w�����_r�綟A}6�~~l�=?��?z����Թ |���Қ��{/��/>}��3���1��z晹��������X��ά�PoO��Z\O�"�i���|���TC��
��|�]�gQ���g��|�{[�Rr�`�L�w9�9�&�٨� ��������Q��(�����<wy��-U�x�(z��`�e%�,�@���905;�sqB~�A�L����ʝ"��!��I�^۪��`�VG ��a(�yx/HφE��4�]����(���]3�\ �{�.���u��<��>S����F�$���P�80�k�s$f���[�1��0><�+Z��@0*t���j��G����Uo:ί0 �����W�^��꠫c�&����M����\���ъ�rI%�З.�� ����̔,U�0�W=k]V���0�F?��uת�L�d���J�T>�aV�X��@J*��p�"\�PrA;�-�Ȋ���'8OP��@��ɠ�@�\�Q��yK�E�5q,,�{A���$�#��[1O��"j�\�������h��
���A�+z$�I�S�
�̛?��p;��*��+���Lڽ��>�f�%k� �_J,�>�I Ae`\ug���ѿ<Ax	�i)}��W8����o�a�{ϡ�Q�}�k5C�Z�	(��]��^�N��*P.{��L��_P��p�Ko���-�#�3z�I�����-t~�To�v������E���L9N��29=$ug�Aoã�����_��+.{ס��w�"5fy��ɗ�Y腗/=���W��;wnG��q�Y�״Z�]�}�?�x���ܷ{w������[������K/=3����'N�x���w>�QnҸH�M�9뢼�>�Ӽ泬��lP���Z�y���g�F�:D�3b�:�I(�P�Ҙz��<�(_xǈjrdn��Ȣ$+j�<�1�kHwQ-v��ŵ������"�Y8C0������(
O&;Є�	6�5����ρ48k��C���yd�� i�����}����y'7: ��V)�F�Dl���e�/��³$�ɂbڰ6͆j�̻��B��B�\�� �MJ��򦳅��b������9��Ta�΅�]�Ej.�#�DC�#���8���d�����wv�65��#c3n�(��כ���]�N;.� �p�-�ȅ�v+AN��縍 /�'/�_��N!���E�N��5�k$$��Ӑ�ňI@b��B��P9��$+	�o1k�P�������� F��6�.��2n�S8Z>��	x��"������@I$�;�U� L��;ĜS�h�D�� 0�Q��`2Z���V�8IqTmEsqK��~�e`�|��W/�!���.�U`������ #��Q鮚(WO�څ��U��vi����5O�{佡@�����c� �H�b��+�pr��'sz��#��_���;pXF�Bex��$n�+�(�������"#!BK����J2��~��j2���C�$|���rY���o ��X�N�{X�W0T�A�de���J�8O:[VTY(�FH�g�YS^���ę��o�ˋ&���5��m�tp�֭�l��}���5�{��G��~��׏�ʜ;��j�;�Jx�d���ɉ;n�����W9S0_}����~��Ԟ}�D��a7ǶD��"��~S�<z�w&N�ܩ�_����F�m�c��pࢨo��\��6]3F6v{��qiY4����i�N�܉~/��n4�	�M����#��=ٮ�"�"��כ��]��H
Dq���V�,�m�?g[��B��ٌWvh�\XvE�9��%���4�K2�Z��/NAб6����(b_ą����!��CL�?"<���%&5.�6�g�;�3���tX[3跔� �9�x%)^��@_���s��rNi�
��/��mDuȯ�V���|��i�D)9C!�a���\��1`�����2�E�I���Ys�g�T��BT)�321|8��#E��P8J��� s B�"FQ��՜z����!t��kFظ1lay�i{�Y.�mx��9T���b,X��D4�0lE�ͣq �0".���DF�ko��z)�h�ȑ� ��)�=�'�������@�� ���aQ���c���K�$�Y�QdAܑ��Z�>'�b��?ɽ	,����B�ZhvֹB@������P��𜧀kr���	#��/��
,A�\9��a�)2�N1��Ȥ!�r��������$Չl9F����� o�Th�3&n�<d�9�p��o�=��J��>�QrE� �� �r�gR¢ˌ�X0HhB�g�f����ןk�s�Drm��F�Ϲ�� �@J&N3"�#��R�!�,�8~�ș�0TA�%�&b����b�����y��QV܃���n��c@ԩ2�z��n���My����J@�r�J�����t �2�e4����ȵ$@cjΏ�$�C/��$p= Jc�8��&�O��ugNN6�4Mk�^w��k'����� FIrzr"1y���m[�}���_��[o}q��������}��������!o�i��y:���'ȟ��o���j�>���Es�����U�$��o����o�Y�`�$��"���.b�۳�N0b� !�\�V�L�� A��U���}�4���I�>�,���Ȋ���(�`���8��(q6uI�Z
v�rʟ	S([���0 �Y��aG��`C#f�a��E�s�9[�qE����S��6Ϣ��8w���l?G���<*��ߋZ�)��]\7��=��ȭMS���yƻa��
[ �g= ����H�v9"�f���kL��O�M���3�Cf,�h�K �rx���|́�9 _��ki;�q�ω0o�&����5^�h̙��pP����I� �~s'zdT���A�Y�<��涰��,��(xip��|v�0�Tc���=�@� 2$�P��e@:�C�L�mpM����HEB~_K�B�\M&'K ���t"ɜ�鬘T��h�+HGFS�b�5�%�T�� R�X���̽������m¯
�Ho���p0®`����6b�q���+ؖ�_��5�8��̋E p�c��s�@�"_�>���j&Q�Tf� r>�-w�8��f�YK����ljj��n5N��Ooۼ��}���O��{Fg��t慶�;��G`<�����* (�t��"��1�u�� B�Ѽ��@�l������Ѽ�)���C��. sd-�������.����s��hPG��L&q�Zzt0%h:�q��$��lv�,� ��#�j��\�Km�"���,r �|�'
��8���ˬ˜�v:��3B�Y~�d�2X�Ke�zG?'��QA,�%mT�mASf�md�l�dm�A����s��EĚ�wQ�fS��k�Ǒ/ QY�D~��x0L�
L���E���XW>�!H���*B�9
���) o����˛�!X)21�޺�pqL�rS� �R�ԲZ�L��XX�ۢ��H���;��(#���|fo0���Țy_�ٮO O�dH��n���E�V���5wn;��}�굽[��Ʉ�L7�x��kY��_2���G��7JV��ug�X��1�M�9c��3X �C�h���e��H@T���^�w�+bT��# �@e�����x0RYr�`� �wE
� :�,�e���{��wiV��u
�[{~�>��d����Ҩ7�$��h�xhӡ�q���f��8����(�C���xT"���.ק�ut��E���s������}wΤ��V�h��~�����#0���G�8�����S��x�#0�������h<���xށ#0����>>���G`<�x���8��������#0���G�8�����S��x�#0���������Z�    IEND�B`�PK   繆X�=z� C� /   images/9595c21f-5942-45df-b2b2-1a139a6dc1aa.png��Sp%�{b�c�c�fǶm�c�IǶ�t�c۶u���TM��<�î�j�~�/��ZQJ
RH�x�   间�
  ~ ���B���JF��8'imW  ���7`�t�� ���/q5Ϝ��_���Y��|��;N�G_��ȩ��)��Njhw��(�H(t]�~��v���OX���`�������<�rX<��#���;�x>v_�]w�"/.�%S̸3|nw�>�^��//:;���w|-�i��o]��M�N |H�ƶJT��u��?��ʽ?;�>����\_׫7=�m��GI&Ϸf�����r���N��|}z��(~g��-�n�㏽��+���zD��!a�LY��Y\�ۏ�Xm�~{��R�3���X�Տ�'͊W���g�>.I��uv�~��Ƴ��˳����kC�����S�#(rs!�T*@'u�Zd2o��Û�x�}�bҚ��>
7�y�W��؞�O0���y4W��������ꄸ���f�މ?P�/��<>n^0*�D�h���?�
�Vmi^v.�H��G�9����P�vK���ˢ9���A��I�r7�iӞ�^�9h��ѷ�Q�$����e�s��{���}��:�L��ʓ��9���kA|�gN��������u�x�k}ӛ��G.񥩘rJ�o��TEH��*˗�R���b�$�˥Ow�*�`������o�ɡ���/�ީ���K��I�B';20sF&;l�eV7W?͘M��Ca�&��(�96a�s�t�t|x�	`:e;nF��� ;���N����x!���Ng��a���Y�#�z���F�+Φ��+O|O$H��?x�Vr���)]7+E�:�5�.���9� T8>�'H3Vv���.kL>`K^�5�*������r���mh$�Խ؁��iv��3�w�Y�}	�s�2��\���o#w?��Ͷ�"�Zr{�
��b�[5�t*�f����̊�wz��3��z��x��Q� ��J�yI��z�N��.z����tm(c<|?��H�t�M�!;�ޑ\x18�N�-��tM`�8uG��j[&���!�/}J�
Ѡ�O5�^�v�y�a8
3HSm���|k�(nSY��>'[��]�1�<f�^��ٞ�9m���hl�8��tI2w�|�Ԯ�g�:=��i�a-�Φ~]J�u!���M�S�2��&1��p�鳚dK�4UM�mZ.n��i�����lP]��������Ӗ�Uh�4
x
(��i����HE���{�[����)ݤs?�E��u�~k{%��#�wG=��2�mt����>�Ŋ	���y�	�]�1Б�b�z�D�<���&�択�s88�¹���|+�ݥ��^�1�hS}s��f뗱{¿"�� �ՠ����"��rD����u1�l�e�c�1�����` ���}����O�>�?+l��x}���|�|xX���˫{B�Pڊn8�n�l�9��������Mo������e�Xq���+&��'I�q�:D��C�@�hw��j��<���� ������NQ�{�1Nc`�S�R�v�l��kU�T���*���E�j'��`�;d�����0̵�Ky������Y� �c���k� ,�1�&,�G|��y����t���u~Zh�m�y{�����w�̌�<1�Mqˊ��A�L�`��c�Jsu��j�����{���A��r�ƕ��2��J��!��{2i���	L�ʰ�S|�ic��P��@�T�Q�� yO]�o����:7���������y���E2�>��܍/�
zϛ��Ӱ�YH*h]�g6m����1���$������^c�]�������n0����J( ��:�Vz�Sޫ��T�"���1��YȤoa�I�G�=ce�#ڊܮ�W�{
�qM_��["����qt��W�C3Zx$*ًփ��^j��c�٣�aZ��!�!����U�g�Y�?���ĥĚ-��r�3�(�� ��ħ��+s�fyՊ� ���9�l�P���Jz����+c�8���5�o��慚?i%@�K�j�7��4�y�	+�Q�Q�U����Y�~0���+x�D�=��h��3Ȼ��*u��@�]�Bz�6�C��ŭ�@#st� ��������>��$ܪ��e�s>�k��>��1O~%a-Y]5.�LD�Xτ�����]�I2��81C�e�H;�>�B.+�_��n�T�Ίp�6.��{u����{ ����7�n)q�����	�o�mO���	���ʏd�fU{���j\���ǸRq>U-�M����{D���0콂`�K$w���f��:�sˍ�4)8A��Xg?QvN���iN�T��t�=C����Kѻ���sg;�u�����_��E��.����~��Gc�C�Q{�R���O�T%��J-F�G���a*����eJS��f�)͛H$��8ߣx;��t̓��:2*;��(q�1_Y Wp�� ]����"6݋�e��=�3t;^�����p���نVb*�E7
7|�#U$z�g&�"��uɐ��%��(w�w�[�4O���~[���+Ψ��[����O�;aʔk�Xb�e������!�������ۊ
�d�����G׾b.�K�U�ԥhfo����9�y�G� b<��TMޝD#�Yɋ��W��	�2�i�$1J!�w�c�d��a�A�.>U�C�-T��� ?܅���\V�ʑ���;�*b�Pҫդ�OnU�Ji��\G�u�]���@oC�b�ʿ����}V]�Yv�I������2��oT�;M�3��\����������f/ٸ�d�2�z����V�2Uy���cdo,�}����?ڔ�:o��;g�qOc����>w�Թ&a��T3f�C�R?y�L��������㼟��e[�b�N�P�.}[��yW������1�f ��(�޽!-�7�eW�,�fSv�
�EsH����j�@F�N(�^nP�K�Q���َ] ���Aݠp�9�<*���}'E7HFF�����OGXй��I=&2��P&�B�LHW��\��>�5�LD����cQYͩRi���_D��� ם5Մ��8��F�ض �==�L�a���F2U��	ŏ�.�l�9^¹�
��T�.w�u�N��#.��ܧ:4T�v�6C��nŮ�Z]q�bl��D&�
6�O��8��=��Ӂ��S_Ε�}��i�6AfO��{!�e�C~�gY��}ݤO71���w���|~]߁r�ֵ��P����v�r����x���{��Y�����xK(�P���o|�݈�A�g͖�5ʌԔ��
"F�[{#j?J��c�ȡ����g:,�i���1�eRŋ�$�(���*���f�C�����v���UI)��
	
�e�ʧ�Zk}����2>���n��EK�S�����M����
�� ��tf賁+�я\jl�L��@����,�_8Q7�/����$N�0�Q*�g1���,�Hl0c3np[��AY	��/�ֆ��D5���[�1\I�W$�ݛ�1o:G�(d+��)k
�m��T�ýW�Ep=��mT%��C$nI>�=b�g�;���`������-����=�=�
ͩP��d���P�2�^���bw*����]~��_[|=3�ktiI���L��I�ْ�oQc"Ġy��E{!AMh�v��a��7Ȝr��)�
:wڦŖf����Е����+T��Џb�4>0�%K��ԟ�-J��j�����2G�Pz뒣��w���:��dI,rwu�Zj���}_��cđ
\,���_�X�*"j���AIJ��(�Q��K�:���8Zj�ӨSQ���Op��ct����7�.SDc6�Fj�c�ҿ{���
��CΡ|Bu�a��"�;m�zT�3��Ă�9�?[2��	YgIY��H����q�ҖȷU`�bx�	����2���(�,�xN1W��NB���v��<�����c{�cמ�jބ�����m�� | l�Q�Zv�qe3c�̊L�'Q()-�V٢R�<�BdvG^-�*��Io�B��%l?�NfF�"[�UL9������Ա0?|q����p��%N�;����.ۮ�;��R�a�Ji�xǍN]|��s���r����g�HC9I���擦��V�K����.-��D&�3�w'0@[rJ���b�p�Z�;���y#CV�+:,}ӱrxo*�P��D`�/���p[����D�X�':w�;�����t�)�6&�@�.����sz ��Q����e�0�ޓ,�Iq�u�}��}�KY�(mO�ր��L�����*�`�W⟞c�;ߏ�����o����epɌ���������RA�Щ�Wbq�t��8I�k��
�(W�WR �㟍��&�U�W��y�N5�[Ɛn*�W9ܟ�&�_���=AӶ�1*$�(�ZzX�k�Y�+�ɠ�|�ǀ�р�\���������u_����`��m��mꒆ7W���y$�"=�}֥\gv!��E ���/��`��fZ�U�*zu'�����Rmz�#�;�HZ��Q�Cb��`u������������&����	��%�����Kr>�7VF�߄��b�0��L� � &$ψ��Xn����?1~��:L郑竦�C�����gN�.���������������	@� �`��������M�Ӳh7S��j��G���B�r�����m�[�l1&�Xu�Pō:^E�{�Z�d���N���ΟkpAj�<C�c�@z�ɷ�Ͷ~�����XI.s�>  bR3'���	������������&r��3N}/�����@c���y}�Cσc����'�s�f� /GZ<$\U���RM�V_(17���ĢS��q����^JH�� �����^}�=$�$�;�Ar�7�O4���y�Ȃ�{хѦ+6���k�0+��U��[�T�X�������aă�
dyRm��b���8,�|�9]S�
�`�<��@2�y�ڥ�4yd�һ�MZ�I(�s�'{'�c�n�����(ۗx[� �����6M3��⋦�򯻗�3�|k����S���ҍ@�I�Gd���w|m���5�Eӑ���b��\.�S$*3�g�%/#[d?����T9�#<	���HȠ�O1�?�~MK���r`�J�IҢpT�ۧ �B����rI�-
��1�nLO�dQ�=��� �3^���Z�w����;����_U;���Py ��i���{F�tm��~��\�J�0�������L��"�hO�c�#������)�seX��cA�F�q�kj(�!�y��0c�?f�vlu<^��j8���R������jn�$Ja�h^P��(:��.��A�ҏAA�1�8&�q���"�"�P��e�\8hJ���c�U����'�H��X�ϊpP�ͦxH��
�g�Ź�:F�z�;okz	7�o�cE�J6-?]��h�����4mkS��k7���tץ�}%,����PR�>�Y�0yٲ��FT.L_����v鵤�,E��cCeҶU���4�nm��ep�:�E�{i-��h-֌(~�A֪�
Aګ������4���Z/X�i��˹�Ӟ�Q@���
�͑�5K��6/����?��h ����t�zlܘ�/q��e]ɱ�Ki�Nig���+�9n�pA���/��ݺ�^�$'�Ib��s.���t�%mv�غ�$92�p�J��|y8WJs/���ش��������L�e��SU�^���o#ƥwg&�K�����ASD�J�ڞ���e	*�V2�n�"�d������}�fo0�����i��`"�6�'�8Rw�����/O��|���|n�z��g���UH�\-5w|�Jn�aW�����p��!���v
�ɒP�^_낟�� �J���Py$cǾ"P$�7�/�sC9፯�H6jy`4J��$�PK�R��k����Y����W�s�v��=�Ͳ����҇��L����g掚AWk�'�O�7�&��|�t�ˇט��G*��=l�Y����CxE���Ѵ�����A�`��E��׮u����b��0"���/��:g�6��5Ju���6j�;=3��cA��B�^�~!��� ����Wَ�v%S���i{�tU�Jg6\��<�0��h�wdN��>]Ti�W�eT�s-�m�Ĉ�ɯ���fˈ�[c]˵%����3ak���9P..�O��������si��[�0^�f�G�L�lxp<0]j�摒A�J���db�\q,44��2-��O6ڦ3�j���X�ǿj_I�JW�q+��R3��x���u��C��%B6(~fk|P�7r2�Q�U{�XZ
������k�܉X�ɠ����+�	)�Q���ֻen'k�e�LF<�I��ή��(��L�6wHGM����	X��uvˢ�
��3
P���QB4mA_�'���c� )���e@	�ދ����M	Oai
vA�jp��J��jo��97fIY!2�N2�k}4�|�؆�̟���{�[B��K���t��ݱ��N5���K���#Z�����6��)�:.���i������瑺:P�ľY�G�皕2����@��.U�%�9��	IJ�Y�\4M��H����J#k�
��%XG*�)����(ڻ@
�)B�d�2L�\�L
F��M��!c_�$���H�s,�x��G��N�"Z3�x�#_ːr(���R����w�?�����d_|W�K��Dζn�Jeļ�tZ��GG���?蝗�����y��0��k��	������*�|�c��c��"_�Pb�@lX��)���}��΄���]����ɤ6������@����|���v*	k�-�>��&}$���I�ض>�{�e�!K����X7�m_;�8����1�/�٪��9޹�e�1+�G.R���B����'w�,��M	c\x�~��R
#��EJCQrJW��P�C��<�U���OR��՟b.�7TgN���#pa��c�9�xz��<O��s�y��~���̭A��)қ!;{�9tt;�P/��e�L��@�Ŵ��)
7WA�EU�? %O�Ո
}U[��w�'j�)����t�};�=|�EW�p�͈�Ȼ�>R�>�y��ȴ�<_�TO�C�&�'�{�l���$vsu����� >�?�$j���G�o�5%��=�
>�b��2����%��"l�,ӏ��{8nA�s=S@�J��wi�3�ҋ
�}(�H�.m��M���h>�)f�3��%�ZS|��x2��ę"!J|at�Lx� {�sN��~���C�Z��%�v/y������xְ�;r�ԏ̪hn�ϙA A�0{	;�U�"�A	�ܶ�&4����~ Zl/>�&1Xe1���1��VcV��uǡ�Z�n=/���Il�>��H/��Q���߶��ʆ�o��b�qً��Cѯ� T�cO�"��W�|����/���M���E��1��)3^�s��Q6�X+��'�]o��SB�)�0"S2jwز�L�G��5�sW?����-��xոѸmۅKK�NhJiũX6tx���^�"\|�F�a$��'<s��vƬ]�7���'�f&i5#Ǉ��,�����\�y~�LU��'��*jes���=�#�����v$2	!)^��ׯ��#�x1���c��z����+�;h����}��d�#sTc�J�:?J܋ߥ�g���:TF?�Q
����a�q/�5�*`�h�񃃣�pV�Ж=d-�����t���u�3l�D:l��k�M<�93Y|m�PGTeX���ʏɚ�-\)�mt�"~-/�R>��j^��aDqo��0C�: E�w�L���;���&�w��{ے����������r�L�p�as��a���FG�A���45a�VA��'��0ZQ^J�2<g�=��d��9?IK�V�|�( \�0��>����!J"���xY��x����\�c��
�M>�='�&�Dx]!�g�b)���O��3�U�{���Hn�����^7rٶ�N nF]��*���h���]7}hʝ� ��d�j��E�f��JIZ��'��\�U��Q|c!>?�4lEu��èǲ�4���:��g��d���y�Ͽ������mM������Ro�Mʡ�@�LʧpyL@�D�KFdVq�XT*�� GIS�q�(��$-bjb����w�b�]72�Px�N!�S�&�L���X�ῑ����D#��cL��ʞ��<&�f�r��簙�"Tl�	x-&��f���e�VlˁK�}�I�!	�G��<up�����>�����1]xr��g�i��
��얕�j�&˅
+��?9dYHZʣq�㱕��iF'm���M;�v����V�"�_6�~�ko}{~r�1|묂t)Sܕx�� �a�� %��Ǡڜ:0�T�}(/�j�	.t!>Tx1�?�(p�ϑ3H�d���񛧨s�xd���*�b�I�!�Jy���|�M��`��V���weL@��-�.�{��&� "c�b�L		��9�u����ӃQ7�;������MXL&G�΃�����s���uw��+t]� �۫ԙ��4�m�v�:V���B6�i������Bk�)Pq�p�mᨦ��@�^K��p���;�QJ���m'֝h��F���M򆘅O�R�T�?n�H���սh�__�H�'���*^�N#OY*��eg���c�$��%R/�o�,��$�$�\3�u����njkf����#ȇ��=�9l"a.�*��"�*����r����4�~p7�����Z'�b�J��0���Y��Q�0�y;~u&���XNۏZx�-#�6V!n�x��N΋�j�,�؎)U�)��Ю\v|�ܡ��eQ�xh�e��7\�Qo�g�����2�C#�@6�o�@KyG��e0�8ǧJ_ ��+�:�x�B���5��u0N�xx:�o˚�w�G�n��9��a��I;��w �**����F��������x91ģIȥ����$ǁM��VAz
l��ZG3�:��T��.x*��++��M�
$��}�Њ���BFXN�Oa��b?�DSH�HF�Dfs�'[��� ���v�%�fSe8���e�������$���WJ��\�<��g9@-
2�Q����^=�����m.�?���d�|b��rm�oJu'�W2s$� �޶'�NA,�?c��L�IX��i�=�~��~o���!��W��ؓ\>�vB-k��:||^���.���pU�bI
�:J.������su�X�!�uM��վtO�l���>C�o:ﶃd ^�$�.i �0��14�g��El���\���c�f�24�-;������[�Ϲ���ӭ]��ж�'g�R|�s�7���6V�@#g�N�ɴ����`JۃڹtRM��LIN����z�v#�C�������XDm�䏛L�X�zԛ���G�هW���\Ց���"�H`m;-.���^]��d�׶�i����n*׎���߭g��>�f�����gG�-�֯
��zc�x�&��ɚqe;9C�)�Ћ�x���s`��np�0^�Os�jp��n��H���e�=m�fw�D�Z�ŗ,�y%�M8�O���"y��#��ú�>c84t����s�+�C�,n� ���N�����CǷn1�z��Y�����h_�Q�I���0k���I���Fd��j�Z9촃?.J�cZH����;��Ʊ%ǁ[p�i�4,����G***���ݯ/A�OG�l������H�0��A�S�����jjn4v�R�9�<H����rMGF�e��7��3��:h�v{�t9���w���ƨw��/Ϻ�+�ު`ަ�'��~�d�np�\V��	��X_�m!¢5�<N�$ij"v���C%a=*��$J�6/��}ˋ�z��G7^"�v�(���u�~oji��:�,w��"ރM�+d\ʀ����:�F�D����;�W= "�|���+Q��i��3X<I3܂���ȢC�H�/�]8k�k�鑌�8Ğ��Bbg�T���ث&��B���/T,ܮ��1����D��}M������o;~L-�T �+���������>����sgiغ�+��F]��2��۰�A)�Wg�N���,�bqM*6o\ԣ>�C+��T�~c�M�V��i�S�~w6���?�L�
��՗��7��c*��z,ޠ�E~�9��x 6O� ��3�AˇI�W	ϹH&R��8���������E��ׁ�e4�����هL�(��sd�r��@���tZ�Lrψ�?��>8�����Z�>�0d]�Q�_��eA�$�emjc��AǤPHCѝɨj��Ƨ+y�����j.ݟZ��SZ?G��6I�aQi�a�� `�#�V{���8s�l�0�"��Sj'���v��U��_�Oy5�v4��i�{����"4��s
R8>}�$���Op��O���-\��@�[�?�~n���q�qG0�Q�%i& ����z���leMs�oʿ�M3���޺�hX�� ��}���!
��;�sc>̈́a�WO>�ȵ\��Ǫ-Y��A�4��tGN����^O"���<���<���z}����w�|2�YԲ�̿�"^E� ��k��v�UF�n�(����ܷ���I�/��(׫]Yڀ;�������8x�)�D��b>n�3�~Ʉ�`�!-Ar13�g\��A�����K��t .B�H%�sV�'��(e��qAk*���l,�T��/�OG�M#hE�@�.�b&�R[b��#�D��ð��s�y	�)�o������y�2:L|{��r+�O���U�1�_6u�G��V�����[3���7%L�@'W����@ L� F�'c�$�����]G�������T�e<DY+l���#�����G$�Y]��y��4�4RHLD�I�&��`��G��rbV2w��XN��H%;�3T����B�'qm��B0)�WF�2��ꃚ6�1���L")_��hŝ�(2A�h-�j��U���s�rY��>���s��}����SWQ���X�Pq
)������C��p��H!�L�#E�ԏ��W+�}�ݿ�2�`ޭvvK]Vib���qds�#�CaZs���t�99o�`|W���~-%V�=�)8ؙ( ����\��r��1� q��b 2vO�@�9��)ۿ	�qF�n4�i�d麗�H�o��;,�_�b�����;*��M���.ޅi�+Ƽ���}x�cَ�f�Tӓ�SO�j���Ԃ�,���Yqo�?�gO74͡!�_���^6kL�g��*��T�`�=��,Lc��]�J�E�Ϣ)`�tca&P�4��BB�Ly���TY��M;)����ڃ(�P:c��hg�za�k�@)<M7D�,,�� �U����ˀ���3���ȍ<�~���y�b�]E����r~��^���A�ޟ�;�Yz�9N��pA���!F�����Ql}c+���v�~�^E��up0��g�K_J�<�@��)�b�O��%�K�&:�e_���e�������íI4�E#1_B1��Y2��J%�?� �[�H�D
�P �Q�˧�z0EPt��>3/u�-b�?�>���{VI�RL��A^6KDS?sSO�����	m������G:�?���6$��Ԟ�/�~��#�c?��$g�-1"_��|���(,�vbp�?Ir�1o/�8���x��)L33؉IwwJ�d*`<��جʑ�����*C2�G##iF>2�H8]���6��]�]�/7ۉ��d�TLGrqwU9�IRzиE���.eM���R������<	����iVn�=#�vɩ���L�T�>�!ϑ!�8!���٩�>2l��/l�����nϯh�i��v�����)5N�h��Ί
&�t0�s n�n���hًTI�fq-��w��"�ȱ�h��9���IU/����#�]�'׍���${�3X� >����ؐT��m}e�����k����J6m�N:�R�S��iV�ב=��)���f�p���ƿm	����PE��+��-#Sxv� �
)JV���d;��2D�['Rx{TS�H_��~j[C����Zlu�o�#'���|m[�> �B�v�'$�
^JLp�jDz����)16�Ƃ����
i��y٤qTݛZo�Mo*�wM��*���q�>�V��3@���F8?��5�=����e��C���8A0鰘����±�ɞ�Wм�H�C�T'��[%�[�r3iz4D�x�Փ�0Զ����zl|�3�$ޥ�]��]�/}6��kMmȗ�|:X90e�׀P�{.�D�=�ܻ��2"ms)*y<rϳΓ)��WLR̆�%õTD/��h7'D������O�'�o޹�c��Zs� b�]��\|����Z|&�וGɦ<:�.���Q� �m���R�K�v�b9/�?���{�}C����m|H���������V&n)	��魯b�aÇ���Go�����^`��]hi��;�i?l�ܔ�Cy��#쏝�}y�.��i��1��߇�}�4���=8g�<�X�,�| hH�ϙ�d���C�W]�	5�E�^1�����E1���a5ɧ��ҕ7j1�dqhUd�лb��(�;�"�mYR�@ç.U�p􋋏v7�X+*��g1^I��>��rf\��#�|)�ĺ[+�n_���cS��@���gj'z�7I�ffL��&n�ϳ�q�͂+Kr���]I�k	>��\��6*���Y_�H�/Ѹ{W���>�b��QN�;����K}"���a�GΞ	ƃ��7#=�ę:�y-T.�A�1� �5(.��x�TT�{�_�����§6\1����?مn�O�x,>0�ӂ�r9`O�G�\t~4�H�2k��P
?&p� M�v�ӲIC?Wܵ�������u���c
�=}`�9f���Z�3��l���H 2��h�r)�YY�VM��PE0�"�,k��	ׁ�b�K
{�wkU��I|��2H��DUK9"���T6E;T�2�ݺ�1�L�x$?�2;e�+�j������^�I��V����i3�х��5k�_>��F?b9�|;PM'�]�옼��}őT&@ �����:b��B� ��Npr��c��^5�y����Zk|x0�i���O��������t�-z6 
j�u�cT�T�Ի|,GxOsUN�0�Otu&XN����7<����{{*�>�l�6�����{^*'@-`O���DuLL�b?l��F�-�	�V
�h�҄�џ1�iцJ0�5ͤ&VH�� ��[� _2��8ź�:j�3�r�X�.8��[�:>PSp�+��33Jև��ȤiGaW�C���ҽ@X��w��tGC�a���A^�9�b7��b��[=�k_	�#S��Z���Şw!��h;T��XЉQ�`���~S\�6�cQ�����K����<�:�IE�)�w��ģ}��D��宵MLPZ����t3}��ٟ������ԗ.&�
��.ŗ�3�1����=��	9d�ˤyk�|Q�b��CU޸62�O����sZ��6�E\v�j�\c��=��W<:���\�o���P��� �º��_���wuG�+����Lz}O�ġ��B�{x~��"㬄����Y��q����>����3����\h�D��ۤ��Ц�G�eER��з��C�\,�It~�oz<PI ��x��.c^=�2�Y����eX�"�_�(L�q�!�
�k�%Ѝ'�b�#=�q� ����Q.7*b�т�@�
�B�oT��#Hb�.}�������f4iM�����۶kz�3���	yژ�b�{yl,�	m9T$a6�8��r^�d9�g�`����p<��dtn.���5�8��آcQ2Ǔ�#�ĥL�oM��1χ��;N7�_,�\���m��-wV�,_��A PJ����X�s�׿�f�����i���)�.�cd8����	�t~TNRX���'}��_#�p�J�d��%DՃ�D�Z�dt����U�!�{m�dJ�A��_��m2�֫����R��EM�T��-4�c���ܭ����j�p\K,Hi���-����2����N��u��͙A�3�9��������C���7\��N.��HтV��5�f�;��w�h�I��#{[sp<F�y)�p6-�NIE̟��֎�G<uh�[E���|�<b^D4"��ק���mg껛]�q�����l���0*v�5�P��C"mU�ٕ���\�h��F�"I2�Z@��,��R�s8�Ƴ>���{F��R�P��R�>9�@F�A��W,&�Co���ch�,@�S��K�G�to*)�����S�jI�3�M#��N���}9ܠ�)`�p�G���̥��r;���\�P�N� aR�]��)hi�n�E������p�jn�҈�Q'�J�(!�$�P�\��vZ�i����� �����[���gT�!<�ο��'�r�& ��D}���Y��/Hک#�-K�<�������ֶ�%� 1ι�����D{�"7s��H�F$�mC���G3ݐ��*�?�.�$��j��3���"V��������G�J�~H�)K�\��	C|Og���n�����;�'y"�5A�_�_J��q�7����/y�h����!��mS�����y6n����8o&�+����XDW��-Q�5�r�8�O��޻����>b��T$��y��kѕw��T��wo��_7�bSlPxV��N�v*4��Snĉvz|��Y���o�wv�8��^���=����}2p�@nyB�=�|ߡ�E-��^��]�9�
xM�R�������Fs�V ����������x�W�5�֛�����s|N�"P<c��O�1�(�)����IO#N8�"����i �"�˸ �{��v�R��PL������םHs��>G��*���"�Xy�0�V������S[V�)�����l��@<-1���Z&!�F�F����?Τ�k����$��d���t�l�#0��d��������7���e�fC�6�k�[�N�M��� �I#�Յ�}rG&����+$́���L��uŻR�M߳�����VT��Jim\�&u���~���9����)o*1�Zy��[�%)
~e<���߽5��:�\�l�R(��7:��T> �v\����
Z(�]9l�8��'��T��w`@��o҂ `�Gu�g���~�Ȼ�\�lNVu/�'\(��bR�r9$�<���lU/0�X=J�M��q }�ZF�j���P��Iנ�=����qw5c���Z��G�x�����٦�D���Z�~Ʈ쫝"��,�L�A�t#h:�����1�-���%�se��R�ۼT�Vdea?o�=��?����6l���̃�u�}F�������6��b&�������h�/1eV{*L��� u��6s1(F;��-w����%��CR
Ro|���JV��_[3�M�sC���L��k�'�X+6W&��.��Ԩ���=�ZW(f?cߞ��]�2-�(��27b9�YX���vR�7�[���%ۘ-,\O>)�"�ǘq�Ih<ű:JL��d�c�%h�ZB��E�y�;T��H���8u66�;���TQ�(�E������W�Rָ��ES-%Zc]�n�������*>��xl������n+n��D��T�'S{��z���ٹZUQ>�"��Ê��_�|RW�����[�]�z�ޣ$.�	�n��TW�gE����4��T��*p��i�`��SsG��(:@��_�1�����l��r&*fW0ș^�h��Xk���ai��֦�ei9�(NF2����=1\	zA��I�)�n�&�����������PiEJ;^���O��9u����
킝�8���Vhw����9E�s&�ȫ�zA�٫a�9��d���d"�H�J\Y)���g��ej{"~�{��{'�x��c�wl:&^T�S�,rwp�^�xVpU@l૗>i�Lf�Ѯ�e������B���������Xl�ԥ�+���,p�����`U�c�~�Y�f@':P���������o�=��GJQ�yFDZΉ��r"�L;�UO+N^}�5(���y��a������v���i��R\̝�y�w���(����OI��Xݭ*C�T��ݻ�;�RԿH8�I�8���!�؎���h�>Y�c�8 �r�*^=:��JM`ٴ9�� ��
D�~�]�:�=_�w��O>�h)$�z]N��� @�y븑���|��r��+CX=;��_ȧ�-/^<g�55���8��������ڛ�nuIⷤxH�2&�v&�,D��r�+�T���K^��cn�b|�"����l��ǟΖ�s�����G�'��
P����A�P�Tƽ8_�	����H��y�&�r:È`�]�0� �	�HB�*��]��-V��L1i-����V�zߺ΁Й�o
HR���4kE-=�2.��У9�{�7*dgo���Q{"Ϟ=%)��՛�wM���u�1[�3�涱O����tn���BL�Qt��f�)I�A�.q-5���z�#�bFTzs@�)g�j����&,5i�����s�8@<pGj�߽}�9�HkZ�>gچ�yeݨ ڻ�0Z�z��M�+R��t���D��]��������335�L��#K�t��9�i�����'*����1*��׵�c��B���+��/>��yCǕ˽Gc'(c�;$(���YQ.����o��!HIIz1�/kz��y�r��}��R1c�-2��EBH���sxT�|�h�V�*���E�NcV.����l�Dq�bGY��`��^WL*ݫI�7Uv��S%����~���ԯ�����D�J�.٤P2���bL�C[+��lء/̉b�!���!,�d���g-���Q�����s���*��Q�S]��
έ�nZ%�ml��^��߸Ȇ���)]� S�� ��n�.
cھo+��	RL�qv1e�L3������-�ς̄��Uض��x�i���t��S�_�.��B�JŤ�$@�4O�0�bޠ���.+IɤMv��5=Im��ɥ�G��옇&����'tdy��rq�@����z���&���ڻ�8(���� �c� w� :��2]52�$c��=��;�D�5m]8 **p�K�k�k[��;��C㕥��H(c9�ؾ�Gg�>��s��"L��4S�$��Ĵ1KS��4�i�ǉ��yJ��K���+��U�.n��y�͓��� �/���[���zࣘ�Rf8=z.��ٟʗ_>a>4�8�^B���^	�V��h�j�Ә��,uo���P6����ߕ�>�H׾�3gJ��z�}�8:�MEm��:�ֱ�"%HQkx
�߿��w�����uCe����_�&�
R�XXx�4��EϏ�T�(Xl�XoW�f���f d�:�85.֒lM�Kk��`s!��Y˗�ղ�^��|�':	f|�^RRpQR������<VЌ}H޿#k#�� )�#�iΐ5�i�>0��9U~8�O�B����P�4A�ko^���/��`�t����ݣ�
<�����|.�Gglw�k����bv�Y���y
.��B׊[w��]��_�Llid�Uv!�C$����R����#����ԗ�Fy'�[����/�R�M5j��}�h��eei.�
��`���K����m���{wX|>4Q��rj�"����<W;��M��~NZ`ڠ����a�ݤ���u��^������1�-�)�cca=������8�BDoA��$Sv]��nޕk��p��t��)%�I��d�`�'��Rl��ǒ�aE�.5���x��Y��O��ds����a�v9k��g �	=�hI<],�%v�b��3�)1��A:����DN�N�'�/�r6��w���y��ߒ;
z�-�-�t��NVX�u�i-E��eݭR�|��~X�(��^��:�d�lbc��j��荑�rw!�����D�4�;��Z��GtB��9H�V֠*f@*_���mb�T�۲�eV��8����^�L�ō������\����|6��m3�����'�ը@י�u�H��H����4T��5�t1�����Rdy������weG�0F���e���4��\����@�Fݺ��k�������%`f[�.1�4V"c��=��fh^��?�X���ה����`xKl����1!q�S�2�Eχ�\D�����h�鮩!�۳yh>��h�~��Z�����n�L�;��!X�;��rs}r�������a +��p�27x��$�h~8�ъVbΖ��_ ��^`Mˣ�T!�^U��Ԙ��2p$���"���$GWXG	�-
փ�^�lu�b�,奈�Ȯ3"1�n��-��e�y�HB��o�,�-�����������$�r�:}$��*)vY+4+��߿N�~��Š��h� 	���C�*�qЏ�4�]İ��S<�跏�x�J<��`�̀K��j�c2� �Q��N�8i���R�|���rްH!��X� P^�U~A�v��>_Q+����t����N� ƶ6wx�
'�(�$Oĵ�S�Q|���Y&�	�<�Y��K�CWѣ@�G��Ia���;6��c9�M�m �q�+����7.��L֕�.�̬����J%9)J����e`7�һ�8Wm'���׽�Qj�L	4��]�^��b�>~,?�?�Ac���>�66��9B[BFj�������ɷ_{U��{ g�_�{?�ioss"35pvxH�m:q3t
B`�_c�P��+�|�`����������\�u�D=SertrF�����ɓ'��+w�ʯ��L������%3�c��@��)O{�/��ʔ�,�0D�R��% ��e7O��K����v�k�α�{;&	���E���"V�1a 0f�����=� �g
^0��?B㓲X�p��,gG�z\=�?�~悝ĎU���`�c�sx�= z��v�����=<���Tc�My ݍ�=�q=<>S�`��gn�Z����E+Ν1�ً��(f���!��ܾ�2�R%�#ځ�.(O�E��*��)8�7���.��o���{��M����ɥvr�Hޱ�:iH��z��B�D�z0�������F>GT����'�Y��c�&Ye?Oo�2��+Ё��cA��x���\L�l��D��z�N��]���c�?+R?�fa:/ktόX���%E�s�b紞^T�Rћ��$bΙԐ![��y,~(
�b���mgwK�M�U�7S���q�T�sF��`)hG�ё��X�YQK>�n�}����j�|���X���C+C�|�=��H�ӱ�9�C�e:�ڧN)1����s'��Zn�v������\�ݝ}s�h���m�狩̗3�p`����lkU�`u1�S�kUl9_�r�-�m:�j�ϔ{�:)a��-����9�Ka�a��������WeC+?�9U@�֭�F6^�]ʼl��H�U7��E��W�*c
'��-�z~c�f���srΦ|sÑ�̰��b������ڈC�Z7�z�;�����'ɾL�0����O]���w�p�Be���|��]���F��,X�_�wO��?�u�M_��o�΋���/��6q⡏�*��0�⋧���!��L�)��*l��#c(���һ�=s�:c�	^�>�Q�N6vHA9�pE�`�P��r,�I9R� �.���A��Q]�k�����\V��ĈPwn�U�Ҙ��tj!=z9��.��\*�~���a�PF/�zbs�aao�Rb�g�H�\��L��6 ��bA*�|O��.Y� ���kj�9�<�aBUmg��Yy/��]?��d��:��p_KEWG�I�����^�t2�?�m5f
�H&�Bϭ���D�F�?���v:'�[.6-{�v휊���ňE����r�QX�������4�Z��>Zf�H �h����@�2Çfi�N`F��ƖU�Of=���u�bwo���_����Ƀխy`��me)�K 0���O�y͇f�[��-�%�(�Q�)�D����5"
3[�Y�53�O�{��P^(�C�WՈ�l��ӄS۾�s���Px��-�@���(Wc*ȍ=���ű�
I
��d���v�U����J�FѱG�u������y�on��ߒ7�ch��燌��<8�.{��e[��gg��}S~���ы���ǟK3k8oS�۾.�ױX,\#��C�E�s]���YE5V{$C�Љ&��n��gB��n	�yk��e<������ �c�)��^c�7D)7КM��ɑʪ`C�Jr��r�|Y�e��uֺ�9IH�A�Eo^Ԑ��.�V��{ԒV$�ot���w�(�<::��7o(�^Pi�����`zd��Beh�4<Y�D�ѢM��щ��U�Ҩ�T-���G�*y���b���[��e'�*B��p}Noo��s5H 8�i� }Ό��)�g������)=D"=D����lx�=�sk�c�@�6���V㑮�2F���.<I�gt�BQr>�%C#8%�"������o*�L}f.����>�d����Uan6��h��Bav+�)Y�f9�g�h�1ĕR��H ~`��4���Rڨ#ht,ZE[?�ۇ�mv�C z���0S��@�њcid(���S¿�q?x� խp��#o��T��9�r�Q�����1��]���A#�~Գ�>�{"�^�F�ў`��o޼-�ܹ#���R��mi�Wyب=��٫���F�pڧ�֐ ):�!� �S�������px��3�0`x̑VWVS��ROJ�S��u%u�:�E̤|}pm����wn�/�~[. {R�ƲQ�4\>��#�Q={��oO�	a��.�&�y(�ޒYd�$�V�҈S�Z*���_w�)/�]���ea��4�3tM:f�9��Y�j���4�v�xN@HX�E��&E�Qa�� �!�������kj�������(�����b}�\����lu0�zF�S�qv1�ǧ�4��E��h���L�
u�!����[�UxK9��e\�Z���0��t���C[�4�wz�,���m�����z�v������5(�s��vê��i���!!� �]�7���)�n2� ���<�f�S��r�-p��*;UF��,LC+�\�9׵�1T�����S��`{�(�QT��&�`F�<N*SŘ�.v{GIBw�z�Rᵳ3��]�6/b^pgES���Yi��8��'[�œ	s0ť7�8R�Ώ����D6�R�ggʐ������a��M�3�o����� H!B.9���Mgrv�B��si��kjTj䀣Sw!z����{�q���f��V�������c���%M*Ǡ�Lg�h4�F�����޲��Mh��чy�>�L+,�ь<3�(�$LY?�%�����[�d�5=�W@�%���i�2�*h
�hؾ�E�2�#�H�}�d`�����)F��`^�7��.4�Q0�p���m�R��u��F��m��WH��g�Tr��5��_{�y֩�<��1�8�a ln�и:9���1N�8e���y��1�)��v� .���ޕ����,��x~���<z�U������_ɫ���.���Ԏ�r�{z;KM�v�k����mp�	|�9,W���{��u���T���W�Hx�NF9�Q�z��W��s�ZJ�#z�޶��zv:??��m�<v���aDm�(�4��NA��.��%�j���¾v0� ����h�A����/���/�T������&���\��H��,���5c�4RZb8>X-ƞ1��˸D��:tl���H��)�81U��v�h��,��rK3�MG�[�:��[�*OmZ�8�¥^ӫM�j�%�N���c�uv�=�����љ����)��F�����o��($���h�N��Hc�̅<���E���:|�x��+����1]�^��*���'��r$�P�ئ��ݙ�9a�֘� �0$�q�Y�D�ݲ�FJ
�]�� ��-��I��a�w�jx�xF�\i��F�5ޤ��o笫q�hm�w ZG�h����u��ʣg8������y��Ag)���*��gӅt����Z�IB&t4�>��L��7ߔ{��)_�ĳ,���?�g_|)m�i�aG��7oܐ�vO��t�������@A:���#������'��koȷ���ܼuGe���gJ��hsK�T���B�^��I;���������7�i��eŚ'8_��n�P90��������҆�|x���?|�c���^'ʳ�z�����c1�չ�_+z&�����67���#��%���
ͽk져q󝝘<t���Xk�׼�Q���#F���v�Fp1C�p/��u<�����\�"{r~�~g�'���飠a�n0ki]NF��u'O���
��l#�c�+��-p�F�3���V;`�y�!X�
��u�]:9҄SӦN1"�~�L!�ՁQ�-�z(�=�C��f����QY����ÜR2��'�7eU��c>�=�m�0�����!D>(e�b3T��M�t����;�A
BFb�q7�J.�����1�}��V�w15�
b�ċF��*?,��{��[�(S_#�E����C:99��
E4��c� t9�}/��N8��zoe`�ӣ/�O����.� �O!�` 7a@�y��%�><e'��	t�9U��g����HC;����]q=�'�ـ�p��v}���:S\�ܖ��g/w�`��lI��1D��|q�T���)��]����vr�5�6�Vt㱁G���:QbBíy�\�4��ּ�M2d_ɗ�h��JR�Nx�5]򲅈M@\>DĠE:�(�����+mA��~  �
��lɯ}�-������O�m��!�|���S�+a�G7�K����G򧭥���H�c���(,�s�.����x��]���_a��O���$G/N����j
B�� �T�{q�ڋg�il޿uS����4��ɓ'r��؝}�Bi�Xש�cW�.��^Z��9��V���©�����"8Q�����Ö,oxe��H4��g-�CQ6��@ ��P�(E��Nɭո:Pe�?T }�Ӄc,G��k*Y�k��,ڠ��^j�6Щu�H�Y��k�e,�O�KH�B�_R�t�V�O
�c&�l��0_���:�:j` w�^ɲ*	|pws��Ӭ���c9��:B!�q]���آq8������ ���a�c'���'qƇ���n٪հ��ؼ��rS4��DD������!�Wp���$�q�{� `�P>>�w�K4jQ�l�,y��Gbd���L�.}t���jz��a��Ox1X�`l�ַ 2�.)V���hj���鍏[��
Jǅ��:/%���c��<x	��!������f�3����A�IH���=��/]�>�o�3�����/N���uPܭ���&b�!_�BXKw��N�k2$��U�Z��v��˘_pOѹ�1�L#9��T ��M�YN�T*��h;��p� ����?�@�����+�*������
�1�;w�Ҭ�G[�T��<�I��p�kE�ԡ�r�@�����ۿ!���������;��>�S�#5Vyl~q��8�.ƅ�j`T�5�@f�H���s*ʒ����D^}�Uq*�>���l;�&	c5�G�6��G�O��f-��1}ga�;6u�2�_Oe&3��ε�-�9��n3�IJ����Xo�"'ġ:�Ve�,�MK��/yL��#�2ޛò��ո���T���b3;�����yE~�t�_\f�����?|��a��o�:�F���,�lł�y�yP�2�oOe2�R#l)9=��Q��jF8)����O�>��*����c�a)s!m� ���5=�d��xKg�g�R�IM̫��b-�b�5Oeۤ�E�v*�e/񬈹�:�ª���-��PB�f�q �+�ay}e}�u���+HA� !���L��[�U�Jf�E<r7n�14�`�7�ĉ��Hb!���jf�\�+C��o���2Uk���)s��壏?d�-�͂�p_F���NH��5��7)8�w1?��~���c��&��:6��(�y���'M�W����{��Ɂ�3~r�B΂E����&�T�Ԗ��)F�m��d��y�����ڝȎ~U'���[�6��;��¤��T	_�/��@~��r~�d��u��씸>ڈ���j�G�YA1y���Eꎵ(�*�C�~�֑gKڋ�׽�l�h)$I1Z:Z�{���8��^c�B��}�����!��!�R�����ZX׃����Q!�nmPy����3�����/~&OU��q���
��Q�h;�SYUP���U�q뺵�ڔ��=�v��"�_�jb9��^�~����F<���9(.���8r9���l}o\�F���/������(����6�w����z$+P�:�i]"�Ν�C*`2��?>�qJ�	ki6a�v!��L�C���X��ʁv�/�8,�F��#o�����B� �q����7mo�$Ǚ\�zD䞵�� ��lv�[�HWf2ټ�����9���ѴLj5�� �V �P{U�q��/"� R��$�X��\"��?��Ǐ���>Vg��6�̐�m�|,�ӐB# �N�"�l衩_%d�>4l��)2r1����)Q����;|O(°FbjR���%����2C�^q^8�o��[f;]�tЄ���d��I�z���T���kw&5(@U@v����)�χM+2��3�syZ�a�,���Qam:CP�![qg��65;c��#��Y!�X��k��y�x�p�!pbC��P&��b=gsky�Q�G�B�	@�A�<�bN,Y�t��^����FZ�:W4�|a���"�:�9C�7�!��FP��	"x�%c	E�l�{S8}��!�w|x ѤNg���YǺ���e���𬄍�^��T�pn��������:��/ΌD';p�s�:��E8���.j�� �^�-�jU��(�`�y�"X(�0���3{���qt|,?�����آ@��3�o�[�y�`�c�������E��qj��k^�m�Q�f���h0����=�	��@x��2��LȽ�{� �&��w���Ҭɽ�=�lE�1�l�Ĥp!	�S6KD�\���eG�٘��tԗql��t6(����G�Ͻ(���5셣d#S�a`n��׭������b}�cN�.'�e�K�Dm�(J�s�9.�
�QY���T�f��A'E@`kè����4E���|�y�(�Ӵ�&�f��7}�?���G7nܠ!�Y~�������dv�ӯ[I�3���6R��'`̦=�����bs|x���g�\���3�i��2��p@�q=h'	rC[3C󓚧�C��s�Ru�����Y���#�D����'��Ya�鰺�z@�A����	˶�־\R���k����i=lj�b
� �1�aK�̥���}�ۉ��|�ᄄ���� ��HIY[_a����M58�p� 	��7�����|��Y��ݷ�ܩU�z�H����O�?y,�O���?D��)Kp���2��hvH`S�����@.,]x��D��&�uD�z�$i:�����P<d5	�������ĕ.<Ŕ4� �h`�{�C�[vD��S� ���n�t���׀�2����o?��gh0��Cp�w< ���҂,�Z�k�_�W/�!����L7��`��č���>C������D�m��t��)v-�$.�P���P��p�B���?p���^L���������z��e�3�f�&֧�B���Vgx�S��_�8^��k4�y�*�/�dөNjtn����9{��ױDӉ�-��v�m�1�u\��.��jj �Բ�n��v�����t�=h�||�3B�#�S��'�tt(�O��px��W�x�����c;����Ɩ�	J���wZ >�MvN����'��]��^���}U&�>O\>/�n��a�*�V�[��״a�yM��'������_R��/Pǿ�,�uI确c�ZX�͝}9нp��R��MlE�A�6��tW�p;Ѕ�l�(�:b�!5���B�]ak.g�P����?:�8L	�L����Aj.�(�Aj�!?�v���(�D)|�} �����]د��PG
�-�`�ktM5$)�Gl�Ŏ�{Z��KZ D��OBG���=lB����,�s�ߛ�8�kAaD�x(	jJ�h�8b�T��mAO鸄Z:I(֗�p�C��"�N\���҇�ڗ�����um��B����X����S�ڕ����Z'�{��tF�������#]�CRA�IL�{�����N��2�Y����ֳ����I*O=�/>�S.u{S��c��'^�1x���u���(�NWV��XL���������I+7�
74���4�<Sfzj���3��֊�s���+W	P��Cf��V(����<��g'apرa�a�,��rK�j2hx��#y��1�AIM����׺>_jx�"���;�?���Y�K/�3�����uP�t��O��n�{ǲ��p&�n7��+������!d������ܰ�:}���X��}f�����H@�0�o#R�j�Q��t(<�(*����t��r�S�� �O���:�8���(5MS?/K������Upo��L�]Z�1T7�4�cd�5w;�3kF	@�Z�ao6Em�Բ�l����L�yAOF�O�A��:��%B�<���9݋���d=�������f��W���7���q:�b8��i^���ҵ���(h�<��S3�s�	ˋm"���Kb�_;ٚ4ޘ���xp M�Z�8v��@��4w�%�'�bCNӢ�;t�ʍ���4<���TY!�<��oRy&�g5C�p�H�;���0^�F�,�k�AEz��S�p��;�
��-�W$o����� %���*�_����������5 �"92�B��aF�IG�˗�SOyu�%�|����?����oh��V�hu��<���n  �q��u�&�O��aH��Sds�x4jF$�u�.��n�� �=X.�=���a�}~2��b��i��I�RQ��0xBZ<�,���~��Հo���v|C俵�ˢ:T��xA��Qc����[�|(gO_��}��������F㬼�VѠ^��4'HU��F�]��ʜk�"h��O:�|��+��?у���q�LB���T� ?�7u#�Q��e-�
��Ad�u<(\("��d�� D���Q��vt'��'=(����@qqq�Z�gN��%]s�^���ﾕ��O?�Dd��k7x(?�ڑs�Oi����Ij�zX������hp<`�1xUQ��ً���m��w�-�������]v��ȣF�6���4�gQd��濫��&p�}��H���R/�g�s
�B����9�r�	˭�<s�˘'�&Ȣ ��C���_g�q:szU���z&�U�����m/��QCbcmTHvy%���I4L�'�b�����bc'<x��"��
����m)t�A�i���������n
'٤i����Ñ�HVRɨ:�k���o2vj�pO��É��ȥ�B�L)t�:y��,o�s{�RW.����pY�2�7/���t�x�ǩ:xGꌍ(j {UGM�Au��A�&�o�~pb*�˯ٜ(֢Df��5E!�'/Rh��_���Զ�>�:�4�g��7�ɯ�y��OA�c��~��pG���h vȵ�����s�]�<Ks�~S
�+�<����O�e `*��ر���mz?� �a��(lյ�� k�����2te���:�ŵ`]�|h�@?3�QZ�u���P�w�I���rM� l0Eu�]�z�ܾqM��}��塞? Ό��L����=fl��3k�#�۴Ld=,X��ʉ>s�Xvv�������> �}�g&�������S�tϩo3���s8�m�B��I���2�5P�,˩�e����>����A�����u�����M���B`Gn���#�a��z�b'Ķ������&�I��u�&qI���1w�1?! ^��V�r53B��xڀ�D���Z�,���B�İo"����GY�)�ٷX�z�k�V�vT*QAa\�O�n�E�D����̸?z3���z�Y~0�e�4�uB�6�*o����0�3���7������2ʀ��c�+Z�\"R�#�tLf~�03��&8sZE�b�S�L2���_��RHG�Q��O��Hwg���A��iȩ�j�aga��@#V����`B'�%�D���z���t�V�@
1ς�O����;f�D�"���R���2��mF2\u�Z����r��eY^h��o���������:�+]�z�(��	R�N���|��T���90���ڳ!sQg���5��~�� ?5��S��<4�Q�`��"�Ɓc ��-ؚ��\zr�3s�5�4�P�����Ӛbmձ��s5�袝���B�)W�����;�{pȱE&ƳYoK�]���@~�������S���������Yj�"�qƼO��]�`��N'�%�j�~���5?t�)��?��xM�Ġ[DV��"~�1�Ŏp���Ňu�@9�iz4��j��eo�Rd�0�M8|��Q$������*� ��:x&�.��aoȃ%O�0P�����ݝ=iw��ܴ���@a�k�Ro�RS��YM����������bB�r���x�Z��6�'QĈ����)9�q݂�����_��@k	���m��)2��U�*�K�(8��GdVD卺�J()��u�F�aG�߰^���h�jVl��j�e���i����۲��"�u��~�ߏ7���J�Q�x��EX����Fl��:	�#�~��"��&�Z^��g���ܙ3��k���3g�w$�|��:�yº�1��i�{�	�,!��VsGsۈu�q;<<潀��9 ꮁ��1���Ƚ�y>�Cq�����<��`뭻vx]�sw�oi�r�o@�;� &�V�*�U ?8/X�;c�����l/J��0�1��VD� eF�VAT���=��&��%~���[}�"��W��z/��
@�������  �H�3V��έ���;o�cޓo��J��LGC����1�{����qO}��$'{lYk K�I��hϚJ��46�˛�t��w��1��J��!0B��M6
Te�p�5c֧�e�QX?��)�
���4�&�X�Q�]��4�iB�gc�v���Tv���c;[��QmS,��s���,k�ϐW~��U�nC�$t�1�X�8�<y*ߴ�l���Q_�u-̍Q1J�L�AE��^ֆ�о����)�[�e�����G[�2щB7�Ͻ'�0P{�	|�lO�ҔT�A�7��݇2��r��%N#���)Uhu���<<�aSV��t0oN/C�a��Y�=|�u@�!�Aj��t��'��v�< �K�'2�W�*�]��C�w΋��Y�৊��k�����(���e2�]�t��!���sT��hu���X���Hl�:%7��Mi\��������d�i���H�����l��p�?��sS�+�l��ENM�9���������6���n��I����5]�J>��&�_-����q�&6��`ҎV��C�[H��X�a��������~䳒UP��_n�`$u�)����v��e�8c%1&
�q�U"�u~.DO�&�V4^�Z�(�F.^+�N�7�"�# �n.:��z�T��3p�353�����x�ܺ�)7��� _~�l=}��j4(`�
�uSR�a�E��a�E=+�Q�8.�7/�\�e��`gyiA�P0������@�༇B8ތ#S��c(��U��}��q��8����"�L�f1[B^dfd���x t��K^[S���iY__�u��w|5��@����t�:r���g�W�G�������^�Vٱ"�t��^b3"=�5��C[��;UDΌL��	����~�W-mnND��۟$��<S�bj�t��D����@�%���Td\p�mn>��m�G��G:��yhC���!A�S��ݽ=]�C:����Q����,8y���l�k��d���l-2@Jg#?�,�L\n���8�����x�)����Wר�`HO�2�౮�>�αHK�_��ʚ4���x4�a�]N�$B~�/��QTtA�	�_�����~��g^ynZ<�D���@p "[7MY�Cď��6��{�!�8��;t��:?P�Y]]��C�S�tAH��dF���t��Y�ĸ7�3��i�p�`Ϟ^�D�3�/4�;�A��׮��?��#;=r��V4����Ou���gAn�m�;��Cpα��vv�q�h{�M�\cE�(*t�C�l�a7 �
�P�3���<�]"偪R�1X�j�3����|�������z³�bc�'�؜�j!S��)��
�|�͢\���ٲ1���# �%��ig^o�)9)Vu��霯�-Ȼoܖ�7^eM��_|.���<������׼�gƩ�%�㘩��,#�#����X6qW�<��#['z�P��C3�!).B��r�W��ȶ4h��Ph�c�w�E�tdo��~#��y�@��ͥIJ�H&c+��c��֌[��&k�2��HǙ��Cy����Ɇ�~6�#��3��W���7d��9����~��]67k��F���6�����+ ��l�H5E�]���^�>z�`jnxr�`Q_��X����xi��z��?xH��>>#6�o�x(�}��,l<��@{qE���q�ź`7 |�Q=�b��YFg�^����Ԃ2d,�E��L*��}tao��-�g���L�.� v/u�c���_DU�����?�*�c��
�"����m#��=�)��+s�ޓ���I�2��xLR������M_qj��MYk�Ks����<˾��x���@�z�6���E�57�9���4Sy��Ҧ.�-(C-�*]��Hل}�s���`lQ���qZ���)�7��K1�s�{H�S�%%l%Y$��	�ԤF�/�Hl!�r�~�t�+��p�!���d��+��#w��I�(͙s�3O�RA�j (�H�����0��f��� �7��%"��9'̨ڏI��� p6=��9u��\<'m5l;O7������),5�L/�����X̗8���!�n�<��5��3�;
^@K����W�0�k�ۦfHYC:
!riMT5}z씝�P�6!B
ѠZ�L�t���ؾ���'��@�	�Z)����a8����<8ܓ>R�{����Rt�<��?=������w���k4�;�;r�+Yt��1���"��)UC��sƆ?�����R=��
G���,+_Pt*�p|"-^|�?'����)�2�k��đg���$�#h�"pA;v\�ӭM��|F�/F�H�5����H�s2S8��m7��C�@Z�R�&�ը@
�Kk���������a/0�E�2�NkF���psS���ײ�밧N�u�[��KW�i�T._�N�4��^C7ƥ��vM�5�2�}lJ�gn�|B���jP�J3�r"澙$ZX'�;SWw�F���s��T&�eIc8��ǬEX�����Ã>��4RA����,nCZr���)��:�z�J��GG����:�y����c�m����Skµ`�;�{dL�A\]Y�������N���zA�e����g0�7�$�u�k�"��D��ԊY1�x����w�D��V����a�s�H�c]�w�9���?���
�&%�Nyפ�F�;�! ��x��>�
 �K�oYw��le,'A, #p+@i�.9��LX��(k��ɏ��{!���HY[#�"E��ы�$� �i�w����#O��[M�x��7�n���-:r������O?���4����5�䯃R�3i:��D�j���yFR�pR5�GQ(2���Q)'�{k hth*RGٖ7r��z��B�od}�����z��j3�MZ<��{��D�
 �vl�4'����ԋP�9S֌!�����Q[Ԣ����u"����v�tt܆j#��{H���/���V���ఢwCn�{�(�7���C]��ѱ��Y�E�P�ʼ>ҹ�K��P����c.{4���A�)�c�����5	g:�ȑ)B= hu��ɭf�h=Ґ���bߘ���V� &�*�d��sn�Hǣ7�(Ʉk�[���{�yݴ�Ѱ�}�ܩ8���;W�EN3*Q��?rM��D
5ۋ�-A�Ҥ��?�����{����S��1�^G<)�A�rIי����BR<P�h>j�^qb��$Nj�&�2���+rn@�JJ�����֢�S�e��MFq&ƑB�-[\��:�c)�7��E����8
�w @�/`����.&'Ԃ�h���e�	E�F�> l�l�FO��J����gyT* (��N�`׭����c���M���U��^��6�F��g����)Ӧ7�J3{��H�����Rk���E$����yp�����^+x�τh���С6T�&���Q�H������Kr���s�M�y�u�x�SנӰ=�o8P#����12Γq�0�Xv�Ww/4�!DEW=A���
4*'_}��<z�N=�ȧS��ǁ/Ph��h���O��6p�h�E؍��F���_��I����K��o~+W�\��F���x��k��8��,�x�"��K۰yq`s�d�HT�p$�8q?���Q�C9��q�����������78�XӓQ� |���H&��7�Ӹ�7�׮\b�rkgW�CwV�V��+z�f�T3Æ/8���>w鲬�:˂�S��<~�����@-c�P�u~�#҂�5�Ngq�H�d:`�z�T�;���݇����<�|����=�;��S��������%a���'�"Ϸ� �x�\+P?�\��~�1Ǜv's�#)l^�S�ߝ����<�9sYn�e6Y��N@�I-@S60U���!6�]]���#Bwi7:�E9}��<�;���:�����z��j��Ĩi��ޤ��<xrC눉�8uf]���,�S��u��g1����ST�U��@��Lp�N�����)�@�i,F	i�;��;��;T:r���@�ŕ`¾�t{v�W)�U��|9�ί	${�Ө�/����{HQDG�G�\d�@=�@�$�����V&�;�i�i�P�λ9�6/�b�-Rψ�"� q>s��zG[��^��c�f��O�^�w޾#wn�F��W_~.��������=8���:���9�>�L��AmI�a�q2^��%P|�=���e�S��ș�g�~!;C՛�5o�`|����d�$+l	h* �c�0z��-}л�|$�,��~ܱ.���)!����L�z�u`��:3��L�C�z��=nE�ʥ+W����y�>|�A�Md�ϔ4�,t&B6��,�A�,�Kl�4"�B��!%K��t(21�[�e�h�.��b��@��D�d����$t���&3��ð�b�R4a�w�˩�z Ml���1�qΚ��z���2������j@��r�Ù�~j:���r!sڴ&9^X���$c�s�rY��%������q��v@�34���C����[dg��|�	�	�#dm��	qP,�'='Y.7��:�o!�8��H�e�"B�b�$#�(qB�1�ׁcIt(oM�y�.�S�(�J��L��[M?GfD�i���ݚM1�%���F���
��A&�ܢ~F�3�Zj2(�D�p�*��Y��
�&)�����(4ik��!�BhF\�qF��t�th|�.�?5�8�´!0p���Su �Xή�����[r���dkS��l$Kz�� ��hқL�� e�ZEN4Ȼ��S:�H=.�a����~�5�y�\�vU�\zE������5�����V=P����]��K�`� �T�̘����meu�_��=�^�&�����ݻw�Ku
����<�CoU�XǕ��cC+��3J�5m�A���s�r d�7���iAV�`Mw��9�}��ܸq��~������G��ѽ�4�����I10���G@h<B��N{!Q�`׊c,H<���7����NCgHN~�q��;�n���!8�P3�W�����jL�z:Nǲ��ݩ�g��'L��ZS��T̀�t�B��=p��.��S���ݹv�W���e%_ၹ���Q�����@!�C``r��4����@����s�t�����a��v8|�׷C�T�>���{R-h��^z���n��\�-��,%b^�c��G@j��JF�e�{��H�Wy�whT���K��4���^IU�-��#{t�c��vaq�=	::��OѮ>�ZU:���k�nʫ�o�3���T8���8��>;��&C
��%���z t9��_8L�"�/�\@=˾RX����t����rҬ��
f��O���,7u�L-! ���6ԭ���Y���P,	�yf|X���z�N��I�#�`�	+kW���4d>?��$c����B��JA�#I\"02�"(P-t�#��މ�uP��-���sg5�j��p�(]ĵ�z����<A\O���^���(�x�v&8��S)��9�2�a����v䦞�����I>�����?�֓G��yR�yK`��8��`d9��n���0K�)�;���]Y[^a1�=�� �:��j3V���3!0� `6��8������tal����#=K7���|�%�=���mR�h�"�M�/h�
�d��C��D���C֝��m՛O��n�3g�ɭׯs�77�3��`gh�5�]�N�lf8�4T���+�W����nҙI��G}3i7"�Вt����r�ČQU'� �H�����7`�!�%;�:�ŧ�U�c�q�@�ʄ`PL�����)����^/k^F��(X��|�>�i��{m %��A</���t�%a�PJ�GY��y�{�Q�������[�x����:
Ǳ���E�=Sӱ�o�7�nw�Icvd,sLik�c{i�~�q�s-k4ʬ�ϫ��	���;��qř���J�N��,1���*��61�B�2F�k%4Y,Q掎i⚼�#	�F���<�!�[��ȣFF��iF����~�b|�yDh:�X�Ylm��>�S>
�U��؏P9dk�ŝ��M�>��H�!ZB�ה�.��ic�)1d�̥���u�f���E5vY� ��34���J���u�|�,�������÷��l����n��3;0Φt��;�p��s�Z�jl��QÛ7o��o�-w�ܑ+�_���O��`D�:�OLI��4/�b}/�n�8��yV8.��6e=��<�̢�)k"2g}j�1p��9�~Fn��&)5@����k�ꋯ�,噦-6�²��j�Nsd�L|�@�n�s"Qo/QZ���( ����?��R�o����r�UJH���Su�ՄBP+�٭�px�T{zAa�QL�������#O��ZW��JJ�J�Ƥ��*��'�'6��:�&U��D���@{�_�8��"�2�S=`����@��1�P�G�vkw_�  u�7��+�w��>�˞:m���w�R;f��L����Kc�3�66ecs�Y��������դ�������2dU��C�E�",���x �yhD�^0*N*�IjB��H�e�U¿"K���?����.�y�_|M�~���d+�Dz��F��糨]x �`>p�O��2)B5�(`�i�P�����4�t�{�m�+:n#�Ep���h�Ș���MK�.�N�!��C���5�y��tKj�����op��vb����I��@&X��\M��%=`l�?uڑ�Q�*%(��x�����G�m����8(A��Ƶ�-���:�;�53}|S�IX`����7mB�.�;��%Ś`f4-�0F?3@*�K%��ϋ�����1���gN��<�&W��(��iړ��Ӭ�@���t_�Q�g&:U��#��Ϭ
m�8�"����I@�CvB�ָ9�jy֖�|��f�M���ťEy��y��u�#�����O�M�5П��)$�չ�� �$>���{䔥ܳy�b3M��s�,t�_#�r�իr��9{��
���^����#��hW���k4zFiEfZ���5L@�/]� o��&��w��gǃ����ӧr|�3��f���V�=Ã{ � 2� $ Z�� I����U�b�׻��H���?��\8s�ぱz�t��nF����لg+��v����S��Ļ��~ƵA�5/�o8}� z�Q�J3dJo�A �έ�~-��U�u��Y�ep#��⁰�� %q����]KH��
{Cue�O�5x�x�lf:�F[i@k�o�1j���ِ3���\
�Arl��s�Ӭ�א:;�ਖ;H�ԻĲk3�94g���qj���37z�%r�b���t@=
Y�Q��_ܦ��K��Uڲ(�1��U�r���RqV����"Vd�h�c���	���]X]"`YfN��ҙ7lHô��<�f2�!�$)+F0��i���-�(��,#��q�Y�,!���u�E�9So�L�
���MԤ�y�)+�vY����A�4��sF���GS����L=q>�^G��R��#O9jŅ�?�x0���h�F;��d��%y��E��=|�<�Ov��M���ԩ�$�����G�{S	f�t�ź���K���GjL�s��6=�a���t8HDb�&��T��0�t�U�y
�|��UD���H�q�_�f0�4���f��t�Q?��������?�O>�D~��#�~oʍN�$(�ԅe�ي�d�MS����=��� �m!����e��/�Q�2��޾����E�#������e�V��� �Ex�پ���|%P�|U3H�f$a�EN+��iUp1;�2ZX�I�@-���cN����s�̳�T���r�������ɿ��<��u$��Z�
7�G�f���F��x��X\Y�[7�`���o��V?� ��s�����ڵW�+geY_�d�H~z�L=;�t����b��"�%�PL��e˝20���z[�Hz8��d"�FϛyW��y��<7V6�A��ب8@ʧ��Ea�C��h#�����B���A�46P��(ϬO���ٹEuj�RB��$�wyЃRw��S�[����D����FGb M5�KDN��(g�e����<�P;҃T�F�����GR�r]��t��Z�bJ��d�8�.�<J�RE+���(��h2��)�9Ԁ{meA��ك% �ep(CJ��%u�Y��6��νe�2�Q��}	���>�֣D���P��{�P�;�`7�*��;ƾ�l����u�-���C<�u��2+i�Om��9�G{{:�SW'3KbN۔�)�
Z�]Sc�y�qe=�E!6ճ���a�it��>@�y�q�fA�5��Zh5�7o�[�_g#���J����e��#uXl���]7�޲�)�Qy�z�:w��i<�?#�'�����ܾ��$�%�������,*8�p�)q����9u�.�v�&��~��p"�C�Jb�^��;wA��kx��	�@z��!A���C�9���}��p�E�d݇�s�t䜵�X�nm�W�"��zC���d��d_��O�.0��Q�,��Ds�
z��,�/�Fb�"{�/�υ���&���'�;˖��9��ϑ�<6
���������%Y{*f�-������ ͜�,�֪5&��Oi��nWfƃ�C��[� �7v���fA)�j���Ɩ�(:���>Y��O%���85�;'
�Nsnj7���GN��~)�^�@��jόb��D�ăq9�)�RhF�9����@mX$�]��5�Ŝ��E � G�X_�Y�vX#��쾝��P�����#́I����|�<l�"]�CzY�}*xW&$��mr�b�l�?G2-ɰ��5��z��T��������qA���S"n���Ih��F"PM��K�f]�(���ԣCF���ER@R3��ߑ/��B3栣���aA�#�Ln�ߴ��R�\p�P�i%��vh,�����)0@�?�'{;�-�us�L��4�N���������l]�p�4�?������_���% T�GDݭ���z(� �icw;=�k����h!�~nr�xfP��J��	�acGH�ޘ׌W4��u�������0�����`��8���7��1h?q��S��,-�U�Q��#�~��7���s��o�W�~#:�c��SǄv��r�.��f��y(2	�#W����C�9I�q/P�"���2�8 �/+s�Pc�2��e :�^"�T5����a����r������~Z�%.;���n4�u�.�� ��ss�Jga���
)K�ntW�X%r��e5̆��	Ym��6��^����:uʚ�@VT���qO&�G����bu<���w�~�������8���2���2�Eb'%��ʣP
s��bN���󘉄���!3�F;ʠ�@��'@7l2o��L�B���X�'�
�s�dހ�!�b@�ו���6ꐢ̬�j0�&FQ�z���~�6&qۜd���̻�2�YL�>1�e{wO�o����ܘ2�c<�hn�7l�:D�)���:,�Ψ8�c)mP�M�VB-�fs�Q�K*��<�_ֶH��
�")�4���v������2\�:��ܨ��W�ӖV���S�o��yV��KǄ���r�l��z&Ru���/v��܃�	�����ϸt�ܾ~U>x�MuH��u޿��K��ڒ��U���;��0@��Ԃ���A�Pg4hs#;��ݵ�S����w���ߢX��8.Zԣ?����4���IN�VBDVϜj�Qu�C��*	�2A�\ˍ7x� �x�����x�x~��@�=ᾩ)���˨����;:�Z���G�S#A��3��;�x=�> ǜ����u4d�U\ǚ^����{x	M��c�Ҁ��� �I;���̀����V>%�
e�g[��@���27�^�f@��,�3���WB@��NY-���_����2,>�!���p	T�?DjKd`�}��_���2�{���f�Q�Y��5���s�9xpY�:%�5.�Nj3�b>�x�"�H�:�N)���v�a�<F#��#�:(��)g�-h�f:�� ��sHf<K*]�~с�$�F(c�Υ�kj&��G�H�4�8='��9#8�Q�&�i�@e1���qi+~�د-����3��9��ͅ"?�`�1�"+�3��@	��;�L';���Q�p�-o��s��\�g3x�AR��є�p,��Fl0��k+��Д������O����	]Ϭ1K߀�לJ�2"h�'��;�Cc�֛�(cwx`-�����c��,���A��H�R&2Í
��B��f�+ʠM���Ug0��׆V��<8�@<�A=ujM>��Wj�o0������?���?А*3fwO�a��� �;[�p�p�)=pPD�͗_�a�_��_ʍk�y-G�r���C���d���;)Z��9�#~��ง�#��/>B�{B����a0F#db�G'�fCn\�)�Ξ���{�<�_�:͘4��`;b�Q��1����<z�)��}����W�\皻z�$M]�gN��ߡ�C�r[�*x�lأ��]��NW�)eT��}R4��r�2�c��
�bؗ?�2��� �<��_v�mʿg�'�%s1��*"�NUA��M�V���y^�8e�5Q\�G�I�%T7���Xݯ���1J}_�R����J���C@#��YVԀ �gz4�ܹ���8�!-[k��|�eM,C�S� a���M���q��h ��-ϟdx�/���b�յ%/b�a`;�Y�=��j(DM��pP�(8⎒����G��U��2�D�
�?�/,e�e�s�d8C랽��x�)�u�����ﳎv��1��{zDde�Qp�=pJ%�b��;�V�۳}V�ҞS���@V���s��My���A���s���� �O7ȁ]�T�FM��{�����*�H���H��k<p	�7�~G����^�{�=��o`Ӱ�q������:�Y�0�!`?ύ�K�2YAz���P��9���9��� �Mu�?��S���������F��ʞq@l��	��\���$j�j T��7�C�7o��ɵ�7�y@��~Lۑ�v�����r��+�|S��YQ��I�Q!g��$������?�>8�S��s��7oߡL/�x�C��4��=N�l�5Rf�� �<|�k�������ϻ�R:�şQ��/q����p��}�HJ{gud,/o��7�&Ң� ����L]�:��%�� Mjv���!�v��y2�He�8�)�1m�^��R��������hp(����<(����z�<F~��Հ�<4(�&ƍ��"�䅩8���m�ek
��q���Y"�6,\Gˮ܊"�wjrci!�t)�z3Pb2W�11i���[�p<(*��&�:e�7R�p��&[�Ǿ��r�![����k�@{�H1��t���\*�o�yAU��8\3*s�hؗY;b'C蜣�Ғ�v���+��>�2�@0��~��E���~-����t~͢��,��AI���0��騛sx<���y<�|���v;{��?�c��u��68y��������%+yp�K|��ƃ�����B�6�X2Ź���]T�g�1���� ��G����dmeU=xX�V��Q�>����ϝ�E�٪�������q��KYhLS��`@�SOI5��߽9�P76���R���A=�P�̴�Q(v�ё�SY�<���f��9j�4��G�����]�ݽ��n�����\����y�-����ډ,v�$����~�d-,/�����3?=| ��-��=ٕ�������{�����ӽϳr/V���5�ҹ^���.~��9��ߗ����OR�AGW��&v�c�P��_Gd�)�)��<��E1nl��AɅ�p������7��9[� D=hoE�{&��a�ZRd�x�N��]��G|��f!0����ށ|��Oȥ�s^y�<~����$�vf�՚S�	N;�@)!1�sՖ�}E*E�q�����]�oE��,3g73�S���n��hJȬF���33{ބ�C}լX_X׈�F��� �q@�M�������޳��w�z�K��?d���hnuz�{�OjE��hOS9��&oݹ-W_�B0�����7_~&��w���(7�5����ӲK�-�>{��._�"��-���,1��Af���Y36�G�3pvT�p�� .��K�\�A�8QJ�1�x��¹hr�����o�C��:�}�<y򘯁����Al�X�k��M����gO�D4A<�ܹuG<ސ�6�B�/ �(�}�>�M�� ��N��г|hj3��5t<�\G(�-��_;�u�n�|]�}��=���q��~i4�s_=��,�?��˫�q�ۈ�����f�*T�_|�����e1_&���¿}N"��O�\S?�<������a��ԙ�X�'��S�I�@��*5���-Y��<Gn�iN����g�����_�M+^�㟡�d�J�Q�Q2 O#�TT�����q�$�Yi6���0�Dp��֯f����#�y�ԖG݋�|z� +"�L^��a SYh �=�!�hZ��(�B%,fp�GCC����b���:&���\*d�|�R�PhP�z���A� �T��
#[L����br	�E��<��wj)73�E��o:��ؤɞjs����n��#��2�|����
TJ5-�8G��h*++k���}�m������>1tk$
�X�-��8��!/s��gԎ�Z���a\I[VU�:����J���\p2��ݩ4x�f((vD� ��!���ۿ�[Y^]�������W��u�g���2W���2��wt$��1�b���̨P�6�:�Т������MLJNi@*��H-�3犿q:[@~�x^"�Ŷ:��-5}��o�ϡ��^}znHd��P^����/z������B1"��3�Q+1Ev�Z��
$�1ڍ�����^ϓgO�ZQ5�Q`�w���5��ƥF0x�6�7����5�Q��T��c{)�y�|_��uN/��`�(�!
�w1��{�^�S:E󅯹�Q/+�����g*�̣�F�s���c�ڔg��R� ���$vi���bC0;���]?uf�Q("��A&� �t�7�֠�M���'�!M"��^;�r_��um���w��F���,H�CE���:܋�n��p����WvhN�A
y&jN�1P��_�BT����� �ڬ	�S��TBQy�;���ȋ�8��B�-P�9ˋ�$�j�>'@����rS� %%g3��7�N�d3�@���W�İ�+{DB�|%����b����gv���ڕ�r�ګ�HN��O>�o��\�=~H�V#�Ys��k�M��AI�:��Z#������tr�}���G�!����@Gt�!_kskN9x�x��Ua��j���a>C��׆��N5�z�� W���>`�ߟ>sN~��NKd����#k8Z�7�ʬd"!�����t8a3@�V�S���#����c��l*�0 A���������ߕ��O<MЁ\}TdB%4������4N�V$:�,u�Mp |��H5T�P�r���3�T�zKu%;����P�r�EU`�J�>�/���v��sc��@�\2�%̟9{��
/t���H�j9�vKϴIή�uHdd2�3[�w�q�o�)�
0 b]��R���mz�s}f ���)�10Sg���x_����m>�-jÙotԟmQ>ܓ�L���	
���J�o8��� N�Y�K�(�OJ1���in"��όx�=Nz:�ƟSKF֊:fz�*�Q��Q'�]7����?���}~��6a�����RY�q�.�IweA����u��k�XB�U����&klD}ȸ"f`3����?B�u���d/��y#�ܹz���Ԛ��D�\��X��|��p4qx�l�b����e�>8�0����կ~�/ ��eX�80c�hDŁ��6g���ݪ3P�����tuX�/�����{��A�<Whiij){��Pt�D��x|�&���/�w\7����ԃ�l�{��,x�@ӀICW;�X<l�!��k�4d�x�(0+�/���wA�q_�U{�|�G0aUS�_y��/f��\�T�;|��ò�Q'-aLT���j�5�fC?�b�.$�����$�V�u��N��[�GB��Ç����,u����cl��v��4-y�V�����Wc��촊�L���b=�}Ԧ̜���2���cî���7���ߢjq��X5s�Ļ��v�Y��CeO>J���)OVD���+}e^`�g��&fK��������u��<�Y����)������1�vnnL����ʙ�,R*w締g�6	����_�&��!��d!�w�6Rv��C}�?r��K�T ��J�Qm�|c�+l��tB'#/��gM��L�]��Xc][s"���&ʝ�bE�U�`Pݔ������R���s�ź,��4����8ξ,�+����N�Y�Ŗ4�Kr�N1T��P���o��H� �ݸaΏ�~��wQE_�qņ� g���Z�;���s��j��ɷ_~.;��(��{��ad��<��6�#gwl� (�1�;sV���:�]�A �"\�&�V�z��ĉb��Q�gL���[9�����=8�U�f8����/H�)��b-�R�yAG}�N����ں|�8�1��8�(�(�  �&�ʹ��?Q�cAgJ}p�G�j��3|x��eF�xB�
���d �mi�-Y�ug֥*= �`��3[{3v�F����m����?���ff�7\ƙ�u\թL�m�<aE`���]�g�����'0V��5����D&��O���6���3�x�"�8�����<���γ�tX�CУ�cyyU�W�demU�N]ױ�.�P��h0���>�� [�?��T�j�*�a��g�����)�M��١Vb�ϲ�~u��fcwm����0M��9���|�m��T#a3vyxru����L�a��ӌ���)[���MD��q��mVŃ"QO��Pg�]і�˺at"N���ڒt�����PQ��3\t3���`��M�UZ�A@��&<5Z*���f�"O���^.���|P�P�.=�a������#���hw[�>�2����Ȩs�G���/�[������p�Á�������2i*��nP����B%����T�����������C:R	�"�����?I˩������������w;�l���7_�;��UM���W�{�s�1�Q��������?~'7^gt�8j�%[A�B���=����T��"����y��������f�A�VX����hYn�4x�y��.{8PqxBѨ��`��l3ӰF����k
]�jhhfU��C�t�5��j�`��?���ΎLu� �,xN1S5�J@�Q ��XM�<F��бv�����	;�/[sy�r����{nE�tn*��@��3�G�z}	�Wu�*�QU3>P�<��;����IpN�A"D���W�D$��@x���Da����8m'���zq��-� �wtD���jZ�?��4�"��V�;�+al���s䁔�$VT��B{Kk����OL5�iG�CfVQo�n-�84x*���B9���}J��y���s�B�57'��&	�_�k��P�Z ��wd=��$w�]�>�L���GR^
�>cv�5'� �7��w\Ԥ�^�&��d"V�M�3������(
Y!�q�HMr�#����q��r�%�A���޶���=?��Q����7�	,��2�P9����<O�ܾE�孷��Y���`�V#9T(��z\fMُ͉
��@
��xΞ��������VgU L.�YU]�Bo���g_ga�4�c�rb>^�z��3Π�?���������skNgr�M@��i� Շ�f�F�2��)	(Fu��$`��l(������ه�˲�4h���<
�1nh�6N��m�ۡC	A��²�=��@����cu<�˺1h��rp�!�����R3����a]b�R�s� ��]r�F���8e�*� ���+ֱ�����h�J��&�Q�M2����w�'�[���Xz�?Ά�rv}EN�/�OE_76j��]�ۚ�������ٳr��kr�r��r��˲�mȶ��3��(	gJ�������I�����_�G76,�E�4�vW��"�v����F�Y�����=~�5�?�E�9WLyL��ڵ�� ��-]t�[O�;���x�B�&����3Kᦳ��G[r�|"O贈�de}M�_� ��\����:R�)�쀈)_n�<�^�K�Ƴ}n�ɔ�����5t6�z�_.5\Ѵ$���pD�{:ؓ��F�c5rq��Á9)�,'}�s�����L��k��\��85%4"0:�U�e�x�0DS�9��W6F�G�O��䠆4ux�j�	�A�ćt+�Ӄ��H	�A�w'g/�����{��i�8�d�oQ(w�I�j��~��4;�{��l>�еr�҇�l��E��d��
�>)�x"��^�RU��G���m���
��g^V��OPV��?��"ϟ��N�Poj�5�u����ހ���"�w[��'��$;��=�"%JW��ܹs<�ь�13Pe�6\Q{:�r��������Ƴm�b�c�`!�>v?^pN��,q�,��C>�oAb�C�_Ooz�oh��R�]R_'�GRq�3ɋN�\B��p���BS))8��ǋ�<�ػ*B��v\(�4��X�8렊�ۤ������@(W %����u�,2&���u:���9���D̈L���Q�^�g9�}��ɂR�w1npʁ"���G��[l�������W��O��{<ۖѝN��UѬ^��`O�v_l�w�Zj�p�rϱR݇=8�!��~�����\�:�-�+�`�zS��B��חE�~�Ś34��t;���@Hss�!�jL���K�2#��8�1jag�1�
'�~�@/��:�(�v椪f�D�`�K���!��l�6`]ΜZ�ٴ�u�g��[m3hOd�M� ��_��SiH&�tP��li
.�PEث�ˢp8�+�NY�P�](v����=�H!�QE)���\(3YQ��5��C����v�|���5:���$3[��e$t�}�����Ԇiu%Rdpt(���?h��cu֑U�X�g����(2Ϊ�W.���"��4 ���� bF`
2�������tjFwkԒ����sa���pN1��7- e��&��YjM1����W����?��.��jբdR�r�ʈ�
0�������TP�������P:�T.�zA~�����;o�B�A�jk���s�zmʏw�ɣ���������<��������;��W��s9w�U�Z��t������lY��� EC��	��S+
��7�{V�FI���FN��v��ַ{��8账��wxT�(t���!���hM,�"ڷ�´{��e���0"�h����v{�ƿw�/;ϷdgK�v7u���٥�}�1:H96KdV�Z�4��耪��h4��:	{q餭뤭�tS�������&��L�m��#=��Y�p��y���^$%�?�>x.?p+M�Ģ�@��=Lew[��]�4B\jZ�,6�az-q�0U���p��y���h0�V(�Ǎ�F5�M��d6�� �~}�6g�nO܈q��u������F�܀%��g�0�E�{E;�C':8�C7��igwC�J���a�A��B����ߥd��!���@���h=M��z[�@@�"��L��RǛɠŲNH_7����~?��JJԉG�T���^ʃ���2;�T���y�Beކ��h��S����F��b�D$.��(�z�m���5�8[�^�9����%��)6�l>ے?|�G���pn�������G���u@#[+�ʣ�-P���3v`�|��YN����`������n�����P
�ښ�PL]�T֩Y��^G=8Y�����NeP�dc+���bc�:k�AD;�����$8[DCgs�^�ƨ��VQ	}.r�"�g̲ԃW���
t/�>�)Ф�J�����z��rp���<����W'��V2�'�9ް.��Y�'�l�&M}��\uu��t�uz}��t� ̨[�G���b�JJ��{f�3�vB�óeQ����#Y�ԥ��5��l
�n���,�����,��t֣��\Rf3+Y��ls���g�E�C� Bx�!5����c���ph�.� #3�X% �QdN9�.�[w�]>C�E�T2������϶Fx���$˶N\�5RP�IrJ�72{nj�fK��?w��XS�mXK��i�m���c][�<�k�+��U�6&�c�<`_4�QB�D	�����{��*.�*��
:)�y���QQ6�C6$o�W:�d��6�!�os,� P��y;��e�f�^׽�wb�T5��N<��J����Bǚ�سk����[o����|���T�b-!Ԝ�e��#(B6��$H٧��TVO�㞂3~����+v��R�X��/�ށd�e���w��s��+�ՙ_��˯�q�p�2�9�b�y�5�z.�;C9�Xs��� ��F�_ӌAZ4�&J��S+c*U3���.%�
E�9�g~w���ģ��ϩ,�����Tl��bmϜ��ѡ��X��V!׹��+�?�'��p��:�CYԥ�T[���$�z�c֕���-���+�V���7_�D����X��t_�������N�f����9���f![��?�t��F̲l�`E/PsP���pLS󣬎���ܽ����50k4�c����� k�F%͡Dz�@z��}�(���	z��e�>����`f���e��Ag��y����h4��{j���Pϩ�т1i�i`�@��SH�&�ҽjۈ6M�7r�gqu����������ʆ${����?�FwM��%��Y�Чf8O��s�z�Vim	�ػ�ѐg�4	�Wm���s2�a��OgcknD�#5�qjp(j��a�Ì�Qd���y���z75�^�&�!�2D�t��z��?��T��gըUt��:M�=�C@�b䔒�SFg�_:�amUQ�*:�pBߚ���̃Ȁ��N�����H��F
�p��#x�ވ¤&�j4�Ǽ��4�mn���Ӳ��h�!y�t�\v!/���}��9U�[�_�?�s��s�8����q4�WQ�h� �;S[3݅��8\/^8%�:FO7�b')��~_�Q̦F� '4 @��2�r!)���W�T��Y3��l�d8�B=ae5���:4�\�T�M}�GO���Ξ�Cѱ��dd4�[�Ɲ�ob���cD����Ej���PD�ԭE���t��"8���#�Ϝ���d��0�ﰦagL+ش�q����@�FZDĀ;b��8*Π�U+���]rs�މ�uP_	�!if�:�4�`f�2.QH�0 ���N���w�G��q��eP���n�E�@:���ς�a�;u��K�1��Ӕk	uL���Q�zVMB:9f?�'O��=���y�0'�Ü;R-��ޭ>��m��զ�U���2�'�!⎠v����*�V�$Jaː	���^h��:�ckp�!����7¦/�����98���,CK�MԮ`0c[����ph`0˭i�D�3U��&M��S:�PN�6�|������sk��k�o���kEwm������������߰(38�@�	� ��uv\��.��վ0�E��/q�x�|Vϝ�Nu&���յZA�1�3&�\5���=�-cY#�b�\:uX���*����@�ܩ�v]h܅5����d�;T���>����8o�1��2�j��cm����hY�67��ﾖ?��?����.W�_�z��:�����;(5;�#�?�尧�=�vh� [�QS�P�O5�L&��I�.2��?B�I1y�C�_z�����*s{�wV��j����頧N��l<����3����ԌY��n�ېv�:�_<�"N��R[��l��HMY]j�|����Uy�x��ݪ���mK:��O�}#��!K�ΰ�n �#n1P�o����<�	u0���OJ�(�� |�Q��_��*e��]��Xx�.�J�DZA�-x���B��S	���_��s@~�O�$6��ߓ���ɞ~���rG�j�u�;j�r�Ԫ,/u�Ӫi�Ԣ�2�������W��a1��+����������DU�><��zG���)�ŉ��՘"��l�FEz8�f+eْ���,��G�Psw�B۞�u��P��Ð��w���F�Ȋ1ia�4MA�����7ߐk7n���
i��7�Ʈsm+H���_��j�1o8���&�>#�e
���b��B����16
�H���e��nhU�2b�$��q`� ��f��d�p�V�9��m0�(���`L��׿�3��'4Ufx��!3�5kA��1�ܸƸ-��%Y_]�3�׹w��	*�K�e��!7N��d�<��8�;*�W��BP�ª)y���H�U/"��ԥ�P�eX�o�;�٧�������6��������x#��'�I*u�0�@>��=����w���>���Z����g�y�����������e��v��ZKs"�T]Ѓ�H+-��62@+p�hF��a�>�[[���?pv�=R��AK:�7b�������3`R���C��Ag�c�"z�z����	/�F�l6!�BR�K�� ي��F�+mlZ֘�;��,�^9�l���Cםw�
���T�@n���t��)Ȱa�ψ��' �6��� �[������萚�uG����L�&䫕YF:���ޛ�d��AZ�`��V��鞜����e�I��*�T�=U)ȗ=�NB������w�|� 6�鬼�Yq�4����V+jx֠�&8��]��j�̱�-$���!#}&#]���K�M�������]�p䑁&�"s��P�hԵ�f����o=~${�k`�������:4@��3�s�:G^ �Cd��$�o�ƜwSf�q�o�Ԭ������f��΋$Xp��� ��=�<�I9�����a��l
UEEã[V�9�-�?��ׂ0��ʪ�!wW��o���g����|l�:2��X���kd�J_����3�9��OQP���"�N�:W�O����.��~�(���W�?���o�~�_~�����Pv��`��v��4f�� �Ϻ6�t��O@���й��ܡ��l����"�'V�^�yE%M��c%�p��s�"/�xZ ��p�;�{�0�q�����˓Ǐ��_���&}�S�-Yj�Թo3�]� ��c�"�+���Ku�GVc��Ǳu�oj@�.��c�r�����n��i������~/I{Q���w�|ꂮ�L��Po���+��_�Za�v�6v��n��n7&���Y~��A�+��	��W���TTT�GќS�C,�)҄�����C��eU�Q6���rﻯdg�t4jZYZ���/�r9vE֗�4:�ȅ�����eT
ĸ]7�4��O�{6I�%�b�3�2KW��bD���.(`F�������'����b�;Z���ݥej�s�ވȜ��ciS]�"Ľ��ݏ�MS���Q�H#Q4����*7����U,gCYEܕ��o�H��׮���hN�O��J���o��IN{p�OiƗ�9�Vb���}��}H=&q�9�4� �*	Kr8n���P������R_Z��T(m��������ji���rnE�;���\m��o��@��Z�6�����D��o��?��uU��`��-8�oF�{�� p �''�^p0��>�ac:+v�Jb�p\��4�4��uP���J&?V|����Y .��B>�X�E��]#{�{��f|�4�)='��o��L9E?��������?+�?��x���ez��J.K;K���5�g jf���k���@��Q�����4 ĵDS�H?�{ֵ�/����s�5�y�F��׿R ��D���Yd��W��߱���� �����H?w�k�ƵKx��n����ۓ�O����!�D}@:�(�P/����� ��@�|[�Z��Ts�AW8�) H`R1���ޮ�e�|BV &��Q_Ϭ�!��MK�T �ʺG%�5�M��R/�u��	
L�?"�K��8V {�wT?���t���E��ǥ U���ٴ�ރ5���h����^�s=@@@L�3y�ЭCS3s�ԁw��$6�d����L��	�1����!��R�E��������`�C�o���{P�h�o^6󃴍d>�����������@c8�#�i@~��)�xJ)3�!r���;�����J���@=0Z	�Eg�}5��P{��H��6X
�BM��b����ￓ���H_�|����y�Gbt)���$m���wG��3�f#���ƃ6�@˵���O$��[��a8_�l������z�]�m?B��.Vb� ~�����l����¿A٬�3�"����m����ͬ��Ŧ�KPH�TM�T��MIU"�Fm-�7��~�c���uYi����k��o4�ؐ:zܚ+e�"���QB\0K$�4�-�d��m���\φ��5}��U
=u��C$Bg�ǰ�� M��������S����'���H�%-1�$��3��*~��B��X�`Wj�W+.5J������8�4��u�u��\��"�/�$M�47��ɔ��H��ut����@Ct_mS��@���y��G� Ui��r��P�-ڸ>�n�f�mr4hfF�L(�?4s��̤ ixA�E�OQhV���<[� U�dZ�5U�`NmE\$THH�gXF��R�|Pfh�R1�#TR�����_~`�p]�z{��w��k�r���[����ŧ7S���Q|��F ��� 
�����ƪl�/I0�TiD���tusE��y��7�!����1� ��l�!'A�"$pY�=(^.o���i�b����t�yeR��R.
RS2�.���$�M�H۵�s#7V#ɥ��\�,W��R��f�U8}b���F/�&E�m�d�S�*��th`
�5�3�XI܌�>���ע���A`�oY`�ʨ���7�w�,�"��DF�`�^���*�RV ����OI�y����a���%�	���M�0<��` T1J�(���B/d�aÅ�r�1��g{�U*�!PX�����b�PXG.���HM�9�D2#��\������* 5k�y����y2��.��8&}d�T#4K�Y��=�iw(�V�蠦������Zl�@FjI x���AF����ހ���jX���뭖ܹuC<x@p[Tu������=�����+�R�� (�W��|�upt|fSC�� 3��f�	<SY��ڕY�4yMpX�j!�5�rn����T���{����ဥ]�jJSN@��Y[c0��ٸ����D^��7��45��;G�܇l�ו�u$�l�ı�����,��kH'e(�
l_�.�IL�R��~]���ԫF���O�*f�G��� .�S�qZ��~��4��olt��G����9H�Mt�������M�t�}D>xů��&���.������?���mZ���WrZ��>���b�x����I��C���F��η+U$UM)W�RU+��GogS#[�=�����?}hYnP�J&0Pr� ]O�׏�q�m�5wik[>�{W����=�}Gm~P�f�Κ�6R���5ܤ\�sZ
�>��K���_�;��	�,�	���	+:a�{�l���^�����Ha�Kj}q<ߋ���b`�����Tʩu"i�M;j�{��������Uʕ��������99L��۷o۠2�F�g��Q��hB�M:�K5��֒��p�]���S�SC5o��{�$7/�ȥKW}"?��H�<y"��^����=jJ�җ��b`�5��P�XgE��WA��aVÁ��$�6��VUJ3B�#��`E:4��t.V��{��~r*~~ox ��8"p�,����M�wM�o��sy�3$O�d��Z�.k�5Y]n�͝ia�i2!_]i������ܐ���N	���iɰ*�����+r�������G'r����hW/z2ue8�ʷ���/�����yFԊ$e"Ђx\sJ�B	�VT�	LFR�hV.d5?��r
r�g��ȗ9��B.f&����I�J����2�PA8�h���ݗ�����*xo7ʲ�iȭ����o˵K�`���Y���-1�`�U��Md�Թ�\Z�֍�P�z�P���#��ۍ�<����|+{o_( ����}_UƉe�3%p~�<��g��[�i>�'+�:�/�L9Q/f&�w�i��3"`5̠�����#5�-�A޹rU�4�Ѿ8]�5d��#˞Q��9;6��yaT9��-Pf�QF3��&�f�o��P�*O��7�YFJ�#ov�W�^\S�,���kɫ��3�כl��U/hL�%�0���ޟ~�@���X�_�o�t<|?2�O6���옯+a��l��X>�Mo ��;wA^�}�LW�|��L�|��2Mi��<>Mi`ܺ�Q <��.b� ���<�
��O?�,ti�������/w�{�����O������jkcIn\۔��Q_-�}]����� (�W�8_�zY�\�����?<��ϞH�ߣTװ�g0}xT�P]��Z[�O�ޑ[7�ș:�'�~��k׮����޿/_OrisM:j�O��e_���kP�w��2�a�;�.���&4�w������ާC�o��V=����Vd�J����)�xCu�o_����#h
���	�;�t:��]�l���B���,��Ϝ�R���taP�jPqx������^�~�,q� ��:�mEڝ+ hD��hwF�*9�K�-z��`�jjO��\V��jR����鑌u�0Y��!��$��g���8Mt���-�nT/N�vt����퍢=�ۓ�_L,ڝŽ7_e����V���q��8�q|�K৩5�U3��1G���y����3L^�~-����n��5j
(K����.%ּ����=�R��S�w�N&P	"U2fe{g��k��*��I���E����J�?�O�(�n�ʀ-(u6UC���~M�Lt1#,d�0�[SpN��U��*��=�>�v�{���"�*�G�d�!�d��7~�)8�/5�cR�� ����~~h��GF�6��T5�����T��B#��?�*y%:-q��0��{��Q��'&�����c������R�``�;#�n�	�3R�� q���F�5q�<#?4�JFC&>o���Wq}�M�n�E�B��|(/��CAɭ���0�4����)әli�x���@���X��������nH�^���/��ߑ�6	��&@���ʒK^�`�Z���..(��ڐ��˂ai�ǧ,�*�7y���N|����|�fC|�;����S��r|ڗ�L�M��u�8A���t���c�����x��0�^�^���-�/� ���I6��<Ƈץ����X���{E����v64�Q����;r��w��ϮF�}��,�j,wC�8*%�TX.[���L�������Tu����x�����#=Vd�����Wu�z��DUi�mua:$TjP���fƅ�R��$5%�\� h��u҂�1#$����^�"?������)3^����&�[;��"�6B�j#͑]�(@��p%+S��@�������:(��͵��^r��2�s� <���e@f�/@s��Kn�;���Nϗ��[2UH{���].��NOt�#�����N�x�1���)�C�w{^��UE R�,�_���G/ ��#, �퇹D`��l<�S�O�3v��6���x�����$>�t�7�˴����!�>���s�:�/���d..��(0_`�6Yȋ�3�ï�
V�=j�ٓ��L�4@V	8����XnSj�;�5�m��f_A��?�({��Ȩ�~VJe��5���K������7_�E���[����4p�h�0�H�{�y�_��w$/�����MM.EʡL�403�U��4��֦,�y���{CG[,[N�K�E���
pC������.�i<��2ԣ!��#��铒��#}��7�����x����뺶�߼%u�k����ta��>� �Ss+�<�Q����#�H5�Z����W��&��)�>��EU?��[T5��P�3�e_����Tz�&FL�z<f�b��RWm*J���d:G���[�Pn�y��,*�'ٶJ-E��x$�u��3�0��0$����u/0� �B�+��y`�����֟k���-2�c7��E}[X7 ���H�����:8Q �Q���D뼯�ˤ���VMG��L`�ސ��ST��5�7�B�S�lhl)�������e\�7np���`kA���t���\�dz:͵�I�r:�bu�_+�>1x�lt��Y��U��W�U�9=$v�3�f�9��@�r���K��g��a��F	��0s<[�D�|��1T=�G_ڋ��7�'��M�[�#17���~�����\*e��hd�-�f ���8La
,��������_�?d�h���3S(:
)��<M�N&���}bM�����է�7M��#?�W��$�eٞy�{��>h��C�����Ӄ=Vn�/v6�r]A��>�'����t�5h��t��0��<�Ȃ�j�*�P���&	վV�rI�bK}����Hj�f���Np���wOd��ޓM�۪4�5C����Y�����I����J���Y����A��E�E`ɉ��R��	ȏm~��~�w8K�<Iy���1̧Ǉ�����^[�V5Ш�&7�^�;���i��Af��S���s50j��QoQbQ2f�ӊ���BQ>qYAĒ^�:�S�.k.#a <�ϟ�c�c�������)�0�Vn�K�_�\)Im��7s�q��79Y���L,S�X4)��z(4�q.1�nY8o�"6�a����\���چ.���B���ۦ�Z����ƌ{�i��a72
��m��3���	�Z���g��x��%E)7�y���ۯ�E _���W�.�<Z"�;���|�߫���������\<����}|_��|a��e^��'���WAb̨�@5%*4�z?������.ӽ���6��;)h�&V��*X��+k�Q��7�(�(���y��S���IC/H�Vg�ߋ	{����$V��ݬ�a�=V6&��%�&���?#�8#�Gz�*�\S ��֤�{fucK�j� �WuOoa�����\e��Wb�$2!�)�s�j�ИY7R\�����<�>u+�i*�{��፥��s{c]�
hAI������xL���n�ilY��:�;"�R�r�Y�f~���кxf�t:ss��L�v)�Y2�hJ䘋5,���$�7���78?9��c�E�A9>L��S��	Uؤ�\Z��ܼy�kM�x�+#p�L��~!����<@�r���7�.�����1��qd}d���)����e�!�{�σ>5U���+�j졛;��t���}L��:iT�����2�D���i�Sz9�G���Q��I��Y�=���]�BIfG�L��A���pЦ���+Ib�����s^b�R����I���_>x@j���g,��uL����T����=��𓜪�D�	�^X�&]�X��h�jM���hh@u�Ǝ��w`�s4�,(��.--X����*̫���s�.�<f���H��d��M�ũ޴o�Rv�	&3�i�{�[�ҕ�[��,&�J.@��f	��5�b_�������sjihÃ^����>���;N\M�U�$�QPdէ�\�AF��a��윯�s��t���O@�R��� [@�3U�
�q�"H����vLX���)o��9NLIJ� h�G_�/?���
$ɒ�~G!��^i�_g&y���ĄL�%l��;ˡ�o��c{��AAnY:�c.o�����������8�p���b�AW��21pZ%��'>dk�^/�dj�l}�]��*�8fQ#]����{t �4�h6:r��=�^�jG#�M��$u��a,Q����/	q�޶�Ϧ�t������?rDt��R��jpBC4C���\��G��.�醇.����3��J*v���>�ς�Ʌ:�����l��Rez'�H\��!]���D���QO�N�Ը��U� �ԙ�xx}dJ�i���z���+gÀ^	��j �jT��i��t ?=|*�ޢ���N�/����SF�g]7`$� 27�棘Rg����9$I|�&�͂.h����cSjg�!�)�̮y�are����0A�K�|G��敫�cj������E�:#����+
�P�蠧 Y�0p�Ø���%��q�Й�v ��R�Di<5����{��(�ɔ�Y�6��n�	�Qd=h������Ůy��a'N�\mc��c;6��֭ `�c �y��r�� ��T\3e��</u�Kk١�l�I���TKй��r�D�w�{�Bmu6�A
'R�k�c�"������[Ja9>05 K���um���%c7m��:�1���]� ��>F��#PA[c�g�D[_[�N�Lz��I,�����$U}_�Ӓ'��S+���4H�o�d�ǳ�ّ+7�I��D _��O��kx"ic]J��\�s+C��s��ځ�Prj�g��tA��\ ��JIA��iO�G�͜W/_!ȭ@�O�Yi\�Iu"��A���,���_��㩲�/��=$`�N;@��� 1q�6�@�0*�����"p��k��c�T�['֠j�Up�VK��x�=�v�j������=\�Q����`J4�rPB3�s��oZ���P�d�\�N�-*Lq;����O�߿�+�(����w�li���>� ��g���S=+C�fҼ�j6�D.|9d���h�[�J�a�vR#B** ��i���-�c���O���C�3�=)<Xu� �UM9�f?p���]tet��k�F�Ф�g��"u�/�����̆!p��*N�R�aJ���\n>
�DTO�Z���o��m>-l��yŀG_�$�'�2�a�_��'j�sS�ѐ��q���l��T���ˑg��~@E(�s���5��1���5E��]�����1bMP� TԀK$�2�_���:���yW�ㅜ���Y��`_>��=�@�E��l�R\F۬�S�	�Ĳ�7�����̨�9XϦ�b=�����')TU�����WnbP^rkrj��rكX4�}�/�OP�H�D�Lm���4P������߲����� ����Z�n=�V�9P{�����V_"�{6�ѮܺqS6�V0�B}IY�3���2Q{)j�#PNГ�:�ͫ`}N�):1LB��IЗ��C�_c�r�*8c�ҭi$�)�ji�>�[�2�M�I���2�~�.۞X��vU��%�Aϛ�_�lٜF-痔�{���s�vnm�)˕@������c�w����
��2�ˣ�Ln 4�RU�?I��]�R8�k�nԪ�׵<�����C�ؿsS��D�_���L��^}T^ߪ�]� �U���O�[2���mB��Im&�xh߮J��S��@�T��x0*�f�2�+1�q��p�gw�T�b)��f�|Ӽ�a�I��3t��Q�u�C9a��ky���PFF�5��ݾ)Wv��D6�E��t���E ��;ɱ^�u��L��Ŋ�D���}Y�+������|~v��e���<}�N�O�YX6���'�����\n�)�?������{wiN�$,2q^th���ɦ#ɇ�,8r�+�F�ְ8�YQ5#�KjI;zȾ��uf��}��
�Q})��nu�þ�u��(�TʦtA�Bbǂ��Оg	o<ɾ;�H�u�����2���~��J�L&�}�w_F�;��+G�!Orn0@��$���!!鵇��<n}-��^�JMr�D��eq8��&]�Y���`�K�G*��Q���q�,�\EƲA�~�aB���W5�;7���e�kh
��4�ω�&G��d���8͹����ꔂ;4� 8�_�x]���@f(�îL'f_ˋgOx&��5A�B>�G���J�h��%�( �6XM�r:ݨ2���Þ�G5��I"�j0���NM�eS�PY
���.��A�Z�Xv��S0 ��: *iO>b��������c�۲��FӴ?p�����r�`2ҿOz:�W.KK?M� �ȸ��gU��M�}�Z�I�	Ȼ����6c�� �}I����2l�Z�7�|�8:؆��í�6�F�{t|!�,�Άlol8�׼;ܗ��`<���_Zc/>M��͖3;���f�lwؓ��ܷ�3���;ާ:պ�����+�ry��У����5j͗�,q)T'��U��Ō[V�(��n
:�bk ݪ��V�����M@�#e���8�m�9t�L���q�ׄ�6!{���hX�̞��[E�}������*����huA�dyX�߲�A���eP�Ѓq�͖��qj=	~8�}�d�.o3"r�ܤ�B��]j�r%�f9�ղ���~L��B1f5��ѫ�
�L 
�� 48TX�u�	�U<4,bO�Q��>0h�2eV������� 븞�1��:�~����Ln�D���L�KzU^>�L�PB1���	5�r���5�O��̽�����ȜO.�6�����3�eXsK-��S����{���>y�uZ/$����AMR��R��/J���(p�Aw��X��D}{[v����o��կM�e�Zb���5�P���h�����T}$k��WV��� {N�wq�Y��������IO��dKlTPS�T9D�胸��%̆�A[����4�0��䨻���%KYᗼ龂D�����wr��V�aݯ7.o����̍V]�R��#3���̄��V��(�[b����9�W�B����t4P;��"�?���"���w�w;.�B�hoWήʥ+c	�7�.��l1�/��'u�Rk�[ki�u\Xg�sA��H�A����u�a��Ғ�zX��`�/t-	L�������X޼z�����b�	��t:��2�8dI�OH�y�BRˮW|ee���N{� wo�XNu��vcˮ�:�TD8��c
+���cܸ1��h[�rC�+�F�|��e���uB[)p�l9�(�Yr����O�&4��.�5�M������͛����KI=f��%$�˥-���W�N�^CH A:)4og�W��D5\GH�y ��C��HKY4d��9+{/4��gFa)����ψ�Q�5���w�ж�,�yM zpA����t��]�r��%��Ɏƥ�H�� /F�'%�e�ݽ�k��p�s�\�L�5�I���L��7��C����LQA�L��Hk�Nf
�Ba��f�ǲDm����a�d���I��53��8%U�)�kd�|��rOA *>�b��׭�`�;���AO������y�C�������b޷�'r~��zU����$�yˮ�F;�2�f4�BU&tt4N����:ȷ�~+o՞�ｓ���9ɝ�>��ͽϿ�~,9m��mN�5Mm�.���Q����y��5���u��#ꏨxC������7����:�޽w36Oc�W�^4�V@'Ӂ����ʺ,����8�s�7�������Φ:a>�+���G��o��㓞��`jskU�/o�J��kY߳}��4t��V����O�k�P�sG�/]Rpu]�zo��&��o��V���gʝ�5���\��]�ّ�� ���n�u	>iɺ�3�>`5�U�ۡɾLp�ҩ�����9��L�c;��v%�7���M��/ I<c��i�
^Z�f��㵘Bi�Y��}�!d�}ń�n�a����L��S)l�j u؃�)�X���g�F���($S�!Bf;"f���[� s�r�4Hu�>e%�e�B��4�҃ԣ���Az�fjӑj�jฤ~��@���;�T H�e�0��g�-5Z*/h��v���`�	�V�T��7p? ��z�Ua���pn��>�4]TM��ʅ,{�X*2���]�����鞷_\_�����"Ug���6�1f�,2���opE����[h�����X��fmT��`\�3,�3�J���.�gl��I)�)��=�囿����K
 1�}W��5��58/s.P���`ޚF�c��F�05:�rd驜2�Z*9F��2�k[�E�Є�� ױھA���]W���Ej�8�};�OX�Ŗ���Q
z؈&V�S�Y��J�� [5�_����
�O䳏�K[7	��_�,�+���*��a$hw��!���O&��q.��ĺ�����U�u1��!�N��Pl��=pC��ە�^_�z0�)���&ķ�:�.��cO����{Gw.����'�+[�i~���\�b�	�<[��g 72I$xN���΂���#���l�/�.l��Д+3�.B��|x��b��g=<���)p8 ��10ɮ�e;Рnus�%q�f�QO�c�D�v4����S㭓�?˯:�>P\�%j4�e�����H�Z��0���4bp���f/��LU`�&���Ѭ٦�u��
P�����࣪:qS��X[�,�R�:�q�w�>A%@�/2�6��U�RZ>���8�>��>���뽣�ư�[,��b��8���=u��L׾���ߵAݨ��	|��zC�k�ϗ�Y�Fs�+#��y��D�f\�l�Z��URkV1ʕ�c��	�n�2�be6Ä�����4�����S�#CB�ᛁ�4M�o2��iV�WH����I,x��CH���t�A݊�B�L3׷�����x4�Rd�`C��
ơWYr��<2(�|c�a=c[O�3����l�<;�2��,TMY߾�i��<g��S~�q1��JV����o�o�@*��8h˷��Th���:F	3����eK�YPElܽэ��%$�n_�J{p�� A!��;�񙮝󥪴�UY����@y���t
[
ܣj,u�����ږ�mlJ{eEV�ߺ�h����^�����N���BV66Xa6�\��ԫW���~��7��o�����
 m�!]�)�- � �%8\f�=�*$4�V���s�l4��'�-�l'^S�*��nhM�ޡp�o��X�k���u�,-lV�=�ߛ���`�k�WwMJ������L��B�����&�=Ώ�ڗR�5o�ϥ"��aZz|)���ڎ?2�$.$ 7੐�<�UH/IsJ�Β��c�X���>��k��[o_�"�}{[m����c��v��br�8�#�)�����kH�"A�k�$	h*,�~����R ������m��>]�����c;���"~��u��ec����c��fr���b������ � ���$�Z6�ɺ��y���UR����.�F�U��g[�b�e���
3��݋��{������!�5�k,6.e������1�\?U^�p�ء�ݏ�̾�^g�v����N���c9;ڗ�/�)��� �kn������vuM6w�Ȇ��j�m4�R���	�$B���'F��s�L��g=���P�A���\�^�ˊ�P�P?6��MT;׬�:���_��W�/wVhC��-먨*��3�nW���4�4��&�zO�]�$/�>��gB�sTF}9�8�=֕��V6q8q�=��J�a@Q贜� �o�4MȂ�7�=E��n^�"����-v�{vP�e(ؿ%��*�5m��m)`GJ�� M�b�"3�0	M�l���A�b~>$ �YG��I��Q-5��=E&��Z�)eD�uk�Cƾ�K`�f%h~�=�ZwN��%|���i�F���)���z1�#x���g�4Zm��/K{m]aŴp�]D�(,'�n�������4h7�-�\��+��k��+G��2�n��Y[Y�FAa>��|��Aa$6�ջr�d�8����h�g1��ב3L��E~��]q1�O1W/�ʫ��9> 1�h2�Lj��|�{�<dz�o߼�2(yf���S7%�ٹ�JAv|n/�H�ƭ� '@������N���X������bR�����н��@��Bs��� ��5�.z7|@�c�: �:�^�J�ԿC��\��q�,�+���"c��t�{I]_�W�1�A.URk�eV�Z_�B���ߏ�2�w�i?9='��t��cS\*J�e e�Z�C?��u��&_~�%�����Mk\�ʕ+r���vV�f}mMV7��{=��%�D2*3��B�"��i7 M{e0쩍�P�zC�������:�.ߧ%��VdTeY�k�u�F}��4��W�˾��\���ͻ�e�����Ds[�d-�\ږ�z.�g?�=�ӡr��k6gù����6"I�a[8���^3�Ƀ�؀���)>�����^P5 ������ĕ��tZMR*�N%tkS������*��(���(��8��8��Z�0[o`>H���j���<��b"�m�[�J����l�i@�jk���͠�lR�Α݅-G"
A;zPi[�,F^-��Q���TS>Y��ڃu������{f�!v��B&���|���[�u)���gG8���@��"���8 ���R;��H�+l�ޛ7T@�kKe�
��>7�bF�jS���STLG8&=��A.@5a��5�Ǡ"�ﰾo� �`g4��[���(K�J���{�lZv<3�{���2�^��S�|�{�U���Eп�Db��'��ADQ��X(R{j��1_V�����/�AW���o�ח�H��g�����R�C�nI�zMFT��Q�YT����VE�@�j��zG�@KF{��5���2�L
�lTҲ��z�=�-�E�\��0R�w�,"�U�5���c9�}%�~�Q����`O1|߈��1�z�%+����ͻr��ٺ��]�#��3�ۆ�'��Qfc�U݌q��"օ��������>�Ͱw��e��ܪ�`��w�`�c�`M���q�1<?�������0p1������ڕ�JG��W���}Mjg�����y�LN�O����LU�����m @��$��	�CCX��4ϣrW�LM��O�2��`�A��>�c#@� e98X6�����]�Ԝ�I��j(rt�'=�~�$���LG�m�O\�ܤ�+��,(��K����n'&��7՘Ŧ}��VN��E�ְa9����g̮nlR#uT�'���/�u�J  ��IDAT��/��|Aп��"���r��ǲ�}�Q�p8"_�Ԛ$6�#r�ؒ�� ��jK�,6JsK��X.ѹ���w���p�e����lU�l�o��dce�(���@�g8ܪ��mѐ�5-�� @�X��Z���b�َ9%�9��a���,h���}�����ك7���������@SaMɲZE��Y�({��u����%p��M��ӵ��W��@�ƍ�
F/sJ.L˭���P�L�Kr��O��Gwd�aY/d�0��ٳgrp|��!u4Li���[��`F�c5Vp���BOY;�I`}���_�j�֪&�
�1�� d��@a�R]�h�f��d0�����D��/@��)ȚA������f�Ne(d��4GPH��d�*��r�A7�2�ݻæ9�n�в���<}*#�N� ���Ә&.8��Jp���9U�$�����#��o䛹�p �l���R�~���A��7�驖p}t]uծ�ƴؗ��M�Lf�l��V��I���P�����=5�T�{��,�
�Ȥ���x�Uw�}�ί�L^d���m�;a}c=!;:�2�Mu������u��R�^wU+Ӝ��"��Zx�I�~��&��?f�u �ڊ�����^�ϭ�+&CG:]�j�4ӎ6j�S9�ߙ�ڂ��aA�z��������)����#�'l����т�]�A�	��Q�1���;0[ ���׻���uu���ukkM��?��b��2��N���r(����P�}�ԓ�3f�z]��q�o�6�;�k�M���8]�?���J�@��T��W�b&�޼h�:��!U�W"��F_�h\>�u���5t���v�c�NM���Nՙ �#PF����;��zT�̯˲Osu�b�Z\R�V�Y�w�3W��9j��-`���(�+E_S�G��8�����b����"����,�+>����o�z�RմRS�޸*�����ɭ;w���?�/��?MP�AN�f���R`n�����N����|t뺬u��F���H1l���}��:a��X������=�5uc���6f3!\z8�Ѱ��f���	̔���b"���|�J�,����x����l�!�z]}�h�L��{����`ު\���b�������V�D��)�6M��=Տ�����l�.˵�[�^n�� \�$n-��&����r%Ky�%��(��Ql@�������GO���������U�ru[~|R���%K��GgS��.@+��"���Ii\�;��H~N���&+őK4��]�.��ks%��q&-˅M�1�0pe�5�ߣ���0ٔ�j�Ʀ������L�M����C�%��&M�D��Ȧ?B��j���hs��t2�|�1{X��޳�L��� <wq�W����&{�f��������Y�^���~o$Fy��]Y���HseC��j�x(���{�:�9����&e�0�U�Z�2��@ �8C�2��k�mi6*V�F#R�8�
NF��Fa�YC�W�����8KF3�T��R�R?��4r��4& m��g*��t�3*�DN����,QČ$�5l	����6��<N*-�����#F3E�#U5���I���cw��Qt{�X�X|���rJ*�M;�[���O���[��,� F׵�ui��A�	�_}񅬴;`���ƚl*0���筏ns"��۷hl�~����G�������Y6	��՘��{�Nz�0Խ�]teuu�eE�c��ea���$]��5��3;�Y��� /���y��@4�S�'+H�n���!N� 8�(�;�[���o��}���r���^�KE�?��k���i�1�2&�����߼y'�����C5�����W��"��5 E�dS��T/���p��)T�Á���*�P������rŚ'�iX� �ә�����
&�j 0��v�������{G@���)U�\���m6c8� �*�����4&+	�:'6�b��
���9�)HW*pC�E*L�m�jlRƾG�;8�S6&۾�%�� ���PǄ�h���9�%E1��f����$�<^?�M��阝- w�� ���-�➮EZ��y��h�֑W/_[�A� �84�!���^7���5��~!Q��84O뱌�������>��tG��W\�&r��Q�������.�[����{��	H0_��d��[�,���9�b��S�I=o���^~
�m�m@�Y�*��t�?A*��E_v߾�s��A������R�XA<z���n�d@���ի�R�?~�M}��K�`8�ޛ%nf�l�"G�;u�g��|��2��&i��W�NxAզ����>�����X�������{�}ɴ�C"������kׯk�ؖ��cy�n_^)�u	�r�[Y_	�;�9A�|p�{���U�%Α��]���*��5(������E@Ǫ�O�%�(���'ΰ�+bSϣ̟N=��i��7�=V`����O�dפּ����X������R�(P/[�հ����o�ToK��!�����T���{��tT��n����Sͪ蚯J=Z�`�XG����}#$����D\Pq�-΂�,Z+��%���~@M�������~�Anܺ�{}]v.�HK�6�CMp���Ӯ�=8Z��V퓥���j̦�.���m
?�5�%�H�A@��	�Cf_���ߗI-�{�����rq
f/�lp(�sҁ��S������D�Q�<:Z���̆������4=9yҚa�Ӫ-JRt�2/ k�9���q�}޸�ߴ(�i�h~l_4J@����Ky������L��㈕����}$G���{���K,EW��W'Y�i�hx����슆D�ƪ"0z8�*e���5�B�ՙ--U9�#�9�6���e$GY��S,<O���ؤ�7���\f�p?�g܊F��n����}�5E�M��F��ǅ��o�2�������#:�:�����4���#�Gh��kb!,q���y��.�]�8\6m�Q��w��:� �<���Թ=���� ���+2��S9U�����������_�q���F�痟ܗ׿>Qpܓ��ޑ��>{�w[���r��h�=c�%p�T�0{g
����
�_h�	��I�����j̸vO���Y���f����Y�����'�\DI�?�Ս���*�x������<��1�HT5i>���p�ЎP���?�,=5�:�>���J����~�g/^3�#�[���A����
��!{`��e�e�J�z�;p}P�@�߿`cW]��������(OUi���~�q�ih���^������m�(c ��l賾�,/_����v���T6�.�O @��.J�̈볭A<u�u��i�wW�]&X�G�룇9���{����k�\`b,��"�$u3,����$��k*��mbS3��"��d�yX�fH�B��Y�W\#mH����T'(!8E%qz��Υ̺C�6͓���]�9����&�����T��vL�����;2�;;[�д����N���a�+��ǰiV������h��Z7���S����ݹ��z�*wv�,�)NU�"�4(%ә�G7J����}�^���
���j���.�4�"�� 6I�IR!F�>Ʉ��C�:�f�������#�P|������7�� 2Ooɔ����.��M.mfԛ��v��)-��be���9*\�g,rыԥ�b���b�޿�H�,��,f���3�4g_�YG��ěrQM���?���C�������7��P�H)˨�W�z6�V��������e�	�I�+�ZTs���A�T���k�31���i?��^�����B���A��g��8͹�S�<�,�-�y@F���န �(5*!T�0���y�H`�1�}q1�`�P�̊,i�І����犓�D`F�9�
��������됶�L���9���z>����!�E|����ǣ����Zn��w?~�
 �@����#M�$��??�ޞ~}����HF�K�uA���4�d�oShl�4f�T+N�h�@����Y��$[�9��J��9��^��Z��)s�L<�5�H�A�O�L ��27�=hj�β�ϡ�+��V��x�K��1Ցه��6"��Je5������p�$�(�W�w��M���xSj������d e�\��k bvJ�9V�4�D���Rs�B)�9�!�`L���v'�C��P����J�.��\�zIV�����Jd ��^��eT�`���2- J��jY4׬�[�H���9�>S�Hm)>�"��9�?����SX�� -"
�h�����h
�qAv\�̆�@�:��_�r}b��3��Y�T�m����Y�&Y)y�d���2(Gl���Bc'�����C�ӿ�Wy��ܺy]��A���Vju9�u�����tD ���
Ħ�s���A���-f�~x�����_�+׮ʝ��zj�=Pn�}��ڑ��V����`� ��Gr1|"���d�����&���e������0����࠯\��߳� �"�����5eP�-(hMuO��5��ԓ�j�{pw#7a����5�N���{=qY�Ӂ%='��7��4'3�eu��, �C���X�A�j��0Uc���ɵ�(���� �=�Luχ���7�L� ߯���s648�c�#�B
���LO���Uv�u�t8y���]U[�N��Ʊ�k���J�����(���Mp��N�X�XT�PuDu}�����3c��ָB0��M-k�L�Ub-��pP�ܹq�NPfɚ͗�jM�l�d�#�����ǘ�L��90k��G�cgớ
��o>�Z�p>�c��S� <x��PYq@	?_�Vq~f� {���[���\l5k��pA�8>9�{}�?�se��,:h'���'6U��6��MT�P�i�Tê����n<p,��멋,a�6�I�ߥ]��1 ��J���~!"��=P��l$*k�FG>�z�\#k�T.��e�������|j:1�U��|�������XU�qE}��יt-�>l�� �[/���T��,����AB��5��k��7!x�� ���!N@`�gx;�}S����N��x��f1���N�^_����餞�K]w�ԃ��(����C�������>f����$66d���y��i�{�lݣ}�s�60�6
ؔYv�.%�¹&����;Jl��v�Ie�P���Bm�oϺ#��}�_3��!� ���� _�ڰ�$��=Ԩ`c�?{�odz�tB;ϣ��g�j�_��}[mp+���Pm]X��6Hs�aϒ1o��GC��6W���xO���{��/�]�5��D����d�;37qU���=*KS��`����r�W����a�0�i{��������e��l>�0�`�	˅�_��8ʂu-gcu"K���������tt%4�.Ƭ�%�@F`�XI ������NؑO�Zf��L��Tz��jH�'3B�M �1`#���å�_}��xz=h�Pj�0"6z�n{n�	ڨj1�����[�駿�ϔg��3ڍ!�&trQ��]��8:��h��j�t��hc��?3�����,?�6��;���{�҈u��t�p:6A4ed�Y��Pom�H���3�2�h�:G���J�ҡ76��3E��o�*f�A�Б��0�Y���.f8��}���%)J=z#Z������N�s噍w�y0��Pz�2W�R�����]����IvdMd�Ad�LV��X�r�edD��q����z�ED���Ȑ.��tLѤs&ϟ<�7/^ ��1�s��YU�����)�/�_���v߽����Z4��?�YR��o,�gM>�w�����C�{YnA`|V<I�ם���X�Q8`�m*m`; �*�J��~��ۆ�ϵA�?PUX�	����z�����W@1��00�p����M]vIS�HCz8pe�$�f�xJ���vmͱ���". ZcW��:z�2);'G���~A����qL5�4)MP�DU"��t�Ը��L�ٳĀ�l�Zl;�ɅL)���"��!{���[9����`�Roe{��b}
h�>~��[[[!�
��Rg'����}{�>?�uO�~�	�+$��i=��`_�7�:a��e݌�Ўj
2U6���5|f��]k �'��?��C�bV-k!�1�l�6z=���V��J�<�� ��=?����7q2¤?�`��p��庳[��+�<��t3;�s�gl��"�:W��,{����Sn1�� ���[8N �L
U����l������ =���ae��o��xt�A���͟�;PMa���ס(�۰�^�M]	��e�v��n���@�5E�p�'#N�d�[}p<��7��}G��w�V�}���o��)Vi}�������@D��oj��=��\F=N~�@��_����9���*�m�Q� ^����F���&�2Mѷ�n�U�ܿ_�)�ˣ'��H�����CA���<H�E L��
)����F�3�6��R�VC�;m�_j)����A���wjc�*P;�&Wf�mb4Al`�Pد	�Esf36�2=^�
l[�獛�dpr ��K��-}	Lvk����m���&m^��g83y��k�QfE�80�l��*�%7O���z�5~[���}؇u'RY� ȅZ@5���K�N�9<�+l���sH��l_�~x���`
.�8��(͒���������'-KvM��[PF� �oVm��:�|#�cb��Z��x�L��z$V)�#�m��&�9��lJ".&���{.cF���0� ��(�ixбN�K��1Ȳ�b#r-����&��cs�1%��|��Щ�=0�f+� ĳ!�6X�U�&�k�r�щn��,U���`<��|�c�QeP�i��&� � �]��!u�P%5�P:Id�S]�Q[6��e5��rikYeq�6��È� g�i9����μ4Y~R9H�5�}��g�=���K���~Z`q��"�����zC��Tl����y�|:�#=�ʆ�9 ﵍�,�&G���ސ��(G�Ȁ+��_�KKn꛸���3��yZ��*Q`s�-�k��!U�����h�	�/ OW�/I��p�����$�j�( :���k�����ɝ[�y�?R��VV��E\r���<T�u�����K �~���?{�����ʮ��۟�.�ږ�<�^0{���Z��珟2���&�h	=adP%fu���[�����Y9��7/ɥ[wɳ�ZmH�����\���'�P�" �s�:AI\)W\����%����;j��zN���r73W�
݈n�n�/�p;��(t�;��^��ϰ
�@V;3���_�G	u��/gQ��#f��}�/�]��D
��P���ɍ�{��[kh��f �\�R�5����9�\8���s�H�]�q]._��,�D&�~��Vl@�9����l(�4Xc�l<�u}
���yk����	�	�Y��^̢��e���^���ԇfA/v�aV���&� z)'�
s䁾��������8�H�@�>��?@P���x�W�Ն>2�G�*�
��eR��=�"�F�@��7���%)�l��<��H���72x8o(J�/]��$��E0-�r�R�xz�{����م���hA��9�x��-BbPߐ C��~�mP!��gCZ�/��K��K�r|��T��:���̏��h����k_Y�u	 ����{��}1��n��,ux)�D�uSֈm�q�i����3��#�'���"m�H�Y���Mp����+~���E�"-���+�,~����"L��J:%tk\w�zY����f���/_�����*+p����0w�pX�J�� �d�C�gM�&�S�'RR[q4�g�I���9�kH|%�������|�t������ھ��g. ����S�cŨzB�vyU�5i�nKC�iXk��y�մ���@�}�U�1�2�ӌ��Qiؐ0L�^Y�h��6B4�P��5V�{b2�T.�5�P.�JN>�&��FE���zpL	,��եK�u'���c9;���Z��(|?`8qUL̚p���5�=޺0���J�?���1��)��5:>'.&� <����a�����MiJ� ���dNl�n44�	m���w y�\G�_�	����ύ� C�Q)�dc<6~��Tqc�qcG�t�Of~�̘Ƅ��R#�o>�e�p*oJ�i�n����&��3��RgC�.]�JkYzC4��^X	S`��>#R��G#
��¨4u#��.�Q]�Eۄ2��gC1�\����3�%?�PQ�%X̒g��L��偹�{j�W�����F�� P�6���l��	��;Ů�"]'u��,���F?l�+Z �`S_t�b�He�B�(<���+MV�����h�t`�%�M�t����[�2�}[����z�Y�G@�T���ӊ�
���~�{6=|�X���?���\�qӆ�8GB��;v�_}=�(D׮�`y���w���CE���f0��p�T�K�iYNN�2b��4S��[��r[��Y�r�  ��^�@լs�$3��7�������=���tT�`�A?Jf�s���$J9��j��\S\��.���m���Q�e�C�@�S}�pr����P{���"���G�)��S�qB��`����C9�Nd���L��Ё�4�
|h�y�f_FQ�����{�}��u��?��Xv��puPq�P\5N��AD_����J�՚^�O?��A�������+���J �}����:miU�TI�Z������j�:�
� _���sf���0+Gyj�5��ע�<@Ï�m̤%V��Ѧ�%3�l�/��4k0r|r��&YUp�����5�Cr�eB߅*KN�2���/L�2� X�ڝ&qf@G���U� �#�񺆣J@r���ѽlЏ��X�p�� �A굵]S��&*�b� ,RAg1��߾|-���6A���C�{{��rƤ.��;V�������g�JWmF�B흮�}�_T�>�~�܂��q�4X�� Ƀu�-<}@�}��E�,�-��Cp�51*��"]�Xa]L�D�\ڲX=Y����(f��V��}`�?�o��
��g/�2O�����1��M����c���^���C�˄ ��Q�*f��_�e��Kjte_��Q����f��1�OZjھƈm�dꦲ"��3fՑÚ�@�b/����S�A�F��Z�#��=`�Q��z��.*���-Y^]W��f�����U&5���~I`��垝�Lܐ���J��Ɗăs9�)���8o���>0ۖd���
D���\��>e�h��	�	{�fN	m0� ����> �5�XB��]N&�l���^�oY
bk&��g��]�� ��� M�8v�,K���Г��A��!��$̄�ƫ�r6frl��#�a��\���dyh�$��[�0�Жƅ��Qʤ���25��r0��!����]�`��bI"Z��5��ĞU"���s>��"4�u��~��D�
��;���8��io_�X��p̬��m��t�K躭���t���L���CDڝ�\��);Yj���A��n��E紁��U8�h8����c��5�QP�12ɼ��^8����*Xx���^�[e�z}��ȗ��Y��F���T1#��Ƙ�5�����|���C�����`X�%냨�d*"z� �h����:��cs�ۨl�����Ɍ��B�:TM�͌��`�#�7�$M�0�1��_��x��S\O�kjm��|��|���� �������_ȉrBV�{��糔��x��e�%�<������c�{�.%���?~"{��̔SƫVW 4f�8G�=�͔mJ���� ����T�x'�jА9�k��$��Gu���@��B�Q��׽l*"l=�,��{�Tkx��������O,x�ħ�����UM,��o~���ޛ����3V=����[�o]���䍼x�KIP�jhkc��lɐ�ð�iV,Kr��@{c����D���hw��q�-@DO y\3>gZ��C�/#OOi�e��������u�x'侂�����JXi�}(��]T�q��'A��ePLܾ�S� �xBGp`���ѹ�0^�/1�9{Pue��]�L�h����������������2���5Co�&���1�lCn<�}��)�l��;"�!_���
PdO/,��vk�����	��pܐ-6��n�v�?���VG�?�%�>�8�d�9��@�	UT�Ӕ%��D1�������x��XR�rqr,O�,�o�.���p0e�\�݋_�Q�J��pM���õg.�X����^��m^ΒI�����9�ԧe�}�)·�{:��g38R����T�������G�,&��x_|�h�u�0Zk�]�����L.\��%��"�A��0���iP��w������s�/�'��( ���\21�ت��o�%' ?W1��i�j�z�y�'�S&�"�桊�ʇ�\�P1�b>�������RWu5J)�7Th��X����;��I��ey뚼~��>P�C}IҪ����uh�B�{v]��V�f�&��5�m����A:��𜎬��ߍyor�{sH\߃b�(K\U�zv/a/�(O�S*g�D�Z*W�z�>����H����7�"S@��WΟ�%��u��KKai�,U�c ���e&$�Bٰ�����Ƈ�Yf�����A�%ƘcC��vv�k\@�x.kWoTZ,Û+Af7����9/�h�(b\CSc�R�}f?} 1#��`黯N�5q�����U�14�~�F��$.�29M�:������;�[�TA���Ji���q��.�ֵ��Wtqi��	Le8 �.��.6����F��s8{L�d�wQkrigSV�-���:�u�卑��B�)6Z �p�&����_h`B�V&�����>��#K�=Q����Z�(�"H�N�+��X����W�� ˃�����g%����:υ/g��^
�w8V���5��fy)ݾ���d�|	-��@��?��
f�I�M�t�2��3�}+���o�*�x�+�}}k[�ݿ#�>�L6�6y����2+�kUdm&n���� �D`���n�+��1 =���˗/y�h�E0<;��>z���A�֋��h\P�Te]#P��+�'��A����ݗW�6yr�j���'`l��`\g?{�yIf��Y���zj3J�Pߔ:�� ��/�@;,��;�4\p��mQ ���L[�R~�ו�RK�F�A�nz
��y�tTb@�O�J���uϥ8�z=*�$�j�v��-�0�EnZ�4�7cc�,!]�A�X�ڀ��R2@��V�L�$�58M"�r8�)���a�
��p~�z6���9)��	�p�T�%�A#�`������k48�+�cf�L ������bS��@�]���2m�����n���h������M�JըVa��RwƴE��w���*Db ����"c�m��+�>��\�3�����J9f`uzz��q"7<�G[� �ԟ�v���Y���}�'�2��ڀkr��@��x ����
�]���5�N��r�w��Eh��r�ĩɘ�0�Ƭ@�˘�  ePb�7C����dp�j����|�z��ψ�l<�{Z���d���N|�və-N�WR}%V
 ���8Hl���>���"��?�����ń��{��,V <�/V�}����פH7����aw��JJV5Be> �M_}�%���W/	�1�f�D�V��0��L�����(��Y R5c�*�ɕ�T�Q��4^�&����V��lt�XQ��&��a�~a��̑�I^)z`}L�����$;��Hks[�n]ȉ��>�V`��*C��
���[K���4:��o�>����{ǜ�ˌ�
x�iW׽鶗�&�3�9�h(g�-��=?gB��l	B�ꍚx��l}��掮�DϞ�f���-s��9�np�����o�54T&MJ�Y �oJ����Ey&���
�$'�yU��Ϝ�7Bd��J����y�+3s �h6m��3)�.����Ո,3C�2;�0�&��<�)�|p3l��Y����֬YF�i6f�����`��Z>��amoneMSc�8���G�B>S�x�m�t��:����3K�l�.B���W���*#�����_M�t�f���g)#l�椶h#������k+�T}�rB���%�@�[?w�F�S� �vj��]w�����#Ǟ=�ѻ�A�Rk��)_2�1��۴Zh�y
>x�m�[���h����gz�A6U-I��JFev\�%����Q�9�I������&�@1��Ֆ����L^���4�ҙ�$-��b���XD
գ0t\V����ȞAQ"q�p�Ċ����X���;�]�٧���&�;��.K}eY>��+�쓏�8��l���7dM�}O����*��qH����z>���쒞�oh�^��ȥ�M��z�s�#6��5��6�VTS���f?w��	�2uH#8�$�*�	�)3'&	"Ë���Y�(3a�.y���FXspD�X�b�m�Q!8����ڛ?Gr&W�yH\T��dU�M6�l�EI+igdZ3�����~�jm����Fݭ��}�}�p�@"ψX�?��̪�4G�`(��8������癩�/��f�����#Q�d��g����}l���@��L�N�l����k���/�N[1�\��ϗ�;2�Y�A�����z���?G �2�}4�6�IQ�b5�VH�i��@��g�@� ��`��z�	F�1�A)��[R= ��:J���` ���j/�3Lд�1x��
<gg��8�"sh�8��؁fݲ`�>�øsʃ��g��ٞ�M��`9� ��fT�=��)�ԼG?h'���/uxM���tHqb��E�][��y4�Lb��YI*�̶���L�X`f�O����;+�a��9���-�ƒ��1*�f���� ҐmE`�cU����9�����zB����`�S�6̶5���j�� �ĸϠ+���ҫD�5I������1�4���_���@�$����E5� ޖL�{WV�Ce��\Pd!��UNP:�������h2�S���cїUt�Yůp֫��+�>c�3��5�^��{�\���L<���gQI���]2$��S7�8fRS}�y��w���ِ��-�ǰט��g�g5�-��7�$-8b�Bš(\h��e7����c�9�Inr�Y6�i��ぎ�&-�z�R��I��g:�<�� 9�9�9_�ۗ���Y�Vc�݁��`��N�!���)�+�AR��F�XO���39yvҕnC���}99x%�ז���7e�]�_S�^�f���HB�j��!�W��	�؂4-�ר�a��_`�5f��J�+���08A�Sy�o��~�(0P�u#��h�� �V ��-y�5��3�&KF��$6�I,�Rm$q�T��|�lBE�7�h�5��̛��)���i�jh h�尥�f#���%���#�ʸoC��p������SQ��%�&�5�5f:Tը5�����WO&��qBc�F�x���g� hU��Co���Js���hT9��'	:��o�� n�㼳A�2M	 G� !�ņ��i)�L�M-̨ي.t�_^]��N����tljhZ�s#�<T����!i �����1�UD�"�I���%��kׯ�%���^�^�q_�t�f�FB��4h�t�rD��,�j}Q�� V��t��7��s�DY��6`�OJP��4=���M�݈
=b��s[�<{ʩ����J�,�d���1G^R3
���Rf�)��:���u�ϲ����ŋg���]w}�ǟ~��E�C^��ޡđ���ؑ{���bp̗_-�5~��:� �}��zy��G<3�_<y,;�8`@�e��?�\�������	��ޣAe\{�S"#YT���:�� HYdͨi1���1z���Pj:��q<�g�K;)�`�Y���AL��="�W�� �N�|�d�|�XF�XS�|����F�L���mY����ǿ���n�9��У��0����aġ�j��ۆ�>:9�ܓ�"���AJS����w�:�����I5��҆��-��Z�
%-�֋�M����3�
(#}^��Ĭ�P��%l�JȥG��`tJ���x`�-��}~�b��΁W��Q�C�somsİť��Q�ʗ5�2�/�i��pr�z�Rk|%+	6�����I5�縰�hz#f�J�,@V�MY��8��4BeדQ��lt6Ȏ� id�F--K��MRK�))W^�ǽ��ܒ�a+(�X`o�6`�.�Xb��ݱI��y�x���� �{����/4*
��5z��\5�2)���}|ߠ�0�>��^}��j��+��·��\�ޫN����h��V�\���QA����& ��a_'5O���ǫ��&׼�"�So��|X��'�{��Zᝨ�0^�A"�S�0��ϩB%����o�.Ь<��������+���to��~�<�y	Q�y�jp�4���Z�vO�Y*�5"2a�����d+��&iK͉�Ӱ�%�(�8��jH}p�1�S��A�������T�V.�����@1�e�(lf'�Ɋ�yR�C���fZ6G ��tC�a�͚�4(>p�b���y���``Uu���z�f��t��sF���Ӣw6I��3|�@�B&;G�bcS��CJ~w/���*���Dj�C�p:�A/�">�W��`������Foi]-�9�W,����-������h�H�L��7#vq�s���(V��Dz�9�M6ł�|��mi��y�T�]��\����!��
4V��P��`�d��)��X�$p��)���e��9w@F���qA馮 ���_qS.��r�XA��9�P���M��.-_�H?�s��N���lSr��qf"fҢڌ4;3��^,��D������:�G�������ˆl�¦���F�d�o���k]Y��k+�<�R�.���� �h\=��`c � C��7�|���C�AV�J��K~VJB�����
^���+S8�3��>��s�a xP3� �hſ��>!��nf�����5-p��`bdc�܁��*($ ��Ŝ���ͻ�!���g�i�#�!K�S����L^�u��MO�Q.��B،������$:�a��l�-�Z_�iB�
_tp�/_��_�[]��=��WB�����������
��6���}X ���]���]}����\_�۷ߑ�k�?T����6�ɑ�����ZW.j�6?ǌ˗_%_|񕮑�x7@ͨs�jĉ�R(��L���PnO�ɥ���*�'6>��pp��\��,�pI^�${h�mX�y���S�A戎�ar�X(3�U��B5F
�YlͶ�(��fYw]��`B!2�h"�����<��@�NR��	hD��2��0��[FG�lW�:�%沧6d�H�#�-�65��S�XԸ/.�hP|���Ҳ��#ϒ:l&�f��uvv�ؑ��nDY@P{P5:R{�ɭ.�s ݘY9҈�&凬��c�a�@ 򭃲�(�L�.��P��|t�i��,5:�ؿ�ӗ$�H��2l�>T��,��@�����jar+m@n�G�Щ� ��*+�_�>�Y�����o�X�N�RЗ�&���+2��!͂�_�N=(SE|_�&_��E*	�AƩ��A���&8�;'��D��2b��NIS��t���S,��!V\���LX��ʮe|��s><9:�@��f���+��E�,) i�6e���jk�9����ή5��,��~�J�R{����e6�c����A�Ь�p�����"i��'}/�MH\q ?PX�����WT+�7'���,+���Q��l7�3�rmG�V	՟���{0�|��`���WU�_�������a�i���*��%:��NSQ����U�������}��y�����#� 4��f>��, ����@aUO�_:��TX $cN5Y��UH&F�J?�=�a�CK���"���$�� �1�����So�ͪa6�꟤dE\�y��?PM@ ��Ww�e�{�i�M�<��ӌ���t���)���E(�(�<둓��㟳��R�2��Վ�) 
@��ߙ�����Mؓ�¼��H��s�R)]��ms l���<x�L���@1�@���̼\�t�s��࠸IfèЉ�B V����H�V�ь�v6Sl����\Pq��qRD�� ��	��
������d�Cw��|r�E�-�.z�!y��֮������l]�_�-k���JG�]]����rJ#,V(��m��!0c�W %6	cҡ��@FeI��.Ⱦ�NNz����T��|Nt�̩waeEV/]V��b��p�Y ���p�E�X���Q�G�e2y]������F��lz�2��e���<
�&�I�=Y�[��W���K�9�<*�H��=�5"ۙ'9�C�'{
����|�ΝbR#��^��JH?4~�`_h�D�	Py��-fU�{��L6�(>��H�!�P�������"s�L&�t%w�.7��Q7��y.�J�ލfUK8��B�h�k��F�6��!��8/y��=����P�"XD��Z��2k��| b�#(�D`�?|�������޵q�0d�N4��������30�9�9`�_���iu��˟��������hRm�>�4l���8;�_�]}��_�tֆ:r��!Fs׬� �WA3J��V��}F�l����R4��:�l�)4�"�E�SF+d��i0�r���[��0��12'V^/��L�Y<k��t*7	A�g�V���z���8��lE=5A�7�!�85���8bk��&vU�&vP��YXϴ"�m���� `��2�Ȋ��==<>���_�w����he��]� TX������x"C� ��ڕ��u����֦�*�w�+�Dj��I�a��r}�\ ��5?c��bF�ⶌ���5'"��[�|y�4}2���}3�d���Q�w�B�(3�����YP��aGʊ��xr��t_��'��iб�x8X�>*�S��ر�ߥ�E&����d�'&"�����
���C󐅌�ѓ�5y��z�sTg jk��(� ��>�s��5��C����jç �96�4�JI��vff	a���Z����V�4�q�+����>3��`� ��p�)��7�w�O&L����J	������B�!$��������{<
ξ�U���<���Y��{JYi��%ZQ�E��յ����ȋ�ϥ{j&��	̇*?���&����Vd��o�Jx�9�Ϫ�K����ȥNm���K�w�V��}+F��wߋ�����J�d����ZZ����<��k�7��:ʯ��+� ||.��3}��-�H�r�����cV�
1�[�=`/��#��UQ{97��ׁ�����0���i�����e%tveMn�yO.(�@��L�wU�9@V��09v��i�9�N4Jg����LWE����d���G"凸�)wXD����ۄ�tV��#�i����]v/ӹ  ޿{SV�����s�~*�8��,�秌:Qrj��<Pcޥ���G��¤0��4��<�R������ږg/�e[�۽�}��>::��FZ�wGn�s���nw0q�9�U��	���!�4%*a� N0Mll���Q�.Y)�h%��"��x��f�V��F#.��\����
�H1@do�����O��O�t�qa����������m�y��v/�Ѡ�j�d	0<���D<���ԜgP#
��p~ �^.�f2��Z�tc��S͂�51S����n�M��;qO �x�ֆ��tS5���_��Oڞ��j�@c*�ft]�i��˲���>S 9 +s8VrF#(�"�t��Rf����i���A;���G5�z	�.U0�Y�������74(\3
>�3��n��cȣ`���j��Ȭ-�4C��GeuϪ�5f��2�����!�.�,��@��,˙��sΊ�+A3֏���I��π�'���=�������/2_�f(�)�y�6����܌��c�TNO�JT�$�zTW�{F �AO��,�k	S*��j0������7i���`\���Tq����DU�@m�>̍2�Sg}�	�؜�$���f��L;d���2`�ft�ɬ�K�XK�eԵ 6�T�,
`�p�� � �-����,��Գ��+�l5����%b��O�m�����T���2��jO��K�:������� �U_�J�W��I-��>8o'�y2 ܻi��� ��1o�q���l�E�����nfj�1%$3�k}�5�����������9i ɤ�<�ǲ�]����B��:},�[�(���GYh~��5������&���||�7a�_�/�1��q �����	 �����#�q���W����Oz��&����8p�V�kk"���]i���^���S��ܻH*aH�7_-�;��= V �{��b���r�?)+�X�i,W�]t��DcbU%0'�a�G���ЬK�%���m�Gdq�W�{�L�����9A��cd�8^$�/-_�[wޕ�����ڔ�ن,-̨�ȼ��Z4'秸��[�3̀�iBa|. <�1�!�k��g��1]��=�sڕSj��Ŭ^���ͩM�W����3��9:=�H����+r����,���5ϊuC|f)ݑW��Fy�q��(��^?����n��ql�2���l�L.F۬�1��AܸM=��E˄-<��V�%ׯߔ�m9R��m��k���ZȜ�uN�C����,c�����|GP[L�pl������PJmptzK�yO���澼P𾱵-G�rx|$��{lZ�&��
<�%N+�֯�M�h�
��4��pL�@޹�����eT�6'���QкE�@���Ȼ�0G):f��|g��j��E��,�s��H��
�^a��9Wu=Ͽ�}����_�� ��w���^9��X	\_<C��~��(6�9��Yx7�n݀V������O�Aw˟U <UBo6,�۷oK�����-�cէi�Si��lpm�ԩ"SNM��?�t<�n� �9@ȱѩ E^+9�ƅ&4�������w�|+��b��z���q�5[`���������,-�9�oaF�EcV���K�Y57�a`�r�v�S�Aj���ϣ�I
i`X�1��|��DY=+748��_|,W�\��/�up��րn�J~�T"�v=�q��I1��( �h�� ��0*4��=6����"Ϟ���E�c6�W��WN�������&(}6��ܙ_���B�,�|�>�X00�-��=�ľ k���t^�A�d+ <���o����n42Z��!3ޠm��� ��'��Tl��Ȑ�����t���>#b�[�+1\���7gD}?V��t�@k��̳�ՆI6���@"���}�>��`�~�#�f'�K5�����}y9S#˜�Z�۪m��O��ܑ�s�}�$�����eS���7�~F�g��XD����C��OcV�3J5dfv^fguM���v���k{sCm��{i���L��>�3��-�~<�����9c}�P�$$R�3�U����8����r�6޹��|��*m�5��!I�J$>?���9�w68$|ꡏί��M���߶N�g����r�E�OE�6<@7E"����&���Țhg'+ �yPw	�5_b=!D���Eze���LN��iD-x���3�@[�s�`; ���*�oZAȪb~_޺7=��)v���t-_�{�v�l�l�����]�奶��˲|A1L�-�]�7���h7g�9�DZ�l�f	a��p�M������tuww_�vv-��0�_����_ �Q��]X��
�/)������Ĉ���^���\IY��YÈ�w�������CE�`���0V_�E;Yb��~"����AsA6}A�ٍ[wd��cy�Q��~v��͌e������?>U�zb��f�a�ff)��r���'�SRF�c�a��L9-��ƶ���b� Gy��W��{�2������B�E��Z�x,u⺍�����3�t�8��D�JM����<��J�z��E9��͚\��*W�.���<�����3z���G#� pxmJP��p뀜v 5W����y����������#`A)F֩?0��p�o86W$��;N��T���]���F������p8X%(�P�;!���`,O�v-����O×M�� )�2V�
��a�r���Y��D#(^�<$GE���Џ���k/�MlY$L��v���A���<J~x�xq|uf�G�p�.������g����O���55�Ah������7B�����jM~�&�S�Va4ٯ�F=p�w9��wv�Fl4��7��\݋gG�rFYO�xۖ�	�x�~���Nwڸw�k��,���Οy-d��j���~E�}g�#_~��c�8 �*Bl����$\b\��jP0������)�q��n�-�'�9a��Z�d��ls*�dl���Ô`m����*�����
��{�@�х Y[�F�0@��4���r�q���-f�8�"Ȥa/����\��Ȉc��z����W�)ٱ�W�xRj��&@_�!^Z��o�7�q���{��wW8�c���m��?M�������7���ϧ9��;�0�p����＇`ڮ����C� ��I�W�]��m���~��3 	����	h�g��Q��������o� [�����X-�y�U� �a>Q�/�1�nY�>c��}�;@Ckf��
ը��AgւT��P22h�;����V�1�'��H�D�{��e�V��{���6x�acI=�t�N�����=���F��*�]u��iMLW���.e W��T}�Hi/1�Y�9î]���5���U;9�4�\D���(�됴�A{ug�
[���k�ee�qDU�j�̞+h�#]����T �YP���ؤT�%��ar�����Z��q��z�JK^������@���s͖|�����o��ۗW������w�3�dyA���'�7�<���XsF�t-���ޅ@�8����+����~��t��֡|�����3y�l]��u���s�|�ܸ��U)�%|/��Hof�$:KU#<�ZV�)��[���V���[-o�uA��q^K��]�����<��Z�e	)e�����Y/la���Ï�w�����ў.XD��ҟ�dqN�(�`�����Ho&����s�!�T��C�b���<ȡ���?�ip 9���+��_ɺ~G@���}k�����r˧�+�v���s�RE�%��<�r�Mw���lG���C��,�eey�
Z�"MP������!j����;7=w���r.�8�8x��
����; �c�d�P���Ǐp���<��D�;>�yj8�� ��gy��c��"�zÍ�dU�Y�yz��X���X�7I�?\u(0,�%�\��Z��X��jT`�����T-M��kDa�������?��I7J�m���od
�A���2�-��������/��w��"G��jV��!��
��шt��0�4l�n��fb����`���)\3
�	Zf=�_r����	wd�t��s8�C�$4Y�K�qpB[ɨ�L������W�$B�ACTO%N�h�s��/ݟƮl�T
ڻ�LX�"G�ŉ�VV�?���&Wn�䠔�D��t�[&C��-!�R�5q�6�����׍�5Ӟc����E��������r����`��s�
2��x*���pP0r��%�cc�&C���#B� ����.01�֮�ba��"]N�ͭ�d����S�ho�%�6��x�Н�_�@��V���?��l0y����� �Ԋg<����_�y�s���Z=�t�1}�����d��`�"����F(ߕW��N[�O��eO�l*0��eQ��m{?WP��|�J�M�� �'����J��>W ���}ؗ0��*ֺW0���6��HTy�.)�k��aO|����j�ZY��K�
���|ZhسUj�g��|�w�^k8����׿�\/+K��7�n�Ҏ������A!qe ��������i��J?bk��_qY坮 ���@b��wߝ�8�'�.�>�������<Vd�>H���u6wc�PN���[�{�@ƮqȪ_�[?{��<�4���ǥ*�teLݧ��4Q�����ND,Ggg�t���;����g����<y��!���C�+�$�-$m��L&*4����z�7��j=�U���M���^�zSn���u���W����?<���<y�.�^��0����U����r��Mŋ-J���pL��H����o�V�q�5�+��[|�0���L7p�n����Q�e�QH�G�2.�N��E��F�n/:��;V�7 ��;�5�9���m��_��tA>��}�གྷ�l��i���~�T{�t�r:E(b�+E�$�,��$ۦ��z�+`���#x?R�wph�ۓ�g��Sy��������}|�/��TQ�,����AUy�[�*sNg�Y2�cf*��B�0"��3���F����r�҃ao�a7dF�d����Y~à��ϟ���E���<Q�xy��棏>�[�nMg���DV �v� @F��;� Ǡ��h��ndu\����`��ӪF�j����M�7���U���:�~�!�d��/�uh�{�P�v�o-��a�� �q��L,p��������*#"� ��(# o6L|!�lP-@�8QǍ�d�c<�?����_�J�i�I*&a��/��N���g|G�G��Z���a��z�pi���_cDՊQЍ}�0bȗb�wԔ���<�E���s0\M�	�[���zp�=���>��f͌� ��A/ߩ8��U�$�C��Ó��"�ƊQ���&��F�<��T�N^p�}pr| ����L��<À*�m�	��H�zbJ�Bk}�L�bt͸6��;'�t��A9|f8�38e,���$ X���e�2n�/�A�\�yΔr�u�m�"� :t���;p��,v���̙��ٶl_K�)Mwxv��/ӋI5���F�42S^JMA�ϣ+��y^�*0ySE�~� �jJi�je�Rp�T+��e��2+�z�����\�7k���t��h��{0�^�VC��cT_�<��B���_R��Ϩ�J��6��]L\MM��|����H���b@*�M�:�TP�м��ONE��V�r��<�q��E�	��9&���9�H}�����Ui�|ݶW恵�y��~�W��l�% 9*(7N���ږ��W���cRAg:s�M�����k�����������1�}w�4:CI�v'~�k1rin��E���ŀ����w�0�	1ѲШM���c�9����Fu�*��Dl���d��h�S*��o���\3���TU�H����OUJM�L���Ǌ���bJh��X��褦L�q�f���N�x\��w8C�xw�����~� H�f�����H8�jV�D�
ɖxdꂸ��]i̜qo ����e9�ó�<_ߖ�O^ʋ�-98:�'
�_l��H����Uy�Ï���?U��(�����`��ǡ�'�� SϾ�V�گw$ʓ�r#�
�-zƺg��0Yҫ����s�x��*�^f����X:@��nN�M?i�\�kgfA>��ʳ�_��'�S��]�(��X��d(�̞�C�8��;��X���Ȃ�!���>��Lr���T��,$ �qw�aWn^���+H}�.�lϥק2#���4����LZ2� X�؀;�h��3Ɓ��W�d}�V���|� He�M5I�\X�*�!�	�9���^J� ڞ�>j'UG��#�?��B�gÛ������J�)���A 0v��>�u�qL�CzFׅ������*����t���kh?��<�&?��'�V��e���g���k����2^&���Xd��*Br�k��"㪆���+��7��&%�3ҕĚQ���(q>��ƀ�S5�菸s��ܸv�c��w��s�ª,�1]X��'�67�4)�yP� 6q-�"���Hl�KfC@����3X�5�L�&P����@�d<T@�PV��I���1��}�]���mݻF�H"��
GJ
Jj���ƛҊ��U0�� �.�p��딁��n>TP�r|� ���?$p�b�LC�I�DՆ�З g�ǞE��i����Ӏ�Uk����Z�N�=xp4���HC0��F�ˬ>7 e�'O��	���L��iY͙Ί,����sQF��m�J�d��l�������"�w�NdO�wU����=f�MŪ����z$�Y�^,�ߧ@%��[��1PfI	�"�d���$O9�5�n)�Y��ъ����x��@��ԝ/앪��	`� <�3�W%�;���O�|��P=�e��\�+2�?�V}p� �Q����7� '�*L����S ݖQϪ�����y��A��2)h2���IА��/�@����v��`����P���=W� D���۞���j�߂/�w�A�/������m�<ȃ�w�5W^ñQ=�?:�/^��&�c�&�,���U��ڪ	���qeI�7W~��k����V�s��j���'�h'���5�;��T�NHM�%�CR�f(�=�U����D�ZM/��+��1���hl;�d�.ɋ��)�o�V��j��7W*޶.p���}�`/�A}�W���/��M�n����K��6KV�/�Ȃ>��v���	Q¦��L����%�2��Ԯg�'���S6���粫�,��/_����_�����Q�.�K�r�{��G��յ�r6�(+<��0T� {�H<ŕ���5�������9��D��=�O?
��K�aD|�ۄ�3O���ZL����T��B	��"d"�(��B��g���r���Y���|&���o��` S��F�D��X����	���%���
�!<oh�����39����Q��ݾ'�>��\�����Y�?P��=�����*���q�4��C)ʅ!pn���HR��@>2U�l��I�HمN�����KT*�x���y���f,�Hl�^�����ßSvɧ��F������
��q/uz�� ީ9�=)�C��+�K�8���� 8��v��iP��1`��.�<�t^������Hbr�������!�,t ,���]i�F4W�
 ���y�6`�t�K�d�&�UϏ�M��Du���?�wf�q?�^��k���ի׸f��_|��S� �.r}������w�𹾫Fm�O�I�H�Pz��A��x�VL���!@���f<��!m��G?ү�F]�V�����u����G ��w4�ѵ �ӭ���
���P���������F	t y]�3��B�����z�J@�xݟ���k���y���ֳ�3���B5:|���9?U���!�^���j3�����E���y�J��¬\S���|���Y��:���[�J�1ӎ�E�0D�>��:�:y5�mβY��b��} ����#p_Y����}�q�3�Y���pP,��bBp��>z�Jz㚜�ɿ�����K[��h�&<�wn]�_|���/.��$Կ ���l��]�&1��[�X  (�p�V 7�e����ܕj��cN���Y�7U�|�L�����4���󪝘.aW��?�QܿM�����]r妬ry��7o��Y���2�o!�C�M�q`ö./�d0	����#i7u} ���Y���=�,`�x�^���KR(�8]�
V٢s��3Dë't@��t�{����l^U>���R����! �;[ۅh�NO
Kf�v����ڡ����>�1$����sb���BY-)�Y�a�>�������㏙��񫴢�D�)�|Ӛ�ﴩ���%1����wyݶ��"�5
s28������l8ힰ�=r�~��q�nKd{T:��/�9?'L��^�-!�ʜp���Ay*�v?LQ&�<��0Wd���}�*L6�4D�pLc
� F&�9����z���������>G�Đ�]Qr��E�9*2��̙"���~%�yń=�9�X@*�
���76��ܷ�xo��{��r�����r��YZ��cӾ�st26Oq�J���Oާ82��'�Lbٲt"�y+�oԐ���9��jC#�LF�Ic�`�����袢9�bFi�q��XNz�tf���G����|��oY�:=;ֈ�Cm��܂�=�VsP6)f��*�uc�.qC�P<���#x �D���.��wߑ;w�]�������Z8�\&K�OBʬA���˩��|�و��7�ᠭJ�뱁w{�y�n6����<9�x�l���v�oE�/D�`6��KK��&�zy�x�&o��SW���w�,6������N����*7����~�4-�e~�.z����x���2��=/�����
�`H٘ku��z5ez��r���=eF�j���S��)(���xG��~q���|��G�N���7�3��vq��k��+	_}���A��i�G_Ae��\�:Y�k[����^dm]�/����-B ���t��b�^'mX�Y������%������$@��ۡTW��V�(�����/!�d����%ۨMP[�Ľ�7��.ֈ��L�F��̜����4�!�BPIxľe&�S�Õ$�pz	A�H6_�����5���P��+�k<&%��K����j����5�;YP��B/�c����Y�����Ay���tXu9�pUA�f�ЃBwm�\��&�+�x��}��%���|H���5pz$�!����~O�gI��< Ҕ4P���L��$����4@Ҭ�P�27b��f���n�gP�*��l�K�ҹ�����;��߬t����i;�`�	o{_\�]y��~�������N��j�W1��>�:z8�̯\���q}�u�K��8��Tdb��;IS��zJ�W!i��g����`����Ë�B��B�R��k$&�1��/�d"�w�Ԫ�U5?6��A�G����/�" ��>��,$6pl�ÿ@���PUP?'�)�D��B��A�g�}ƽ�I��g^*���4]5���ޢ����$  AE���XU�p���ZbJc]���ǽ�ڑW;��Le� 	��_Xϡ�ڳ ��{2�4������i|/��	}g�����T1{��������>0�k��ƃ�J,����TW�ܐ�z�?��ll����_�$��+r��5I�M���j��f�1�o�)�T;���{��K�#�G���<�9�ʫ�-��{�hw�O>�?�T?�;��*;끢6��������&��J_�=�/�B���[|]�FG����|�y�n��������POfK&%�lj�u�G!x>@�2d"5�^�!����t1�z)G���@��n4L>	,�b�C8?% �������=0�55Z�(���c�X��	>�i�.rf� �l4!�5-��d�(3>�����Ф����1AHN>��-�a�9�s|2���,)��9��)%2+��n@�R�ql��n��а�ѩ7��]pΛg�a����(>F̍6
�;�@��q<����j��*Vm���L��36l�S��l��/�����vu�qw#Q]�R����!�3��&��_7��p���H�����|�AaIx1P9Y�����D�O�5�׈�wkc]>��*�\\Y���M�� W3����\]~���<p����2���-{�PS�8�
�����E`
����H����� �P@b��yL�MBٜ��dOaQV.,��w�a&Ҙ��g���@�ƫWs���ck
z�����T �����ɓG�(g�P�jT��t��$A�hh
_XU��JJw*��q^��G�(�N�K+榓� ����y�=�ӵ��tA.]��� :>�b��?!��z��D� *,�������pd��^_R����w9��~���@A5���ζ���i�{����$��!Ӎ�ۂħ����<�{���_X0p�k���z%\Oh�.2� z�I�ݹu�� �?���VG�@���׺������:}.�	pJ��꒸ƆH4�w�}��Ïet8d#xĽNǝe�*�u?!Rd�+� ����`�
����8W)Z����@�M`<�����l߳�߯QX'3�x�	�őU1�n6�fk�d�?��G�&��ˮ�Q���Hn��ʌi��N?��?������QopO���"��;� �|�Z�R��(`X�0�썲����/JVJH:X��y(r}��W�;x�k̺
�7��>�C]��k>LGA3|�=����I �,�>��|���<�� ��||�V���7])���������%�.H�캗�vl���?X5�w��Ҙ�'�t1 ����z#1���3�6����$�����SЗD�@��-���a.��"u������_��{��z]љ�+�8�L�x�_p(�e�V�����h�����ܾ�>m��9�������іtu��V������@����~W��:P���6`�l������� ���r��]�����>"�����O9a��A��Yj��݅9��qio,�8�x5�@�oLb�4h�l%^�v���b^��V?�sO^'8�D%��4p�I����F��1����;?��~�_z,�/�JW7��j2��F�˨9�O|�&=�0�BD�����)���)p�V��,�@�?T#T6����LQ	42����z��xB�8��1X @��*j�9i5A��{^�;���߅{YWha#�:�ʄ:�`�`����+f6P~�s�L:�)B7H �(9�����S�?3���A����{��3�ݳ!��c;���C���Х����yW%Ȫ~��<�L| *DŚƫ�mཨ�DK���Q�\�ʟ:\�9�B#��zq����8%��%�66�������U��Wָ�.�]d;��j,s�'�<��?P>=8�S��R�:3rt�o͗�3w�w(M]���}��k��v}{����	�ByF�_�������N��;���_*�8MC��-+����?�����Yh�1�cvM��ܹ)�ď8�z�Tz��[ڐ S�&�F�U����S�M��m�d0[ _�Hf͞�j��i����X�&΂� ��/>��E9z+.2+��UCv�w�����S�NR�l�k49���Ó���$#��i�!�z�1p�*�(�]b w|pH���E����Ǐ�O�u�)2�J� �9&M�T���}+�~��3J�r^G=�3�1 h � ��d�wn���L^>{.�/�1븤�M���<9?1[�Y`��%g�MS����jTZ6�{ ����>y���R���Br��[��#�jfs:IU=�i`5�`pP�v�J��kz�5��r�jNƂ����$�VΩ�9NWfg�d�Қ,��шY�.^b��P�1��_�֬��&F?�O��fp�~+Ӄ5 �JX��͓!����6{�j-��ͪ����9Y)Y��Y�� 4#Ì���xu��lM�x� � ߠ�����%���~G��_��6�͉�Ze��]mjub_XW��jj���g�?�^�JZ�+�xU��O�%[#�� �0Vi[�oͧ7��� �����Qp����+�4�jQ�cO��C��DAeO�{c���a����-��H#	�l����ϺV5p��M�8�آM��p��`�{��_U��O���?�נ	`6���̶kr��Mj��z�DN���l����M�ÛW[<7ۢB������>�W����SP����p`�����7o�#��G�z� �9P��Yx�pR��޷1o�����e�'0D'^o�1Nlk�4ZU����Kef�����T]�q�	QhV�1�r���'���m��8w�+���%Y[�"{[uq���a�1�ή�A3����_'��A}���y�[X����)��v횴g;<׳�����y��w�li�f�8�WU8k�k��<���Zu���熆����̴#��_)��pd�� � O@����p4����P�_m���ݒ~���E�?�( �1���؜Å����Y.D��/~�f幘*��=C� ��,� �	@9�(H|:�����t ���fp�0�x�4��"��ϩu�2���^�X��L���nK.^X뤁�Y�̓b���q��.�����=y\�}w���g���*BxT)T�{z� ̚�N����!58��Pap��U*�����H��t�@�8'H�Ѕ���5��S���*]O��R�+��7�� 71��� ^�8�.�5��۔���(����=�Yp�d��jz߷w���ʪ̶����>���f�Pqj�a=�Ilj�2�kC�ش�O�ϸD$�Z�Agh�N[ր6�{݁ �"��]gZY#{|Q����ʉW[�B�n.CNB�.�7}� ��@�58���#��wo��w��\ý���/��=���H 8~��{@\c��4�΅SF�þ�@�T������F5�67�@>��c����7//ښ��=����}�V0������z�,e�8K����>��U��O�? ��#f�a�]W�͹�!�Ά��HW���'�ҟƽ�T���z�߻�s�WKʀo�*bG�ZR����զ����"����ɿ�+[R�����T?�X��~@��ySϪ�jo��E�
��w|��Q�pcF��MyhPDu�P�����gG.4|MnR���'�sa��z���\�A������vX�
�6�5.#�=����^���L4��N�A������-���>�C�C|}��3p||��:(F �
����,��nB�����)ֹ�����^�:+��41�Z��6	�wOd�4g�5\#X�D��]�^g����c������t͂��k�c4�`ђ�A��1ɓ��AU,�=���B�[)e3&�"\_R�c�^����X2��c)Ax�S��\f3�0��Uv\�ay��Ҝ-2� G�sp�ޞ��*�-t�'�Tp"�����־�\�~���\���|,��ӳ����&?��0Tʮ(FYVv��u�_���m��`ю�N��qr��B��(.�Q��D�w$�p��`E�N�w?A��1�5�}U��T3��zSv�":���k�5/�Tc �?��0�� ���	�IcN�Zsܬs��8a�����c:�>�c�`l���Թ��������ˢ�י���(�BC��)Q�1�7�  ����"��{���X~? "(�h*32���t$�#m�q�Zc�g!-�)�
��u��8p�a��XO&K�^�t:�{�hྀ���φ{��c���,އc �Ðt;����Bc�̀:|�gK�Y.��s��P�G�9�
�`�>��Щ>��L����bM�!�M�؋��dAi�Ɍ' ��}?���*Go�՞r�0M�}�XSc�W�����1��u�2�hl
-�Xۻ{��}��yh6C1�<s�a���x�TvA���оm#8!��8��`���'�l75��
Z�0�pV4>AEeԧQ¤:Lm"+�����E#��20]Z��Syet&G�99���g7��sޢ�C~�:j E��A�i�r�ѐ���\{F����W ��P���E5��:�S��kf�1U�ղ��I�~�ǙV��h��cD�N��A>@�y���^�g������lV��*S��l��q}�ٝ��X����<���8�=V�4h`x��Gf���w���)�\4�a�a/���\��Q��F�<̅ �
k��+�&j"@��� ''FC���Ѿ���;W���Fxp?1yЕE��:���js[���ȣQb��a���8���Z�:����Bf������S0<S\�M�H?�{�?fk�q1����t#��q��*@��������p��g��+5��0�>n���3�a�_�`<���B0�a�;+{GF�J7��^P�b���¬ ���ng!g��G�aj���hX$]ܟ�ͭ��r�X�w�v���p�{��ɽ��b�~ך�_�^����~NA�τ}��C"i�`�{vN��`=8�{�� @￮\�F߄�v�t|!`���y�m5�4]E*�wj�e�^T��aa���<��g�F���H�@i�z�_�+}�f�z�E��
-�.�Qɩ�|��vҪ�#&B"��*�j�Ћ�VT���6M)�d��Dz}��e��0�����^��/���)G�t]�rT8����M#� ���r��Tσ��f�t�( ��=T �S_צZ"�y�;���`�teM@��,�C��\������$)�@���o�-��|�a���=�<�a�L�i��$�N�<%����C#[ȟ�M���Zې���������Vd��M�G�k�>�1��jd�{g�4ה��YX]��)�?9���Cf�0�k썛�P�hJkvNfg:
���܁����Ț_�q�ϡ����+	J"d�d�~`��|�L�L{�M]F����������KO ����@7Nh\�����Ds��=�C�{q��ЄOOO謯_�)��կ8��y�x9��������D9͔0n ���y��a ���QR��?�3f�a�XN�Jn:�g���{��G��o߾MC��kq|Gi�3��4�,l�;�p	0w ���JV��:x��$5�`�J#<-�f/WX6*Nl�ʞ����8�9*@�O��}�����%��9���@WHbv��dIӀ�O����Y*�$�èX��-cU�Z�Yw�d��o[տu0c��r�Ś�ų���G ��{d�Ӓ��y�ܣ�}6�r(��oT���p��ǁ��ý}9:8dƳ��ۀ�]jk{��A��Q����B�p� �
N��~���+n�q�^ct4Њ��]�,�fФ[�Xo�C��C�dcs]��7Xb>�������kp]�^Z�N2�AGs����ɪ��C�8�q���iO�vO��O�T�T�v�3G{3��, �q�4�}���?RqM�w9}�:�d8�~|�}��{�=6�"p�?�c%�;�*��2�q��P��v�C�λ)��/ן�kIm�HLA�	�xTG����@_0V�~l�V���F�1޻ۨ�r�9;��L�4x{��I�ƫ
��C���o�5����~?%`.U�&_o�̻���)[_T�dJ?��0F�T�I�§�v��y�Fl����3�L����8BD�Ҟl���8`��E�N�&ǥ�{a�X�n�p4Ө����+�r�9��DYDX�W9��t&�ӑ��z��Ԅ`�P��@ڥ����ɦ����L<�.�y�y �*"�SHye_��[/\U��ݺuKn޹���r������D��뀨|���b2����������c2�Cl�Q�q��E%	�l\����+&\� }
C3AABc@Ic�lIÑ���7��$7��W�Њ�eA\��2��<x	�d�I��4�jo�u�$N�TYn8��Qor�|nk�'s8�*��q��k�˕���krq�2���g'G�ՕDqL{�\��9�����^]�H��ud�O�ӄ��v��r�:#���>�4�$_'E5?\��,T�R��NW �[|�w%�DՓZ�e����Kʁs��	<(5�������`ȳ��4����h����,��O�,��!�u���8���d��>?����@��R$x��ڢ��Ή�����a'��6ь��[c��۳��ˌlč��zF�{�s��=���ε�-���{8d )�v<���by���C��.k�pd!��[k�����(�p�sk2�������R�@�]�.���	�#6Z���>�v`�q�QVN3���{A�����+���vP�πQ�s�1 �Y�����g� ������plDd,atq<�v5�nL]c���0����~�G����jQ�l��b�N�9�Z�P>j�?�reT�(H4	�}���p/�.m�2#�m�ȑa�v�����1h�h�9��
G�:+&bf�*=z�D6�=��;rau�ΗϙCz���jP1�E8b}�B[��b�O���YZ1.���F()ꂕEP�"�����a�
�ru�Dn^� ���r�ꪂ�Hκ�\[�b��od��O��o*�VG����&9�}}�I�(Y�G9H�݃0f��!�^���غL���t����>�x r��2#�$B���@&�x/]X��F�Y��dv�)�5 ��縬�UvL*,��L���ʃ�/崧���tB33m>G��_�vE��Z�2+�c.^�hq>,3��Qo���AHK޼~]nݼ���;��(�vz���+#�o�7��dac/ao��|��7�4-/~�� ���M}~g�� ٱ�}�jiF�L��v��_W�q�f�?�� Z��I:�t6�����4Yu���S���Cd��fX�w��f&�U���
��k��3C��@8O�W��P�Ώea~I^�Z�����z!��EZ%8��q�\$n�3�9! (�kX�~�8�HJ���~4�B/6*"�	�8�8�i�ȚNj�'�^���� ~ɢj�M��_�(��OKu��/���7��|a�`���?��<{�\
�0���	)�!�� � ���3�o#�~�ZH��7��WL��챭��o��Iȓ���**�y� �.{���\���9}��s��[ ==�fΜ	kT��4��1�^���E*g��Ը�UfL]�Cu/V-�&�}��羆94* �rH�10�k�}���8
�Q�&i���)3mf����&��l2-�U��3�j�T?ǔB�v�=MX�Ӏ,q�O!�������=�^�(B�R��`�`��`_p(ڨ�cE
�I�̂�Nh�ܸ�)���'�o�L&�
��P��,�UqH��<(�u��R��eB^ں���&�r"�,\؀�\��4�Zjq��:�d`q�����[����>f��vL>���I�h�i��0-L
�7L��D42�4,,˕Re��kڳ�-p��8�(�j�c� QVwh���>$gT�Rd����Cf�jQ�cf�$/Oq�ȘwP1D�s�!��[v�2�V���#���A�9��Û}f(�#{��ec�����'y�g�{&�#k�Zc��L ���a�.*��|�*#a&a��<~w ��v�@�����Gz�c��*^0�0�n�a�`,���R�g�}��;oM�����o�9{�ԍ���tY�Mj��X�s7G��	�Vkx����3tQ�̄ƂQ�$��� �� ��y��k�}"{j���?�'�5�DYouiY�����xgeeu�&v�)�pT��><:���V�����^���:���!��y5�)�(hȕ�g�������U��j��i���5u�T�I^k�ѳ,��E�T�G,G"K�#��-.��B�1ٱ���[�n((\�����9�=y��M�taE~������}9���$�?��o�ɓg�K�K�R���<8�}æ�%��ٹ6�g���Y�h0�
\�I�m8y��U�,3$���2���{�|������}�P�\;�� �jM���ƃ��13���s��;����M�U���u�l���]^X$��r���.ʳ����Ŷ>�%u*
�{#�1�x_�];s�@!;g9���P��EY����ok gSlc�"H2���5��֬i���29р���gr|t �޿+�~���r~aF��!�>q�A�A���< ��*I�fΌ.�AJ�"�W ]>�%�<�d���(��T�7��g*9����i0�z�ޒ0A�˫�Hl`@�ڢ�7̫=ꇠA�������r������h6'ep(2�0�?�Y�*A؁�!RV�ˊx���M�����F��-����<���S�M�=#)Ʒ�s�o���g��u�0�{��̢ܸ=&��"ǩ�Y���	����l�	[1����_ �1?��g������bUϡ%��*A` �L �#���9�3��t�r�y��y�<�08�*�� �����}�>�m��U��׵|vJ�%�ݎ�����O��2���\ˎ�N��j/��JfE�fG#��ݽ=�{���16W�<�"x!8�)�����1��J��8��4�:�;��َ�y��q+���0:���54�B&qLGB���n�;�e�,��I8[�?�l"����r��k�ULC���bҼ�["��q��!�|oL����譠@�����< K���̙1���e�F���}�OH����z��zC�x\��<�T4�ī�����E ;@C0+&��8
���Ԕ�N���.ThPA�0�_�b�F����k*�ƚ^^��L��Ph�d4ޞ�O(Z�wc̔{������y�'��A�7�"+E�m)�)������;?S�tF'�i�5E�.��C�ԍ	�4.�2�d��A���a�;L�&�W' MB3lƌ9@�0����WH>�`eՠbCz�w�B�TW�
�!�7��Mb<,3c��.��EJ�]�`A����6�I4��t���p<�=B����Ѡ(O���8��T���5^������_��O�.�j�P�i�C����7���l/�*0L�#�	�	�Zߴ|F�H0��TɈ��7����ՆR��
Ѓ�@��c��Ľs�|�z�;>� x戊1,��F�h���2���'e���C��J�rÂH[�dҜ���nF�؄�nq�l�{rtv$g�;�9��믿�͍��[�:�Ms����A[b���t���dͽ�}y�����s���������q���3��hc�3^�|�)����,�jl�f`�fF4jg�=0R��4nn,�^������c�r@��{z�sI���jp0��	��S����܂�л@'�u�4�o��:���,u�5[P���2rf(shd��ԍp` �Zz�-�[��q��}�z�
�
�0X�X�
��"�A����f�֖9Dp>P�=8�����n�7`�=t��|��+|ngaNn�osm��XP��������� ��x.��N�]�B	��.�R�h�ҡ��]g�̉�sЈ���DGL'i��kzM�V�r�)Iao?y�Hn޹�������"��̝���F��#�����~y]�EXU��fI}(@YT�(;��{wt�o�ϡ���ԝc�ͽ���1�4ٌ��I��������g	��W�ȉ��V�2>_�5ҙ��^�rU�.��Nr6�7���	��.u/g&2��,y��v�����n=G9�U褠kF�8�W �7�����M=v�j�{��r�,1V�e!Tb�����x�ʮi��=m��Y�o��_Zd��5��Z`#�߻���8d�q��s���]Q����ѦR�F��Td��~o�N�u�M���(�/�7���D��꿇��p��h��{��	������[���M&\�|9dU�U#4��ఎ +\�<�5N��fE�sg��ty	���!�+[�(s�cf�%���qX�!���f����v��8���P�{��M�q���G�P��Fտ8�
J3�a�"<�&��6/$b	�cJ8��H�w�Q��6&�w��/��f\И��B=(�,q�+-I��}`�|�=�٢��0a���Or�k���x1kTm� ?�|8E�$d�}AP����T�hs�I*�'����������-jQ����:glC�Mkf^|x 6���e��j �.XO3�<a���>*�~6�X�<�:!8O��	Y�د;*�JxͨO ���g�9W�u����i�lDS��_�&ޢ6LK��<Y��̻���K�8L�?�@�t�O��1�v��g �0Jh���:z֛:��:]�c?LHuÌ����=%x��wg MA=�#�8-�0�&�}ƹ������C��~C�ߣ�鍮��A��/��{�D�׭!�����a,I<))�'�%v?��"�VqԖa��L�,`�]���8{ ̓G��f[6��c36N���I�w�=�<K�`�������IW׈]��޵��Ľ�#�S@���h�ޡ�~F`����Կ����^pF*֘��L�r�n��
U����Qo빞m��3�I-��"(O0��� ��L����ի�4������"���C &a\|+�.��`�a���1\j�#�˛���S�VK���j��{Ʀ�>*6�̡v5�F�Y�c:�ǁ&z�٦��#βe���c�ST5 ֿk�: ��ѳ�H{t�=�>/8�ް'��{W�߽'�����ߎdk���xa�!`FF��$di��d >3l�5�z ���֮�?|aOc�"Ӊj �%�zA5��aP^N�ȡ��@s���o}z4���Ȋ{��]��&��T�9�[/� ��|��a�
��@"*�+��^�Y��FR�t{퉂��q��J��C�?C�?M%)Ԯ�7+�Tin��Ρ����VК�vv����^��k�co�b�*�QI@0��a }�X�M��\�K2ԉhL_�J@f�	��T^Yp*\�(�� �Wn~�Aw�7���@���:��٩�[H��tV���a�q�P^p��7>�}�W{��o��TE�N sp�= �}���׿�5��N�<��C���~�?��?'M�]�jgnKp\��O�E��Z�B�P�̳Y_}��� �fS� ��P��f�X�P�Ȫ�3��`���,��J�:�{(�����y��'�����4����S����3Pa�ֶ�V1��QF��cÓ�5N~{nu:�0�>G�;�Y}Ν�9������:�w2�T�������Ae$�]l�ہ$	}��z�g�j	��C���K��6J
 ���U�$f�!P�`6���RD�.쬄�2aE�`��=]��$p�Hg&���s�G�xE��1�5v��ګEdE�$�-�J�!
�<��g�[Bi�����l>{ ��ŕ�Th4\�q��ep8��ˌ2 fe���X5BSM�Tp����[x<V��Q���b'�W�P���,����}h4��Y���tcͶ�2�6=6dc�+�!'��0�	��Uʫ�ˍw�)�ưekc�}<��n�{Y��� �8�_��_�Q���%_���dM�T�I�����!��$��7u��.5�5���� F�\���x���)o��E���O?�g����J��߃
wL6VyT4�:����Ue���&��9{�Uz@�wU����="����'x��-A<K��,�����u_�B�TSh�C��p_�
ʯ��ȟ|�+y����BS�(�]���+�>���4t���
�p�j�)|��4M7���k���g�ǳ�>��ڵ����q��3@�$��Z|hXV��}����h��������o��'�z��R�0|��up"��r���re�B����n�i
�S�|p��_f��w���+��Mu�����F����;9,*�Â]�)��GVI5��G,U��v�5̊���":����k�ʶ������Y�B������?�b��ݻ���C�����xiY��k�S��g�H�P��BPqp��N�/�{;���3��=�dG���{�Ԣ2KWWk��d�lr�|�����v����a�0�$�C��f�.�RTʈȐ.�αk��U\��Y�!\�k�رcHf�y�m��5;>:�rՇ~(�0%�
�/8��p-�|�c�\���,MH�b4a�jA�B8޼�*Nb��I�)��U as"ɴq i������lm��k�[�����F�|�S5]���>Ц�]Z<?�O=X���;����6z����/~��m�{��`�����;�&)��\�����Р���p8�P��'U�;���);�2��Vq��`]�$SX�=GX���������jx�����=-*�W�}A����7�Pe�.Px���R����Ѽ�	�#�N��y!X�/������@r
4�a��H�����'��8/�v�O�F���	������S���GC-�҄��R�л�ɋE��s@��sB ��Cefy���F%�sx�R�)}���X����^��f����ʷ}o�5E��E���-��8_�y��\cB��=�ާ��k���Hʞ>��,)��bXgK}���y�1���bL�Y��X�����W��
����Ѓ�dhft.^O	���&�ѷ�5(!R�h0�z7&�u�T�lV����V������[K[��>�~�3Y�ْtj�h�($�E��]�~/��k�l6�sM�ՙjlbA$n6�d\Pm+[�GYZ�����Ae�(F���C\�t:�^���:yɤޤ.,4��V"��:<����}�~���@�.2θUkl1GI��,���Cw/�L��k�]p�/��gbω-Ihho|��]���_�5�@��g@�Sk�,B9������JZ�78��^/N� ��P�qB�ğ[u3/���f�Y����
�ڷ�}�DH`h�� �f9_����$l���{��Y@��FeOY�ti����9X�@|��x�||����y�l��10�pV@�!�ϷN���!"ϩ�f�dy5�ʞ�d�T�<Դ�����Y_�w�9���mi���0��"�˽�5Ɔ�X&&�Ղ���4�
��O?#��M�iN$����{Mn��&��ˣ�����{�H-�=�Teiu��A<E���L��M2����N%�����'�F��*#����}c[VV;2�C�.SXg��SM&\/�d�P����_YV"9~}m~�&�������Tp-�\-��Ԉ\��/R���ψ��6N��3R�F�\������o�L*OV�o�KT`г�#y�*é����$KH}�h�u��3��3�9���/���`U��~��E�_��`���Wn]ߕUM�'㠾TX3�-���>���=�%��/(-�ʩ�}�9����v����_+/���ڵ�R
{��W�t:��(��ƼOP��'�k�_���8�c��� ��\�����{5e��胹��S�Jq�?]�ё��t�u�������=�_~��_��������O��*�oTWe`j(���ֶܽ�l�����t��ٽv����"���Y�\��7o��k7emeI���%e-{�(a�f��|�k�Xı��R<	�=�wD֏��H-��e��6�%脨��9��G��������I?s�捲���Ĝ(�,&G�Y���V��o�&���o���� �w�w�8<(_��~w��>���_��Lp�؋x.+�������l�&y �#��� `g���M4 ҏ��s��67�������)�H��h�?�cF��xg٬�&^�^�)aА���f�`�'�Ӳ .`Z�I}s��^���"v@3
�,���v�/t�D�	�Fl`(��@^>�/���r��=.0S�'(��&���jbi*�*�-�	�=�K_��*\Vu����m��!~#J[���	
 ��w��q���?'M:W���[�esk����~n*z~������Wo�� ^�
5>�Z���|vNRH���^�4�j̆B��&�
�N�#if@9��B�K��^�$��F�2��F�a�O�@P��"��[�XF��!���H��:�����Y(��]����,�@������ԛ5i�r�������{�'wM�"Y����@�)"�S��[�E*�#�����|^^u��Q@=p7��('ᡏ FA:2}8�q��t����+5�dRk�rt?�ʇߑ�8��h�7yU� C��8�\���yx7x��_�@{��	����*1pMT�h���p�f�\M���8Qd�\G��Y�6�4�HN􎃗�2=��)>��koʁ:�ӓ#��5[1y֣�j֢A|}u��6'��a�on�hŰ�.<f�{��B��F�D�ۃe�R�)��:����j�72r��������+w�^�`���Cy��!_������=!���z�(�c����i5�{��oXC+K��߫S��O���E����NE�D�)_������	b�l�s�Aah^ES����YY:�=�e�8s��ī31iyH�^�勯ȗ�����@��5�C�O�\�����P���ϟ�����s�+���mpPu O��K�H�qSnݸA{��~�#yK�Q9�2�!\�n�4_y���;��뫍���&9�H3�\8 �7nܢR�%ę��2A�=-�h�( ^�iѡ%�n�@*�����Lc�|D*�ӌ��њ=[��W�N����k�ϫ'羶�*�6�^��O
����=.#���}���Q��^����@)�\^a��L�ӗ_}C����)�jh�|ytF�t4�XB����p ��=/t�����T����7U4��r�w�a��2 ��y�*�[��(�ٟ�	��'��dlO��O�C��������y�]k�N�rҶ��`�T��_g����T"��`_�����R�>�	vt�^�V�C��Z�령�JW��p)�]bОI9I֓V:�����`���
��>ѕ��F��;� B�\�)'e����!.�r_����e�����tQ��r<aq�ߟ*f�y4"r����dw\��-��B�M#��>�*6�FƷ1^zD�6���z͹&jz^2yVc>&(�����(�I\V��@�8/��A��8*oUj� ���1��k��"7���vUEZ\�{��7�1�w;�͍5=ι��T�3�!��k�]4k�W����<_���$[]Wq��G��v�T��a�Z���}#����i��� K,��"N�C`�/����QQ ��k%�t�l
�[��.�.��
���
`��y&o���b/�H��5�V��}>n
�;HҦf���1�f|����������7��ʀ{߀� ���Q��ꁥ;�W�x���MQ9����V���;b�Ϡ<$З$._���Hv��%U^��CG=Jz3���EPB�҇^�Qr#�=]���v���>��5������y ����465G�U�W���ͼ��c5�R�r��q��^y�
��fD�Ћ�@i]��^=zm&��]9��cm����ĭ�u���g4,c5$WHk�Ý�ɬ�n�>���R�it>-)Eا	�"}pT���Mt��)x�N�[�
�`���&�3�#K�N����|��O�|��7�3�LK \7wo��<M��?�����}	�z�#�R%���BB�D��`80噐�q>�@Ӏ>|���%�'y~�K�������T��� ��D�G�~�*��V��Ea��R �qM�p�� ~x����������� 9��gt���lx�r���������~���SX�h4��x�=��r��{t|j�g�E{rvޗ>���R9���CA$ jM��C�����/��r��}�e�*�*���/�$�;k:a�'
���r��=Q�@�)�zH��Rdj���[�K�{/V��Aο[�]QL��ܚ����kb�^l@�k^��7B����E��E)�X,�y��q��uɩ�=��݇O�j���8gB��pȪ���A)���~���ً=��X�va�i@61a�b4�F��y�# 5q��������~���.7E��S��{Ol;��Ӹ��������7�@�+P���&U`屋S�(%�v	>�C������	�h���q�����^�
dp�a�8zx�fۋ�P�z��b8,�l@��}±��[ �X�	��>���y%��>h0TLjZe��"�i�������'O�YC���'�4��k=hbp��i9	��OYP������D2���~o1���S�$�x�{�b�ׅ�f
�;Pm�1^���Ƅ~C�����0����s����B^}>3�^=T���'>"�cD����6��O��%�$┚��\w!!
�Xl��/����l��VL�G��*e��
x(��B*Ф��M�l!�_f��30Q�;�Ay���K�s��cH�A����CߜYV���GE� bxA�_�6���e�.|v�Zf=�RK����0�(o�e�1�wM�����dqF>�D�/�Iϐ9��ĕ�C=*��Q�-H��N�u�CT^+M�H�h'<?/3�d�����Q;����[�*�����1��`0���y�^���J2�PU�nmy�l0u��/>���@�bxc+ʀ>��N�����86PG��P�Z�*�F�υ�<d�n�(E(�4i�:O�j�q~PoO *Ģ�M���@�\��u�Z9?=&�&34��Ta�^;�H!��s��|�Σv����u'g}Y�X�;w��DM	Z�(�c� �����޸�|6/K�X�D��f�]�`�8CvZ���v��&>WOn�髚�C����� Ù�4`�Ѹ/�l����nk�Oe��#M����t���(�%G�.��|��>��bOk0����:զ�����V�qXľ����_3IY��{
d�wc��&�U�@-Z��� ��U�@	�������������KdM�h����c�3y��_gz=�w�ē�t���	W���8�`y<3	���M��D���ϵ��,�L����O�@���D���Olz�����s�� ��`\���X��%{Hl,P��5_�M�p^�=��$��:ԣ����hy:�k|����t���I�"&aʠ�$��[��2��t�c��ߦ�Zt{�^����\F�/�m�����UY��i���x�λ	��kk��YC��������ޘM�Z��؃b>�zf��� g�W.=M�CƔ�1Sz{��ytr@{o�:M��ɽO�_���' _�B�cŭN��{ o�hl�MF%�
�-�õ�����fSk 
�r���z�n��w=�����ᜡ�6�n�Qfp���~��߳�2��W���|>�A?� I69����}K/�;`�	�&�Y��ں�����1�Fj S��1<�p���h�����ky��������/���	=$��+QUD>���PE3 /��~*�\^U	,���Y��ekz=1P�⷗;��"{^����\��h35 XK���h�A����n>���濃�<T����R���S��a�>�y����X��;�ĳ<H�ۼ��@Hb1���'(BF�!���/��!� �}�Y�Ĥw�?�� �"ɱ������*4M4K� /FeS�����B�%
�o�i����h�Ů:��Kٟ�:���fP��'�pt9���qb��D�#�΃$RJQ�B<��+#�</����C�f�Ѝ��D��̦iŖ��Ʋz ��`p����l>iЈ6��o�aa�
:��J%��ipyQkH�85�Pr��YҪ ��%�M�8����|�	9��D�{xxd?�5��mT�z?/�����a`\�}���wIH ����2��;E4�ൠ�x��Gp�ÇR8���f��{@5 �H<)��4���u��B� ��r�x����tf�a�,6#hp:h�C':�\����ɑmR��+��9sa���t�5�	~D��\��F�C�?�ѻr��'_~���T��I�4zK�B*��%�������������*;�os'�@��u\������g�&��i�Pj�(��oq��Dl�S�ی(��\LC����}.�6R������1�3	�/0���_P/zM��i�Oh��i���!Iym
��O0�O\��U�����s��Q}8P<gҲ�L�ߚ�#���@��z�H�2�G������'Fk�����gO_ ࡃ�	������;��������Y�BDV5�%#˓�]�z@��3�I45`�Qn���U����ޛ�|��j裚�m[���_��#V&c���޺��q�!�k
�m�����5rrw�ݤv4��|�D<�'/5i�^
t�N�r���rkm�2P�}T{�j�ИF��mⴴ8*ݪ�e�w�Q�i�CtL[<��o�z�FJ\�줩N�jo|��J؜�ٌ$����y��l#D��l�ģ�년���fy4r]:�,?��M��xp� �fٴ����Z���֣���ĂA����XJK��2�ep���hQ)ɏ{6�h4g�2ܒݵ����d��@�3CB���<�D�*Vy�D�rrfSI�* )�,.UV4QF�)�/d3�<{J�|A�r�8E��r������W�p���k��ο�뿒׎&V���9��H�\��?���Y�7��� ����+<�������=�Ѷ\H�
�s���뻵Tq���Փ���Ve7�^�/>�F~������#��T?����t_�_7�gש���.�����2��	����H�3Jc0���@®��j�cO��	�[l��>�t�2�����<�{ε��}�S����H%$����/UEoC! ��7&=9��jXJ�<�� ��S(3R5f$!�/�-��ԝs�a��s�h���dD��6�l2�Y�dAl�=��F"���C��V�3����i4����h�)�H6���.sd��be��������@n|dz�@�0�6�J�����\O^B��x��Mo٢��~v[6}1�������[+5#PX�kIAIl�X���ͦ���%�v����1��smN�mp���,-sXլ�TW�� #1e�m�*�&��ο��^:�P�&TJ��fy(���L��l�F���kH��n�)�d����;������W�� ' �Wo\g �6�c޵KOz�σmG��z���T<�@40��<�(�c	�`�������3��d��ݑxoS ������ �a���x�zo���qyܸ�V���"&�����6��k��0C��[���_^�Mk`ee�eV�S<��[݇{�������ٖ�+�l��`Â���/i��su1��N�x��5��<�GR&R 4@�:�G��VC�{��cM"N�C#
y" %����Ta�
6� ��zq�`�ENM�5�����#N!�
��8.Lc�Aw�(e�*���H�L�2�N ��Ĵ��;?�4�Y��8<؃�U��"������mP�Ap��i|��4�=�a�/�|@c~�c ;� L�h�\�X�S�Z"�����J�0�:�mD��z����n�yS~�O�M�<~H{���/*��aF���n#�CC"8��ou-�<�ϜJ����`$gz\/�ਸ਼�|8ar�Qg�y��;r�vVU��ή�����U-"5���N%)��>�(3;\��|{\E���['\��%n�pU-��鶒�Z�ԫ=��H�	���ap8�M��!����:�;��/W��k.˵��P�D����:���Ǌhl�k e�$��*�t^�@Nن-Y����ҿ�RvL��Fր*��'�]
SW��q��c�yߓ�;�?@r?��<0���ʂ��� ����Ac�}x�9&ا���]��O(E�x��m��Z��$^��A�,�]�p,�3^��S2RAv��y�=�W������.7鯭W���ǭ��"��	�%Pq�r�A<���3�Z��L�a-�M��@�]��6��tD�'�U��D��š����~=�	(zu�5#��t�|��UO�f�4k�)[$x�e�18,��R���Q5��T\ڎ��4�ð=@��>2�Ğmb
wSZܳj����z-Z�4�tۤ�%��u:�d��m�
�>���]f	+>9nr݃..��L��S�Mm~L_�Y5�0e7?u*�䱆��?�?�EQ6�'��1J�e]���;ň�<c�
 �f����?B���*[���p�L��dҠ#Ey!�P�%% �Ӕ<�@u`2A�Ve��֓/���Ґ=�T�j�b3�0��s�Z�#�d����hv��?c��X�C��c����Wm1��o�1	����{nrF�d�^��ί�M��K.7��.Q���X�NN͈4%j�T�������F�y�>	���%I^��6͞����X�y��D������O�ܼ}�ρ��<���rcQ�u�A+��qM��I x|G������@�u��=Û!A�zԥ�L�����]٣Œ#�zX�h���%����!�B9mU�aPS!���(�qW��َ��y.u��p|�Q9�7��I�ao0j�ܕ���"G�H�����?���g_~!��:U�+�8��#�ڇ�p;�7o�)wn^�u�a?C99> ��9=M�� @��_\��>(a�����2�gU�r���p��bs�+O���^��D:����F ��O�Bţ��mM�d��U^0�bK�	\�9
�n��:���|$��ʓ���5�UӛCB�h��>M�X)d���ףQh���'(�h�p^hP�$�[�o�G?��&]7������Q'N%84c�>��z��k�9�K4�^h�^"��9ݕ5ٹvS�\�I����t.��z���x���m����a݀;]�B��)pv�3�WKK�1�{Y������UN޿Îlmm����C9�92�5�"ܐ�Y9Ȃ��r�g��U8�ˀA�d:*�z�%!PMB��h<PWL�ݐy��J%-�9����\ypd���Y��S� �Q,��}�ki���fU�-]J���6:�Imf��_�������uz
��#Y^��#��S,�dp|̓�T=���*@��}����sYX&'����HX� f 4ܺs�T:��@� v�Qe�D���ܧ�x�~�p��=��,�6�s}xղ ��N���C}�T�\ ��7�mT�aSX�{�Ւz�ROi����U��K���ˊ(f��;�{�9�'��㱶�-� U��I�<4��;c4�AEoӦ^#�P�كq�w��/a?T�������3Y���v��a[ރyC�i�3����&�j�Hc�y��l�8�6+_]k\%m5+i�V����8V�a�a�|BmȨܳ�$�ʑ8�S�A����ޭ���=9S|��HNO�#�i�C?�T���cbW���Ə���z��#i��RJX�{�ボr��ĺ1y��i�� ��xv�1�oFTM�r$�o���[	��^����Pַ�2�fiM�h�mfRz�d�������?tf']���xvmԝ�4�fE9	�58�LϦ�dļ\t��d6��쥦Ms�8$I?#Ai��W㸱Ig��Rq�ȡ�r[��!���8���Ҕ�(
7^�*|ڭ�Q3�0
M3V�\t��0CPs�aG�:��q-!+z�����K���+7b���c�4#pr�7�� ���G%ѵ{��E	y�`�g�;�	��9��@�q.�L��??�9���޴��T�JbR��y����@�((_i�hw�@����6�%i�i�:��� �#�FZ�j�,W?y��S���y|v*�[��>ٵ0	��� ��8	�@�̉�"���B41vP����G�c?�������&oI��(^7˭w�t
6���m��Gu��U��A;�G�\s+���u� �5���U��1�;�5O�=���wlfu*���p�ֺ����:�����g��\��7����`�Q�:ӆMs�z�L�m��ܦ��M[K&��ay��B[����|y_��޷�jM��_`��F���Ѝ�Y�v��2 q��!�Z�x�L̣q���|��7rr�g�F��Q
�I�b3y�t���x��k�L���=}�$�k[���YZW甛��.(�̲���SNlY?��Y2����1NϘ�C��n��P�5�LB1
�Ϻm�z�Z��0>�MhT�oTb"-o����O�������x<�|�z�^���ϥ���*PG�Y(o6�~|�S"���3ݞy�Ś�U1r�n�$��*$;Qm���u�����֎���)G�fdP�@��\(���94�AT��ܚ�ί�5ľ�5��ޒ�����=��b��&VL��0�I����5WB������ҵ�_忌��(}��Ϋj���a�p����8�Cj��a��}��7�:x� M�X/��!��{�ڇ���A����@��'�:��wQ���vBe��%��R�}f�Y	>h���+^��0 #��"�H�� �;=�)���)�	��Xp� �%؉��[LՂ�����@{�܇��v�0���6�i���"\��}�E	�83�j�El������3Ɋ�]:�$���_��k�U-����2�0�#T&��Dp2��&�:b��ߛTdj���tj��H,�w�JC�P�a��[m�P����)���agq%*$^�贗��2�<��
�AW�d������&�<"iZ
#i(�d�� >���i>�UT2��M,h �0rt=/| ���nk8c@�q���`�0�n����6��y��9�Mn0��e4-f���<�i�� �/𠜏��A|%
�Zfs��o:�h�	�v`��( :�I�ѕ�������� ���Oy�Bi��jT��,h���;�]Ɖ�l2I#6�V��D��i�Fo$b�t0N�5g5�6�z���P�.�O,rlV�_��\��^��,��|!v5���s�<%\wP@��ZH|w��z����}x]�����7Ƣ,
�܇J�1�Ҭ�#w�,){����A,� �v����k�żDa��l��M�Zp#���&w��KD73t�4&�3.'"(Cp�u�im�Z�\v��u�k��,+�/njC�����$rZ/.R]�����g#��6���H8oE^*���s��g�"��!��)h���"� |�I$G��@�D4�b�ʋ�ٰ�ԝ�u^7��b/N�x~+2�)���J�Vq!UR�I>�ŝ<�����'ڮ�y�	��*[#-+W�:���D'��k����nfA	�|�g�������Y�ol�t�^��QJϏ�t%�V�"�~d����Ѱr��� ��j���S|�C��^�~;����֔p^,3��Bh�!#�2 .!Ȝ�}C��c����<GxN(4��\.Գ�I��3�I��k����qA��g�~���>D�r�Vپ:_��T�]T�+�l����$�#�HA�^:<<)�G��I]bJ�Q�����4�wEI����fis��I��`/���6�f����N)���_�?�^4�+� D��E��Y1��1�5������'(� ���k�؀<�C���6�R�)ф�>����)a��Dח�O$�i�d��v	2�PJB0��8��ej���f	�n� �2��<��	��}��G:�9U���c�B�~�I��@��x2�_N�A0��_��=V��6p�N�z��#��?�����cu���w)L���x������͇5���C[�I{*.U3`>@c<��~��&�+h�����eQ��srjO�f�٬��EH��D�!��ф}��:�2V�"&��th2q��c꛷���F[�tD��������d-0���a"��F!y�ŽNO�hra������Sy�d��6������ ����Mo����V�6 ��i�G�����/Alkr��d��.��+�~-%�AN��q�_���^2p9�IV�yHD	4�@�S�1GdM��0��Z{V�$��;��M
]dQV���R١�])K��N�|�'ߛw��%�Y�rZ1���-b�ٱy5�����fV�%��tn�,��h�ZR����Ǟ�t^����O�ҠR��baC�42KL(���gTh$f6
	 �'p�:K���ʌB���E.��P�#��ۗ�
E,?Y�o�lP.p	�hB�2<�UX�F(�nvh~�
��:���0�0D�܇���&B��9^�N�G���2؇�����\�F�ύ��F=@ź�`�9�x��w�j��w�������[9r{8\�υ�Ĺ�����&b����HGQ���q���DX�-x�=����RՠW���Iš��d��=:�N�I�� ����U������_��Ϭ�R�k��L`+��-����Q�cp��_���UP�Î��^T�H�آ�=a�@o�E������:8?���U���j`;4�p@�/4���V'O;4C&�|ѡ�9�|^c]�����j��J��|�!Vă��y��H" �8�k�Nd��2B�3]w@��EJ��')h2������/�R�M����:kR�ɍe*Aa�n�oqb.�lQ�`6�6_�_H��l���A���� ���-�`��p~k��ǌ��!�m���=z�B���ж&z`�d�Zb���'�|$��s8G $X���9)6���K�VBɹ��.>����^�=�^���7��	{�^��v�+wu�&Q�S��K`k���:}�8/ߧ�wn�|\���V⵰��F�:T*ٔ�.#�ӓ1z��xzpD�ѝݗ���α��񅜝��5!�l�˃=�J���#ʣ�&�'�rv�/z�ҙ�aB+Y�<0*H��^\x��� m22R�w3�|�b�>?
߫�|q/V�(�kT��ݠ��}�5P����x��H�TjCe��>����9�.T�=�~�/��\`��+�/^���!I���8�{���͑t|���½tt�~��2��E;���k>2��<������KM�Rr�g'4��I����F��fF6�Mj�T���w�Ɲ7��8�tZ��9�Z���|85��(�9�w9q�g!.�ݮ�B�~�F�ߕ1P�F�߃�����3k�ݑM�8<.�	�A�1(b��6X���Fa�����I�ޯ^���r��ݶ�+���k�>�䪄��,�x��Vm4	�1F�M��PuK��-��ؠ=�062z��5�N\J������Ӟ[TEG��l�*�!]	:o|�BO-/2u?�2�V����%V܀��a��l������5K�R��t(Y�{���'�/f���M�؅iN&d�V��@����޲V�Du��Q�� u 
��2^4롳��&�yA����t�Ф�.�4� �����(��?�ߣЁ�a%��K_\`E\�A^f-��F�Ν[��fMf�,��h�P8
�6w"�!Jn��!9ҝ}~w�0D0z���ܸ�¿�w8���(_�q��F�F9����_�����t\㠝��G��߻R�FeR/W��$$�8���$�$��g�1JL/����!�ԕ=\�ZJU���U��h�Fdn�P6����7oɏ~��ŋɅ!'�������ѱ��K�A���1+x6�I�X�t���*ֳ�^3���1э��*�J�����]���ٓ��d/A�fA��R[���=:ܗ��{��0��'��fĆ���=|Hdؑ��=�#ҏ��>��'"�k{`8T�;�T
{n� �G�Hw�7��#����#�~���&:C��{{D�q}a�Zj�G����E]5��uo�eYU�"l���6P���kPKa�@��J�"�T����}�Tԁ���.�!z��q�}�wo����T�T����M�D�6�_��کNܒ��e�j�Ť�ǡ�`y��n�k�UJ.aM[�_rEE@{����]=�*�bT2�J���N=����@����s�<�~����� �}�bSO���ŗ� H|g!XsP��>�KY@
�g<<M���q	[�C:�7����Q�n={�D����Y��2�y�S{r�?յ|
�
5�����P��??:�A�D&�S}�s�4	h%�Ѕu��J�ώO6�����%8|������v�jթ���q����k��D���Ж�{��b�R��-!���SB��wJ�r��)���O�
�L�h��� �7p{����]���s�t8��m���i��#����gx���c��{�@����x�٤�,#;S�р
=�ф�捤Kcp1���Q������j;���������p���Q�ʿ�.^TnB�\V��l�F�)4�������gX[D�/+���nq>Yd�H}a产YM�:�[l�Q���{L�v3��o�HO�Y���!��VMP�PKm�'@�١J׹�)l=���d��zp�����m`�'�V=k6s�5�qd����ـ �n��H1���� >�N���mus������d[�Ϛ�����Q��Y�������E����Rxd��7�@��?F ������p�E1��2��"�̄sL����~���F��ƤP`T���ܖ�v3Y�z��M�q�1�I@^xW��� ��7e3	Q+"�a X*��δ�rvdes�����,J,ېg�*&�i ԣD$�q")yd1s�d���SA����Q�Ͻ�.��Fm=X���mD����0>0J�4x�����A%�<z(�xG?f =��td���3p2����`{5�)T^F�{8��y�Ρ���pN�AU��)�Y*+p���,d0вRc��({t̀��%
(S����,��$R�-|�Ӊ���5�g��9�y���1��������@�h,Q��p'<N =�������c:Y� éLFSy�A�CM �]��\
�v� ���5\�$�qa��HX�	�b�ZZ��u��;��k�q��%~��7�~hҶ{���/��|���H��N���ů����Rԡ�y��,׶;�:�^o
���gE��7�g8��-@/��^oY�9P�T2�w�����n���Ε�f� �k��u<�s�{Q��s
�q� �M����eO��p�+�.D��3�0�s8yxy��1Ծ��$=�I�/�����`.�|�`�L�"7P��f�y���5�1�{ �M
NL�~A	�����)*M��q��g4#�N�GD��)>�k)��I�� � �VX�<�*�W|�5�C?I���{ �{��@ j]�?�� D���	�ӕj����$���|�=�5����/%��^��Փ�ȯuV~�c&71��'�\�vm7TF[D㼚�%�B��}9��Ent�!���k6'�h��� �7#��k�[p
g;j�SC^��%A<��0�e���̽3�rB=������ʼ��R��-vW1��Czy�Ȗ{��{�� ~���a)�ڰ��5@���������w�ޠ�����u��}�ͣ�t-)�+@�=����鮮��~�E���-�k|������� ~��q��˩�N���/��1�aǏ��=`ٜ�f�q>��[o��ـ�$��fC���i ��@j�|j~)�ׄ+2����=�7��L��g�&���QV�<)��d�y�~Ie,�?'�	P�9l�f5�-O!�ء��l�Q"Ӛ�aˬ	��X�Z�*�+�?��ɇ�I;�c𘌧r��W���iϟ<��{��e bj1�o}s����Hf�1�6��c�
S���AU�
 ���c%ס��V�)��z?Җ���8���C�Eq�z�^FrG��$�g����=�]s��AT�ip�$o4�+�ȼy�D�"L')�[��Y�76�ZY��f�ºٗ;�2�P����ɋD�7l����~�\V�]�{�����b�%U]Ľ�5Y��RAK��@��f9UA�I���\&����	ѱ4^Zq�f�������aqg!8Mu��c����.�9�v�i�aa����h�hJ�F9Nc��BC.w��#y��!�W���-��{��A�?ar� ��#p�F%��_i5p��֛����	�=s�뵭��<]4K��
sjq�Q������P���3h�D���M�>��6� �O��=������'4��9+����;~��z Xr�����UF26�� �R	�
��@}���2qJ�/����B+��N��*HPe*<�5�j�[��FbJZ�V�x����kЈ��U�I轆A������H�w��&���}[��L(M�Jٮ:= ���qr��H��ȏ�#}�-56��'�M��/�k�Q�l�#�'����{�u�� �y���t��O~���y����{���r���quWNԆ5�j�C{C��U�<��������c"���D��gbG�'bc:F'���2̔D�W�Fx��
����O�%k�3��;�{!�[�Yr|x,��r��Mټ�#k�r��&*ЄǾ�-h��X�����k(¢Q���
{t�š2��"�˦���*Vw	���#Cv�|(`!PF�k��2��P���P[=�ٚ�6�'��C�YbibӘ4?���0v�Zz�[�w�{<��AKYZe�ס݋��É�鴬W)
��IDG������[� Iq�������q㹇��G�OsE0���?����2=�l$�6����o��X\]��v%Aѣ����F�����BtvvJ{ ��)��f���A� ���X�lX��0�8�@T;M��&wk��fZݯ�'6m���f��Ɍ���1��!)�s��bWV֤$];�X'/�V�`��r��;Dڹ�
:(�*bܼ�U#F>c`I�I�� �63�x��5�gy5@~a4���cY�{��:�<N�ġ�4��B3�IגS�0�:���/$鵊�OU�?�g`����� Y��k�� ߘ^��?�I�?zH>��t9x�.�dpܝ��Ag�N�`���<��� ��{5�'>�9^m��ד���R$��寔�PJi[�˴[�N�&����?���C'�{�wJ���G��*Fjw,�F%�B�z�0Z�dQ6�
ܔ��8740'�&���@� HG�Ĕ>(E�UHB��"):@NR�З� �0�Qe��<T��H��\KX�Nz�� ���~Cw�����W1��р^!��Օ.� .֗Z��}��+&�%i�8W?z���q�S��3H����{u"g�'&���u,`�Vǀ��7�í]�)s���ڈ��b� Ș����+$�[��jȋ	F+oж��j��m���'�*g�.ɸ��fY�,��MyA��彤�ԁ<h��qh�2��~|dp�psnPl�#�Ԑ�t�_˺��חd~��7j �p.wcfu����:�\�S9��r����b֬F-*��"}��Ʀl_Ӏ����qU6��ɒ����Y����o\N}N	�~c��@D�ky5L�mkf�Su��)�,�Ș,g�'&V} E�EJ���ϟ����4J&U�ʝ8�� B4�K
L�_G��ڳ��t7�`'l����$;G����_�=Q�1$C0v(%�qn��{��x��T�Qڄ��k�;��eU�{wJE��Sr2�J_�,Qy��sp�q� �X<(�l'x��/��-�����#�����_B�7�x2RíΪ�CN+ψ�U$8	3�D�F4�Fg"Ƙoip	�f��_.k��Km F�����"G��;>����v�a�RMG�N�#k4~��mM�;wߒ�~��,�����wl��~�:�ey����e��I*-�%p��������z�Ř��b��9�tv<������7�����k��8GC٬��ߥ搻�Pl^��څ��鎨���;��6�����u�J!�[W�R��ѕ?���8>T�[�5:]�� ������,��!�U��@g�˒�	K2f
���)�Y$�cȌ{����Q����b�y�-�(�c���ZQ�
s�B^�P�"T6��ʹ��.S�����ˤ6,�0�z�Yi'�PŽfcą'ؾ�B�W��U�d�>��0Z���y_��^!����{9����e1ゎ���:m$z�R�`�eIuY�e��ք��**;� _lD������Ҿ6H�.u�^���k<��ȈR��z�l�7�r�۝��O�H�(�ԏA^&�T���I��:h�I�[l�G8\�* 63fc�'r@&~J���`6}�;��8�F��a����s�����������e������Ц�4F��x�:�g�����}�k�{��Ѱ��G������|bo)/������{\Ek�j�ENG�g:B��pj��Z�a��dvM�[}^�'VU���^��c ]��m�L^<�'R���\��,��-TZ�7 �c�����j>Kv�]�u�ԥKCoM�F#i-�˘�M� ��&���`İ���;�׌x� 6r�ݎ ��[���l�(��dsL�U�
�s�E��M8��\�&�K��������;��������g~�<��?oT��4��|�h '�����|N[����ͷߕ�+W5��҇";@�x��eUo�I��c�' ��qca4m�����D�gdU1���qI���#�����*4����W����w�Z}ӽ����_l��,�Y3��lH^�j �}c���zS���C�{� Sf��	7vH��G�@��j�g�����1G�K���S���5�xq��[�B�{��H�%Woޑ͵I��4�0��g#���p�C9���2�2Q|/<Xf+#G5#$�td�`�K��5�}���q�Ќ���� ��A���ߌ����Z��xU��r�]����7L�.5�/k����;��w'��`0fx�NO� . w�~l�|\oh�_�z�i�\��Ə�ʢ���9n,�G�X������.y��*��J���,�mFAF�g�T0��hk�uU�ܺ�F�kj�1����������{���/��d�Og�J$Wwv孻x.�Y�o7�\���-dg{����W_�	kLO��*Q:��*�-��t:�D�QΜQvk���q���~w�k��C���T��T�����w���&=����������T�A�%Q\ynNa���5@�I+��k�1��Q��mUa�tlV�{6.���������o�M�b��0���1��2�'���l�hr��y�����_���f��
|�tf�2̆ƛ][%���7���h�~:�0�7VW�N�Uj .����r�!	)�'��B���Ҫ���4�V����3c���0���Ĩ$P"B����8nT'C !�  �&���9�J?s�{�}B>�ū��<��[��F�:y|z"�:f쏬:Էʏ�CP���3d�B���3D�G@���~`Cʸ-�	WP�q��?*�[q�5yV%H���jR[[���PD��2 !
+y 2��X'��w�� 0)�Q�8@*k��!�i	UC|"&+��k�v���h����q,����`Ñ�x��I7����{փ����tG�=(v���Q��.��稸�xW(��q��7(,�~�)�&t�5�#�"U�.Y�k�5,����/�����РB��.s���� (��[7�>���=ڶ)+13RG�e�������"w��	�<{����A%�Q%���Y%��(����a��3M����Q̍�`<�C���f���@����8)J �^�V���|-U��JJJ�%�T����S����~���2�����N�D���ڑ��e�ޓ+��r�Ҕ�����&6�=�$T*�WTa$��>b�ż�צ���t|�R������Hn<~&���'��?�Xr�s0��WTm2��h8��3H�"��k}>��;O*����P_s��<�m�Q�s�A���e�xq��7_����@�x2@��s٬i7V5����ғ�^S�������⯟ʮބ�?���&3)����k'�Zi˝�my��5�5(W㧛hmy� �`�������ܴo��Cy�Ïd��s
j`&���s�B)4��0X�*����cij�l�N�0$���"4Aߩq��ר-�	|-tQ��
�$�"0ccm1�sgCMV����U�7�9j^o��7zp䋌�2R!���ؿ��u���W���gK�]�����3J��g����XG�}��7��R�ťjG�q�#��1�G6v�RZ�4	���ylm���e��TK�<J��!jX�}v62Ȉ�����o�%���G���*=�����Q���f��:��'I-H�]��s��~��r��x��J��c����d���Ұ$�<��0��40� '3�'0�淿��|��"gβ�pzjCO��w��=�#�������=5��g��P�@�����%��T�<ֺ�A����L�|���l�����`��,������[�#�ڀp��<ݓ�j�w_v�ڂ����-��uY��f4�t$�9�r��L�E�v��彀��J�mu}M:hL��j�iH* ��
2�B,��P�ݤ=c��<r�VQ�*g8�fsVX�G\)�W,fo���' ,D�p2PGl5���W���6.��Ãj%��>b�#�c	�9?bAf5��/��S�x���� Pv[���R.��9�6f�)�-k#B?�k;.)�(u?}��IID�yő�`���ui$Ucsn� �)	�B� KĬϊ�s=4v{Mܬ/�|²�8/T�@Y��5�呮���F�Ĳ)���(�?9?۫��� ���(���_x�h���2�xо�j)[�@���zOL��䢫 ��ze��p�a�]��@��'e�� 9�ۄs��=^�v  >E���n�b��=S@�Q�����������+��s�B���
 ��I_o�Ѯd5�x��gύ4���>��T�����w��;�u�9&���.��|�q����k[�Hۃ��{�Fe*TO59�>?�0��\�\>�=��"�|!�b�Fl:=���h�����@ ���b�f�w�)����.ǒ ���^d��8�LX#�������d.]u��-�ԯ�5�wI*W׻��_�3����[�[e_]�Z��Ɨ-r������6�dI����/?������?��ݫ���jW㶚6y���3�lnP�=~�+���(
^���kN��2��-��ꤚ԰���:�p�pzE@�Ka�WT����zl�3�H�)Bw0oLƋ���$�Gr�r�2�w_~*���d�{]:�D:�X�"(��A��׮v�����r���g��F���f�/�}y���j��r������Hv�6���)7e�����g3���F�(��$�Q^��꼊au!��kv�.J(!9����(8�~�̐e8cL���ݾ��i�h��è�N��53��P2-����#)�hܘ�v7�>T���Q�ԫ3R���h|�����Rw�l��������5�q�������K��~�e���.˛h
��Z6�*��VdMY^䷎}�e,�`5D!�SHC&�� T�V����&���\SGs����G�ɧ�o����p����n��h�||F�aL������ܺsS�זy�?D���@�{�����y�**�}R1L��N��l\]3ޛ|F�����M4���|{������'���5nZ�ZFI��<���be�M�Db	2�{�ȍ��+8���Ld�[���Z�^b}&d�$-&G�;�k2��?�s�6o��>��<~�T�5�z�����ߑ��s�q2��7.�way$��~���F�b�R��@r1�v� ��3m����+B���A��U��N[�i�,��z4A���#�-?��^b@U䔿�����9ZK���!ޛ�$�Ќ�"7j��phl͢
WƤ=7qG��d������t؃�I�!��U���>�����Ҿ5��������?��!�N���f�iy��!��j�l0�uP|b)u�=�	tȉz#>�B]�k��A�����l��x�T��� ���Bm��5���p�����S_�{�ȃ���s`;%�RQ��P[U����� ��0\�W�J����/����@�$�ql���'���辤�����Ɵ�k{��]�	�$?��3�=W��$N�4E��d<�����"|��A����������yೡz��Txc+��c�aLe<�TSWmگ�\�!��-�y���F\C$�����s�ǩ]���'�B�%�.�s.�~�����s����	i�ν�cg�T��#^�}Mt���qo$�ؾ¼�j��ѢLh`fb��8Wq`�jz, E�I���v�@1Se)����ip���
:WX�6['2����Ql��@�},���45�Y�����\�^��V,�M]�^�x.Kq*=4�-�\j�׷9���x��sp�j���fE����Æ%?g�����79<ؓ_���*�[������D�4���}���U�;`c���#����_�6��ػ���2�zy�t5c��򶏊W��'��P��`"![�� ~Y��@����V�C�_�Li}%i��G���XL!k�(��]�����fU���S��Voޔ��K�I(�~�%Ki��?��'�~'ўՌ
�U���\�(���u>�ɖb9@e�Q��w݋��Qh0��h~��[�FY#�@�D�����O�HpF��%*䚇A&��Y.s��%���a/���?<��T�K��w�;=ƃ}_�����e�K<�o�h+�Rq���z�������5�K.uHL]�ƛ����tN���o��@��B"���"P�B��?����A�A>�q�]Ϡ��t�A
4��;���׿}.��o~/O�?���/}:���>��,�I�?Ac�5y��<{�Gĸ�5N�ƃ�c��X���3k��ס��hξu�M�7���r�=$�����@:aJf��3e�@��d�t4�����es�4CY\��xh�E��:+�b:2P`4u+��#M��j�b�'gI�s5,驔��>�+x	�4�Obկ�7^�ĚѰ�a(�<ѤD��;�ԙ|u�5�M��\����?��H�A p�a��Iŝˈ�ߗ�	���!Q$q�dF-�� ��ڮn�	`�)h ��\F�e}m�	��??��0��k�c���0C{�Җ�����t�
�UenC�#If�z
�h$�y�3����u*��� ���"
�G�X�,�s� t@Cf�?q��:5QЮ�[�����Aq߭oƮ�;�(pӃ\&�Rl�o6B����Ć٧u0�<w$2��5��&!x���`��IЂP�L�A��+:	j/�i��A�I^��W\�5$d� �����rT4R+�O�S7�yi��N)+f����&��3��H0����/P����eU�N.m���<��E���0*��qDT�a���:l4Q��_���9>5���A!���w���W����8�X*����{�s����m�IY����]}����AmA� �=�������v���F��@�j�Ih8v�ʪ���yN�W�=�@�t:LI#���G3̇�A�qR]�z��#�/e ���zPn�b��l·]`���	bS����{^�"� ��a	gn��W��j�g:����d��s騱�-kL�1���ҙ��Օ۬D4I훰(���,W7���D��$�kW@S{�ku�)�g�wp�	X� بi����y��;�Rt�v���~�c��g��;o�G�y�I�գ��$ 
 ��V��8�A���e�(/����w9�}5D�lBt�"8D�s/^���ٰ��Q�o�T�k 08�����_}!��}A�akuI6W{�Ԅ㿐����cm;Tx�C֏N�k7�J��C^4(����g�	����Hz��5��l����f������I����-�=�"`�E�7�d6Ik�-�gKX�9\�TEb�p��G\�8
�޲߼2������[�o�y�w����n�]�%��,��6�_�w^����G��;�ݑ��,�}���`�҃�`��yp��q�P8����	�L.�Ze���(e�PG��x��#A���r 6X>�8]����z�M"Xf�B�F�G!x��aN֟����l�➦@�U�`Tm�&!�	����c��޻�P^���dI��D ʚNsYR��<}-�nܔ�+D����+�x�u3[Ub}{G>�ئJfN(H�i�E�n��)Q)�/�� mg`�YT�@��ژŔ�q�4�LP�hvWx�P�(��6ey}I͌�&%�`��Lr�X��@��̽�?.��PT	Z*	�<�̸��r"P��G��>%V��$GQ�0p��@V�l����]����I�z�rp|��i��ĩ�L�r�C2=��u}�v�)�����m{���gAk(3c]@�E����w�[K�.3�F�^-2k	%pPh�zh��r9D��c�DY�c8�;��'�rV`IEJ蠌�?E@�sS�@��	$�Ì�W�62;6[#���s�`�+x���9qO�\ր*ZT����U=$@PF��qš5t%  ��IDATBb�Ǝߓ2&f�MF��0��C�/�\��n�=V��)��k�;� 1�q��*�*J� MTY$��"��>1`�Q�lvI��N(1�H님T�y(�[�l�t�1t-3���c�Yѱ�`�g}GzXY��CU*��Y vI��2����;�9ϫ�h`u]t @���˲i�Y�%��{��UQ�ݞ;�h<��1�mT%��#H���Q g�]��.S�c�K޾��@�Qm]I��(D�S곳Ѿ�o�7�z�d�DR~���"�(>�v����FG����\iR� �V�M� �S�&��Y���������%�ߘz�h0b7�k��I�~2qڳ�2��5�CG��ب�i4+�|T.3B���{�:I��K�f6>{L����[P|��嚐ʞ��K�sR�|�*(РϬ@�A��'����o�pE�s���I{kUV�6Y��r��7�?��T�W�[��z�_kK��A= �Ã���ŁD'�`\`p���G�i ?������������Ҧ���Y@B#.)��]�c��G������T�"����pe�wE�y���̞���(���2{O��u��>��?�D�'G�����J"W6V�����!pV9��A�
�T9b}�F�%K��C��N�M����#���|�Ь��K�]�q<�;�/?�7�/~���9(FOs 1Q3v`gYX��c�������k�gm�j�9��鄳�8���/�q�}�06.T=���C����Ntp�� �c+���B�87bQq�=���#��ڹޘ����s�ȁa��+-8R��I7���}G�ˁX"%"�HF��T_���f��_G�]���'��<+'Ăw�B�sZT�x/��{��r�xlQ%���k�%��ߛ�d�i`w���x�--�рb&?��W��O?�}�5�C�[��zoMfS��|C�����\'�u��/��𢯷[�a�'[��l�՟�I+	h�+�P�,J8�Ͳ�`H�r^LL����K�@�����$���������&�1�¨�BԵ�Y�t���a��/�L�C�k���KF�^���7���߁��ղ"��	+�6=,0�AS5�6�v���$?��/��� �,;��=�*>}�	���-�|pM��u���n@t!�z��BF�#�v��`��h>g/Ean������{��;�{���Z��1�t845���u�z"tD�&&��*!��Z��n��Mr�o��� ���&3I��exQ�t��e�&HZ�^��t/�5�u�Ďh!�vW��h�H}��R�� u�XC��bJlg��yY���='��>8��x�+��B��3�1Y�x�3�,���bT�p{Ҡ��lUƜ��X]	}��6�%T�kv��Q�W��,/�;�<hy7��B�zP��_���*��
BP�V�֙�#��^��}4
&;.?�96kr8'���v�]z�^�^�{��>�M�m��⺃���@�T��W�_�"Z8]�N��y�v! F�%+��h|Gs�O�v� ���q,n�b��;~���*��t�y����z���#p >j5��[�uV^;������v�z��k㟇c@��4&���7n�\��^.<��#T��M�kB�6j�4'eϨ{�	1U��6sxBLZ������'=K���&�ӌ�"��N�$�/2�Ɠ_�$�wi�Z�� R�L��������72|�L��H>��J'���%k2����3,��
��ѡ�1��on���Z�NOMtf�;�fh��E���E?&��N�'��gQ�ݕ�B�j�昋�Q�=OC|�����5����Qt��9g��.�5���9ͼ�N����@GsD*�2� vfyc]D-ħ�P����k�t���<��;IGcT�eCԚ^�uh��Kr���l�6M�iRU��0t%�d��D=�^�5}��7o�εmdO�>���S�y�m��9�8������c���O�z�����1������!���o7"��n\�� ACR�Z�fC d��`�����s��'	u����q7Bv����1}�у�O�ȣ����E'1�_^j�{X���� �K�w�fp��ݝg݀�}P&����K�g���z�@C�_O ��]7��Q��>ϕf�$���7lj
����\�3�����D:�3���X����ņ"�D��M�������i�I�)��M{{����W����+�M��ڃ/��8�aG�|����;�9�'���e�{��9'.Bu����� �����ϟʭ;w5��H�$8"t���$B���G�{�ƊGn��~����
�yd���=a���M���ʚsh�5�uY�D���9���=f�L|��$8+�L�����Y�

��2�̽�9lF�5���(�"X�4�K����c9���D�伯��	�����&���yұvV༄��8�!K��W:Fl|{�a	�9�t����&��j�Fj�(ѩ�_�$*W1�M��1G��z��2��}�F�z��x��Ϙ��~�.͸I�6��ؖ���u;T$V�N�����J��U���1�dk�F�.zP� Z�������ދep�}�>s��r��$�����q"���s�N�6-ܻ�1�6d*5my��P/%z����$��]��&Ƙ��}����`Χ��R�r ���e#�����n��A�yЏ���xbT2�z=�e�\QՆ\a�!c��7���;;'�Z����D��p��3N�vT
����g�R5p�����#�%�d"�*]՚�lr�9��ݝ��1�������5��$�uW�V�3!������TV��m�U���}.�?�%)[��bd����p���nih�~>6`ƚyAEE�� 6g}�i�a=���D�W,S&���{��26�����@�"�z{޼�C�������~ ؆�\�1�;�Y�9|���X� ��?��_��_��_��7���$��-����u63���*��O�/ؖ�y�Z|F���ږ��&���,ט���N낳��h���X��.b����k̄����>���Ą���4�ġ�������$w`=0>r�F��^6r.�� PAm�od�B�z��U�Є���K�jAV!�{u!O|H)��Z�d�_={L5�r�&�N������a�!���z��+�a��~��i<��k�����]��g`��dܗѤ'���F$;ˣ��d�)����e��!�Wc�g�Bz��K�8��n�*C�}�[.J����؍���3���R�����'�?���&�:^J�PN@�2h3k+5ꊢ����rvt(+j`��7kU��=\����y���M�� �����1���X���[���qU$/����\��=5�@�WL.�'�n[�|��Q�oޣZ�(1�i��44��܍/꧒��zN1x���$Y��ˏ"���i�.�ڑ#�a�M1��!xG9n{{G�鈓Z#6Gy�:�7"�IÛ�x��@9oX=R�˂~}�iV�  xc������׿�2��no$=��9�XNF<���<�'~��F�a�=�h�!��P���n�s(�s$��
]	/f�Qܠ&8S7��}3��֔Zp�구2@��&����c�h(7� C�j��4�+�U�L�&N������\kl�065��kP|tv)��>�� ��F�ج�W�j�L���'�59�l���?�CbH�(���;�1p̀&DV]�+��K�{� ,[ ��f��Y�Թ�
"tdA�IHi6^�\��h�D4�L*-
�9~K�����5 ����A�^�o��$�����.BI27!yEL����sDB��zY���Pq(�Pzq��Ej�V1Z�U��D���a�ә�b7G���)w��Q�T7!��h-Hdp����	�Sʦ�,�R�w~yA�2 ��]ϰ���A��۶@	�.��{ě~PnJE�A >��eWH,SWf��+H�)(L4�a�ՔM��~�I	)�n^���|��t���DM�"9  �Ͱ�*���B>��������	i!`0c4�b���~�/�z)Df����)HH-Kb��Y�/������p�ŉ�,�C0��r�����ӹ٠Dʲ�R<M��i�G*=^�$l���Z>X�Gb����I�i�Af�}0>���1�M�4�~�M��0�|E4O��?�ͮy���牀7�w��]�*������7�4��s�s���~(>�լ�<ص�|���_�)ʵ�[��޿�.q���6�xǭO�RަD����0i�[n�6W~���t�%b�2�Ŕ�L, &͏ ��ψH30��kR^�l���r.��~������� 1435���J�f��q�*�:�\��]_�2��LY�-�}iTԏ�����hԽbwS�ڭ��7Ci��C��X[���@�4	랆�.U+���Sl�F���E�y4�$�s&�^[Fj�u��w4��3K��㘌�5�(G~�:�O���۲w�"U�nbT^g���*ˉQ����/?��n��@�')4�b�Ǝ�������3h���˜��@��1�dm�އ�4�A8��^�x.���NN_I�cO��X) �~��+�=���FQ..�9H�׹rrM����f<4{PP&�7�l��!)��d���!#D	C�Ռ/ts��'�S'�.���Bܯ�ب�ŋ��؉q*�f0Q���(ـ?�<�G\��E8od�F��\��M���� b{k��0G�o���Ws颱�|�\sNy�\��0]gԖ�F���������l�z�ˎ#O��������rY��:3�t94J� ��wry��	���]g����8�.��j`)/3_#؜0Vj`�j�K�PB��/(HSv5�xs~&C��V�(
�%LMk��~_E7&���N92��
)/_���:0��^�-��j���g�op!���&v]�c�#h8ow���ԐN	:3�`ʭ�B`RcA���Lԝ��k�m'���>�	���<�%�պ)9ٸ�a�q��\ψoJ��h���rl���w� ���ȆոQ�=��A3 �c��issFN��9h��HI�	m�2��2��vOL��Q+ekؔ���bb��gT9����伄jU��ڞ^��ޏ��U���}���o$7�E\3*v�q$&	���7�ҡq�k �lSC'����ޒO�	�:D8VfF���5�=�� �Y*��������˓C:k$d���,(L�ρ���(Y�K�Mͦ<��d�
,U
�Q@��q�Z	M�e�dGq�fD�C���w0���	�@���B���f��څm@b5sHv�}UD)���]V�;&��E��04�6���SAlTnĽ��X�m�!k��'�2�\���h6x� �{�N������HV�ʞ����l���z>����S�;���Z�͠��o'�K{2�|����{��� $�Dѝ"�ڡ�����#�����TŬ��|lm�����-�o^	-�˹�����s]�yO�����%� �d �z1�����VG�j�t�{s�,�5 �6u����yJ��5YQ?��}�����V���U�{�3�`�!�����ռ�Q��u	�+��0����/B�X�h�C������GTT*��I6�ϸpy��������Z���!����~�%'�^ɸߕ�jA��:�O�ݔ���/̧_@4 �}��_R*��+L�� G!ΰyfS|��\�ϥ�o˰7��ZUmS([z=��sq��{�*�.Fŭ�P��&y�H�;�	iT
���|^8$u��0���W��$����I����e�zI���w惡0\�7�	�y��M�1�!�šDk���|���?�&� {U/F�q��1N���}��i�Ӌ�Ne�Q	��@0-��M:eÔ0h
>���6�W�ϻwnq���F��ǚ�����V4����y�/G�^�ٝ�hn������פ
C �Ϊ$[T4B�j(�3��M�C�$ ��m�nb����W-މ,,��Qm8Z�>��Ư�1� ����.�;BNVoY�%��4�e��ߗG)�F|��{����rоl�=����7ot��#�ȣ�Y�X�d�d�,.���,�De?pH�i��\]{|�V�k�����3iv�]� ��BC����9X�GH4�WWjx:��'RA�c�T0.=D�u6��J�A�z�I���A�B}!�m����?��h�ʒ��Dn���s�L�+���.��S���!hxE���֣��? r��E�[��i譍U'��7�Ǯ�d	NY���h��(2�$�0���ݹÍ���#\\�Qa�YL4�"���&�P�2a�Q|&^+9�˂&� �6�ӧ���:����rc�I/�
ޫo��h�H=�Č��C��&�V��o�oo�������kwr�Q[h�(���:�J1����U�C�q}ⱬ�Ԥ���k�aD�����.��B�h 	�ɐ˱k�.;zR	���t���� b����SV.�"9�Z)���eD���e��bc��hO�{_n��E����ね��_�ҽ����/I��=YF�c�0�$��1�c�Vt�*]���mI Z��"
N	2*XH��.��ۍ�&�h�	��g7,L��,�iξy�y�q�%��~��yH\��p����!�"a�f�Z?�+��x�f?$\�����of@����D#{��KX�XB�6?lH���Ѿ�j�������/�=�#���}����Yyյ�������j� *<�U��s���y�k'oOgЯ{>��T㔳�y��<z���4��s�=�g5�������d��@�'r|rd��2�E�,�����t߁g
@�4u�4�ù��yO �2�<xL��=t �@�A%���1��N1����65p��w���s���_t.�ţ�~�����߻#��ߒ�7�\���!ah2��.�����a��bV��zjSGWrqyƊB:�`�@=M����ˇ|,�{��^�n?҄	~9f�P��}9>|#�'R_���+�Ȩ��Vt��]�h!�|g �DS����H�	Q��C`��L"�.�w=�u|&6��1��Ǉ��n�$T��К�ui�ʲڬ���ڴT��Kr��=Q�7�L��X�x7��=��)��f�"��u����y��c.��^t4G��^����+�y�:�M&��9�ZA�Ꜷ���OM,���D�g��dД��$ck2��f(��{��?��}"�r8����q"�$���M�(���x��~�#�o�)F�y=��G��ˊ���������2}�� ~�p���y
�r�r����������)#��@��~X�d>�Q��:x����4�!J(w%��;�e�3xj��t��5c���'S�@3Z|������3�Z�����9�E���)���/@.�"P,!��0��ɩ�~�B:�6�}>�;?��@�����Z�Ϯ���!ˀ���@��ug=����x��bX��/Z�62�lb�Z	��ck��WHZY �����d�{m�@���Ls��+@�׋� ����5���s�)�9��\k3��]���qjD�S%!���k�v�t���_|���:��hMv-ݳ(���W�L�}]�^#Y�5���[DغCۻ��y�N���TḼ<���g�q`-����ۥE)���ȕ�KȤᵿ���<�?���jﺮ�i,G�/��k-�s�g�O�J`��X�[;���?ecgW��r�c����"�������kV��R�2k��+l���o~Eśa�KU��pJ�&�Ǻơ,v��/I��ۨ��7Hun�t��ea�SO���������]������\�O��|#''����2�W9�|[�%�2�/�\Q�+�s���L��煨'��>�D�����D��&�!y�A�Tq�4�Ѐ}0�ϋ�Za�S�?��h�F9C�lP��mg�n.��`�}U���V�s�oL�����|߿{�6t���_t@H\���Q��W���W�=�쥋�����vޟx=�e��O_�ߓ��ّ(�<��?�:����ct��P��"�d�?�`i�N"uq�qC������WW�
	�*�4������fU|_������!�T�^"uJ�-7�����{�JF	�MvH����>VϜ,��#��ӑɝb��V���]���aEc,�[����(�TQ�D!^)"��h����q�%��[,�2�C�����<{�P��H6�;niR�
��֚tZ�6�c�P��'el\.��'����J�����֒j�q�JCc�j]z�^�s����h�Ѧ���{5��9tw�^$ �g��wK��rE�ET+׳uT��Nӭ�
g`��ti��3����L�1����S�w�$��d���sM�p:c�N��ɥ<{��M�z1`���l��K؀U+�t�	�:뇔Ko��2Ĕ��0���;�Y"L�	�ד�J}��جZ��誏�i����X6�Df�8b��P��@6���T���nje�ǄƄJ6��ϔ1����g%�xf�64�>���gg�,�d������\�i�Z���eҼQZ.a�q_�]	�2�}E�#����s��u�󗓆�w-7���v���NL��Qp6_|�� �%��|��2�3p��5h�ָ�~pt��$��TcQ5���s��0:@F�8"ú�Z	����ao0���ʪT4(Q�`,SM2�T4��������9���Mt�4 �OZ�'�Iǧǎ�+�` �
��	g��p�
AC�
�3���S���*c�Ell�8��t^2܄ͬD�m��84�c��Wž�8������9 �g�F��k�D,->��"Ҍ���͑s�,׻��F�T�o������R���5B�c���{w58+��q�m�^[�����P��N����RknȎ:�O���>�X�bM�<}$j��ij ���o�ۯ�b �����B� �0��ڗF[���Lb�/�~��>���-=$�p$m8���lO�ӎ�Ta�-gkZE�S$x�1��4��z����;6ЪHm%F�'�U�z#il7	a_�&��Ur�i�
6o☰n ��..:c4�.�,0�Gb:�{��ۖ��1x�YbA�bT�JU���Skb��T(s_�.�J�ۀ4)b-�B@��`f]�������w�@�D;�u�ˆ�GW�O��o�싿1�FO�ET�gH���&�(=,�#�]�����f���΃w^���1<����-���x]����V�N�B(����䠢�u�&C̭)�WB|��G���x��s<���x>���o,E��`���������c���r�������<����^i����������5���N)���&WAH�rSU��Z�W�SjQ��{�y�g�����+t��x/�*!�iү�ܱ'�=J�`>1�Y(\y�<	�Ւ��Iaj% ��z9y�B���0_�ؠjssKk�Rտ�)9;�)���R����\��������I/O���vgC�h�ۘN�Id�6J�k�@���Jc� ��+s�Y"�w��CI��e4K��&��3eu��:�K6�~��܃�5��+����H^]�d�d�!���O���j��U�L�I��LCdh��\�4�������ŎC��Zj�ru���� ���ZT��^���R�`�&ra ��hƔ��^1t��-����\���̪�ƨD�;��]c�L.5+��>�&&g]�d����GSͲ4#�,���H�W���CeyQ��\�O��40
�"J%��Dkv:!*����C?\7/��"qF05cF�Y���2\�8��o6.�7���nL���g�����r�7�y�����<�p��x�s���ۿ��\G�Y~��_�Cok�A7xЏ�4���Q��q�a�G�4+����6c��C�!�_޽}����b�Ʀ3�e�&By�Gg	��%@)��Ze)�ZnZ̷J�G~h]��媮�Y� �Q�m�\_�&8-�lJ�9�>p���q�9~4�W灁[[m��&�M}�P���&�(��I��ז#�� Ɉ���?2P#�U��H@���!�����[R�&����c������ڸ��K�,@I�{�)��v�+��-�>�8��N�����I���7�a��lS;?�z���&5��zc��!�ګ}z�՗�ȳOy�|�|��������/�����{�$�~���8��DmJ�1�t��&<�'\K�{��<����T�0��hv�zr�<�G)���A���bWPB�K���5��WoX�נ����f��e!�߅N\��gl�Q�
/p��9bK��ت�h֎ؤ�O@�Z�9��1�E	��58|��A����t�'�1�����Ԉp<����-��0	@"~�sX	')�T�	���/�I;�(�`:����g�N�sub�fccSVWJ�ʈQ�(k�T�:����6U'�`h�������Ar�f��{�:8�=O##q�qҗ~�/H"�.E������s��m;���7�� ��?�)���>F♧��|�������B��ṕN���nx��J~/��������A���򍹙�O���[�x�׿���G�q��U6�T�ʁ�V��h�E�aI$�dR�)%�~�=�^��
�+w/�X<g��?'7t�`���D��Jn��\b(C����VM���
� *NajL���/���'�:;&P�=o�/�G֛k�s��ݹ'�K�*:Ot�` ��d�����S�}d���}�8;U�TT�֐��u��^���7������,�¥�Z�����+$��H0Ў�$�I�����Dm�[����ŝN"+kM�����ᑣE��~�7���X"�nGڗ��{��q�dh�>;��:�kt���Ś0�u�w�i4��z�f-u�(h�x:�XS�������?%�r���;:11���A�Ǻ����y���Hsх�t�#r�j4�I����&[���H�!2�Xl�48�i��G�<(�`W#�H�ڪ����Fij�ߒãcwȊ& ��p�� 5�Q�8�A�q�H��S
�(i����2��k���p1���gu����+��$��Q�oZ�`(�~v���j����@1H��ή:�y��J��KMF�6.9)d���h��_D_�>���y��u��S`~*�_N*������q������mź "z�.� @��"�)�+L�p A�q�b� ;�F�R�ɍ������w ��tU���p�к�"���%o����um#�*^�������?�+M�&z�k��5���*�����m�n��ph��)ц�wsύ}��c6h�!W@z���H`)�
=�zU�W��}6��y$&�X��8�Q4hA)�%1W��P*$��K�A��Θ޶���MPMH���/�{{�i~��ۑ���\s���5H���4{��d��A�Z3��ǷD��%��:A,(�*�	ܻd.rk˕�
d�K<�jG���I*CL� T�z���z�D}�=�֪�}��&e5yp綼x�/���_Q	����
��8��K�7�v�@�j�^;)XCYќv4�w�=�ڐ������mh��G�	���u�C�H�PR*oP���ʓ/�;�H��I]X04	6�%Ek,�s(=�k
��[B��)ě��M(e	��4V�92P5���W��r�+�<fF�4i^����5�z�o_��M~��"�>�mBw6	�`�
�Q9E�	�_�H��F�*V���8�� *̕j����#���c ���Tf>�Ƶ���+@� ��Q���=��4���15A"��<�}KG{!�^Dݳ����@R�����33�,0IOkHv���th끡�ٞ�;~�葬6��m�њ�<���
?�=^Z���A��}0�Q���=��m�^���Z|k>9�Se��r*ly�L�WyJf������Z��w���s�'��ijf��9HO�����S��ڲ�AQ�jC����� ���i�kT9��L	�@�6���4�Ƭ��|���!�#�$=��5M��m�T���:����+�I��^ؑ�1�zp����6P����'�K��◲����J�N �^cSXu�I�����tfT�Z��i]ʺ�#�i���L�)�/�ñ��$;������C���3Yd��=J�gj�$���H��{����ϭ��H���}e�e���+�#gc ���{lM���"B=�$���XgSuK�E�4�z0��Jź\�hC"7)�vL9Wn�#X��mJz=fh�yM4�)�Sr�`�#��
Ԋ.�����+Dc�ںEE����j�G� ��rb�2#��0��]�_��+h�4}5֘�XS'9n��hPd��x��#���lo�yK3�Q�7���A�f_ͦfo݁�P�-rN�K�TWāU�>H#��룧���#� �I�� �"��{�8lq�fo4� �S<�Da��lɆ����l,��STI�L2=������u��n����p@��d���Q� 6�)��R���f���0��`?�Rp��;<���>i�.��'��==�S�}L�V?:˽q���Y"ZX�nR�ZI3���ǿ�-͢���y����!"��Y�ާ�t`��Ӊ�x��#膼����M"�?�=�I��gE���|�:�
{!fI���S�~�΍}��?�N�w�IG��o�]�h��O��?�ߕ�J����b�	n���s������٪�K��&�C� ���7���ܗW��q���/���)�Q���9�ׂ6 �>��K_U�WV#�>����?���3t���XU��ǢC���`��`jk�������C��?�^�G�~�*��AF,�Nc7���s�1�/ˏEN�����-F3HjA���A�R<_`_����ߔl�H?>\2'�VZ�������R���iL "cR��:k�DĹ�OAV�~���>i�O6Ն]t:��)����Mu65&��e
������O�έ��� (��z}��ǈ�P��\j�~�c��v�/�Bg����[�;t�kz���'R�i_�`�;^ ɏ�?S��g��;�0�D@�k�sF��3��6b-��0?��HPg�i�^Kc����S�ڌ�ܖC^3���a�鏠������:<c�'�WC�0(,�Ow�Ł�:#�g�V%5ҐEH�jR�b�XT@o�c�p��]_���w�������B�8{dlʐ�#QX����9�  ��=�%�V_�d=Ǵ�p뚨hB��ZuUٔ����3%�C�ۯ��ܔa{��A����&�fB�^R8�AZ9=��Ն������<��'��h��^�}L\?�	%ɒk��� G��%���+���鷋��/�~�A~�컙�ݶ�\�=K3��ჴ��,C��͢�s���Cy��2'&���d%K@���Mk�O�['^��!�M�c���/6k#�]ER). ��~>Јы4�쳹�u�Ω�A���>T۱&���g7�O�kbb���1�����sՓ
�hS��
g������	)(��`��� �p���t���dR����ӓSy��G���5��5k��!�
�U�fIQ�Nf�x�{�.�7ns�FU���|G�$&�d]�b��5:���3"�]���+�2����:��r~�FZ��	%��j��G�����V������ڭ�\�}����؞�ރ�*��͸O�m��>A�8)3����k�h�@ϰD/`׳�>�>:� b��5�y�$���e������S��"sla ^��ZӼ,۲<[h�{9Pc�� 0B|<�����j��� ���9Р�*�{����C.թfX��XlRd�*dc���U�,��bV4�D�2=�PY��i��)H�s�������V��Kp���m�6�h,&
�a!3xj0��Z��ţ����o����}�!0�1,T� Qrj4Q�������a6��5Ap����Y�5M�ۮ}c�"�����y�ڹj���~-�Rr�#W��sj3d+̥���
IV����?���{��Š�����ϗ�`A���#QD50i�]r��4�̯�DR?��C���}��7�n����׻�h�BS��6VV%��2`�<���`D4-��#�g����t{W4��Ɗ4�6�#����dء���,�*;���}����x�hձţ�TtM4t��~%ߝ�f��8N^�s�5_�o��g���vw��_}.;�ى���F��׿���w�^���C*����b�T!�8��U��o~-�}��������g�YØ"�O{mH��G1��{� �h�:Y�+Q��H����Mf��d����Bv�#�6���5��~ì�54D1�#�k���J�����W�|-��rkҗ�c:_a��t[��>�L�*����ڿz�Bm�L��4��H�B5����Q#�D\s�R��k��{w�Ц��f␊Fcy���*v�M��nb�@6�|�F�t�xڒ>�H�g��՗�����Fq�_8~sh���5����jMȤ�b��Mؿ؜�à#9h�G3��J���Vi��6Oc�*W�}�$2KeNÅT @�7�����"����I߶$X��E�X{�VW�k]&��rH�xj�n�"��4q�?y%��s�d[$}a蚘��rJ�
ՌP���%���פ��3��:���M�P?����Y�*�$�LL�͇����;%3]���>'��sU����*6�BE�V����Ցā@v�,�H�	]��Z�Y�i��.�������Q!bE0���47d�+�3�;�6/p���_?�o����+�/������}�t�|���s��8��᮵��79w61J��j��50���V"��� E�S� ʀky�׸�n�6���Z�)c���Y��&�����~j~ENH��zZ@����/,�+2�Hݚ�{&�5�]udz���	Q�D�u�<�	'9�3��:���~�P>,�5�ޕ���S���fsdU~q�F�+ؠ.�*%&� u�!�PmT�)�8ϝ�Y]i�.���z����+0��:ZC��ސ��75�x������%M�������7T�X}u}'H�0Ke��Jgdc���"���aVEN�D/�b���I����[P��,'G0mBߺjڴI��de��_�I�ذ�%���9=9��&.dv@i�M �p�&���4����@����Srm�+��R6�.�|=�<�� d��֕�&�8+��l�ޔ�<��`:h8��4�Q���v�M�:��/�p1X�m���c���/5xeF��p���p(a�`��Jڐ���c�G=3�D�8Z���Kd�I"~	���U_�<y��aՁ���ɞ���%�O�/�u'��4��	s�HO�r�A��y��b~N�Y��,��OS}W��v�d
�;[r��0�M�C��5�A<���.������ ���7?<��<e����9$�������74ڕӪ�
��ԣ�N5��Xb���uYm6Yf��z�a*�^lp�$]���.��n��k�O�W�k��$\gv��Uc�2~@9{����?��D�h_�Q�\|Haa?A-��MNk�U��vw�Ԙ5dU�ha���Z�:g�О/p�\�znl�F�x��y�����wI�Q�vc���W���"欅�U�|P�$t�����9'��a�f�R�*SU�������s?5H��A��z�s�3��m3���K=���dnv�/�fk7��}��G�LF�3`C������ ���	��W�rK��r��u�\_՟5ٻ�G:K��T��N�i���r�k��{��gEΏ{�M�1mol�̓[DA��vMj� �_�J�3|}���f{��A9�SPu_�..5���Bʲ3��!URlQ��h�"��"w��7u(X(�9h�tcG�
�BO��
3H� 0p�M@L���҆�ep�]�ۜ�(>e�$�y¾#pB_����$�`'�/�X�&E�7w(�x����+.g�\St��SL�����]���-���>�#Cǣ�Q�8EH?x�@���`�%�JG1���z���f~�/*�ͫG��dG\�Q�
U�_�_8FY!!p1P_U;zL(���W��sO��<_
�2�,3�(�%)a�XR2N���'��f%+0*�����,V��}N����u�'����W}��m>��-�����:���d�Qo����jÆfrJp`�Q}d�0�ti�C
�k:��}�y� @���UeB��� ݒ���
�_;� N�O���ɨ19c�[�*��G�8����b!οqҹuM@�P�봸� �i��8�],D���E��ںX.Z�rz~&�զ4T�^� ��gS����\a��x e�8�{#.[�����i�������vf30d1�6�$�׆}X�cb��FO�ጌ�ݽ=K���G5{~���,[>ŵ��*�L���w���������?�d�0��38��w|f�2�ʥ�Ԣ*m,���d��fy3�g/r��IZ������D� �_� A����� ��#Ϻg��>U
<Ẉ��,u���V��V�b��Zg����s��]�R644�&��2c��oX�8v�j�#��7�UnL;q5�1Q>�ԙ��KM60]�է�J��2F9r&��6i��!��	Y-l�������h�B[�3��������XV�������?������7L|А����o�(�������XgxbN�� 9JBi�sY�&o8�U�C�����d�y����B-ɗ6IB��-�|v��}����+ryg@Bp��\8mP��?�L~��?��j�(To,c�j���j�â"D*7vw��~�d����׳�x����ܑ;wo���R�/��{_`�Y�V�h�a�:C<�h�f��=@�߻�f��D���{��Ģ����Q]	�//�\H�v��v䓏�� ��*����6��^���.a���o�"B�߃`˯ ɿ���;���ruy���2��Ѽ�=��?���^ȩ:�V��F:���}`rH��~�~>��!�*A��ǆ��~�e���N�� <X�%9s�تk��N(�W0����tŇ?>����&A��=�z��o��̳���!v�vp�	�'�W�:k���7d�ґ�Q���>é�^ ����kHKw��5����I���6+xHT������ʼ8O��'�F!�J=jw��$o�[�Q�F^��h}(�3A��tu��;�����b2 ��P�`=0
�_���ǹu\W-y/T�T�h����&���öBVwL¤�eD**���H�����6E�'�5&���tap]g�;M
�hx�L@�+��|�����~��9�*�7�2� ���˧����o]��w� 1�b�`���Vߖa�TΏz��8`�^r�b�#�_�S��,���lȄ�L)�*�Ffo�j'�}��ܶ���z����̏I��L��)��u�Ϳ&�����'W!�ټ�߁�8w&�+MRl1��}݉��J%Ʈ����~�"C�q���G���t���= ���S���̂K�f��;���6��P)Ў������2�����u��7���{C&�KM��H1ًv��4�*�yU)UW��	rY�e GH<B�/���L�5N�u�>�wb�E`	�OD04�� �P��k�w���EUEǧ��qܭ0 �`]����YO��֎�ȁ�I��f&���z�x�,�!�}��:��b�����E�����G���o��A���InS��3�GE�'yǞ�L+Qj���nk}M�77��Һ��UjcN�kÀ�D7�H-�:�f�+���M ��Hn$�N{T6(��(��|�_>�ʂ[X5�#�395�Pb�b5�`������Grx�Z� C��^��!�(��}�k6e4�Hc�0Bn��P����0����m��(L��|R4b�m�J����o����oq��|$�n_�?{�F���8K�4��.fʗE��E� *��^�g腣Ҥ��mK���#� i�8y�3<��%&�9�uE�#1B}ko[��{R҄织��� % ���ڂ�Ӓ5  �;�� ��cystl�,4B��&$?��ˍѡ��0���d<���Gߓ+���2�����/���O�|^����_DIP����Vj��Y�Έ�A�����{�@��R1�.�Q
��\d@#U�5����ɟ��w��/��ᇟ���N����7�.��M�Pʅ��No�n��������Id���%���;���d����^���y�����O���lmme-`s�)�u�{R�(�iH����Ǽ\�P��H4�|�"�b��8fN��Y Ʃ���cW"wzǈ��f�?B�{,qCY"�L���σ$(mϟ?�0܃����d}4�ZT&*�jL��^dI����;>� �E��Ly#:�7F�!��\?�y��2J���x��i�{��'e�O��#���WEݫހgx�S[��=R��͟�o(���)��6H�����-!�H�)�@�
��m��#����~��'�¦��W&�[�bjwhvU��`J6dj�>�L�~g�Z��^���ɪi̋�x`�'��x��K�W��
�Pj4(ъ�38�4���%"���y�g�(�g&׃@�W��Ofs����N�����S��Η��U��Q������$�G�d�~�L"վ-��_`F�W��$S��$����u�OǙ|�8}@^p/���r��Gԗ�˻��r �� �'(�*�7%���.Q��R�N�I��뵲�� ������zt����\OGb�2�ޡ����x�W�u�*��3��}T��x'���eŊ�F`����`���\�fUEު�S~+��߇KQ��j�{OFݶ�h�=���T�]�v45�:��P���g4�*!�*U2j�<���I���H�����>)V�OR�������K���s���'�IU�}�Q� U(%��k�����,3���[r��=Vژ!Գ�H�nD����~b�U���񘫟�o%�>���x˚{�V��o���M3�
8h���b��~���x��{��I\u���eEfmSdY�ш�	�T�(��K4ڡ2W���L��&�į�o2�0	F���iP� �uI�����`Jtp<�MV� �j��p�D`%KZXқ�Y�W3�I/sL�]B��~wHJ�R���qCu �����j���6��с�8t���I�!�0���M6*dR`%4d�,	�L_�����ۿ�;��o~�k�����Z��� 4��-�@�������X��3�m�/��rm���"�Azm�.c��gZ<��r���~�_�u�bC@�����������$@���_~��P&A��@<Hm�@��Mn����ߝ\WL�4�Άc���v��KXR�x��G4CϺR.H��Rdw{M��:PcYրy��MEO�D�f�e�>�R�� a��GHH�j�mO�JӠƠI��:�5��oNd0�f� hJ�
5�xbZ��_@_���5�0{;۲�	�ͭ5���۰�0A XA##���G�u���cj�����ȕ��۱I|�Bk$E�B�.��.��V��W�D�&p]���ܺY.���;��}F�04Ծ�9h�1q0��P:qA�?BӮ�(�D�� �m�9����_ȟ��|�'�|,����mj�}_��:a�&�s�N mD �fdh7�v֜V6*tDu��<׵���7���Nh#�g�Q�߲��,�=|��>�@*n��G#���ӭן�ش뭗���Ѡ������Y_C��?1S ��$e" Z&�VԎ���r��|2��<�Ht��&�s�5�3���[QN��m�1O�9�A��`4�G���`�BB �`d�VTG=� ����L�|�����l"�6ŕ�(�S�ɀ�A���xsO/�^7yM���@��\[��ބ�$�G�^� .������{���.4S.=| R�!�:�����ll�ɹ� B���D��Xq4Vg��0$���L�at ҜP��
��%� 4?� ��>)���!�EZ�u������O�?������""�{^7���&,#��7i��c+�J�jҊ6�T�z/��d2	z]9MY��  .P����U�kU����=�B@�8j����A_�~���&�>qp"m�-����`f��^�����Y�~��^�XdskW&w>`����KM�{���)�EU�66)�]jlH�����3p*H�/�93.�%�S�B��i��לT��q��yKN޼��YU�V4�T�ή� �x���kkc���p? ��*[��%�K��@J�\u�jK;��N�ߎ��D�Kf�������c`�z��D�|Ρ))��(�y�X�' ��s$,omq��{��=��us~4Q�8Ǐ��Fw���[�	�N}z�f"���捋�ư��=�[��:���o_v���f��`Q���VQ��\��%�0h�q:��bS]��:��)Cx�Q�L�4P���LM��EIM���!1��T�4��Y9��5�TW�O13u�? �	I��2�hƪ.�_�������䣏>�_���R_Y�gO��e��e.�eem���oI��m� �~�##�^_�Y.[.?��Q�T3�l�� �%����D;uz���7V4��!���&��ã�o_/'j:�H����V���t"��k��dgta��X[��&p�^��'�Yx����y���LW���Ѡ�X_�k_�4^�u.��9��N�F�����c�mꦾN�����z�<�u4���tC��T���<�a.W����Y���� ���4�(lj��s��5h�n�*lLŚ��.om�.?>}� F����t]S��j��R��!����ns�������!�/�_���60��y~�ZX,�[�|���|�J�@�`$'��@�JSGQp%��1��݄� ̐0O��{ٯ�X�P� c6�9����\�.:T��hTSk4���5�Zg�޾�p�	*)�̓������Ҹ�.؀����0�#aE�:�qXTRդ�*��&��'����=�'�vGm�����޸�π��Xo0�� �'��B��<0z?����/!�(��6�UOp���2 A�S��=��[7�e��j��j��Ų��(�&Շ�h�7�M^oC���������z��HDFzM�<}A[��:a�R��jҍ�+�PB}�?4>��%z�)���e�4�[��i�I�,%]g8WNq\`�S࿧ԝ"�M���?|�yqrI���r���M~�&z�м*����a�
q0�-��,P�x}z��&��Rկn47l�����雓��g0�bV�9�5p�"��3���g~ͨ����5�'��-�J��޸�ﱄa�����}������������c~|���#Е�_o(�����w�*U ߺ&�u�;)U	ؘu܈�=�K�}D��ךܷ0�x�&�W/^��F�|''��,�M�������y;��HZ�x���0mx�.x-�2�3���gF��La{4p�ޗ�^�����ֽ���%��u��mJY�4 -z:�����rl V���TP����<���ejӵ�����:�˳H}~���������{RA��V�+L�[�R�s+����p��K �3�����TRL^m�Ʊ':��&NWTA�_B?b�P��~�/��sJݼ����� X�'�{`�.�&����I�<->�L�KJ��l�\�LɅ�Q)��6��PKHU�b���F8:��@q8�@�]}E���5�!h�֊D�Q�4����J���qNlnC������GU��@?�%��z�<>6���#b��{�F�8H<��,.D,iCN���l�s[YYcST�4���A�|����bN'DT(�L4�����OH<lJ�)�@�������C����0@�s���}�������Сx�q�9�PYpZ��
���^�;"�e���w�@�;����W+��ZD'-����h�y���5J<����\��R�I�l�\< nT(F�˨V�ф"b	���� �_���y��nY�C�����ɋ��+��ޔ��ӧz��?�Л�Cܭz���D(HwILc:4%?u���K�j]���6���C5�dJ�L|>�{��Q��_��9qp`O�@k8����!�N������n�����Z_�ɝ;�԰����iV����gp��=* @�
9�_\��9��S~��I��r�%
�p�bT�sޞ�4�.4N�����,�6����z�������#��L����y�fN[M(.�=�ǚ !�*��{�ݓ�|�<���l3��bUQ��'�Ҽx�F�����~!{j��>�

4׋�l����^���cJ<�o�=iBg{6�+M�P�C�x��,#�}�浍W��]� �Nַ6��>鹴��۾����Ī�1ѱ�Ey���Ύ�2��N�G�x�k��k��O?��~�)Sh�l���gl�$������X��f��Sb6�Z�X�B?wbc�3�~َP�A%�u�5�FX�п&��AS�)�/�ip3M"�,��^�5к�  u�F�D@[PG|��-���d��Թ,3M�Z���� 8 ���$$L>�����H��OA!+(����X��9�" ��N���(��,&�o/���ϯ�_�o!��O4RTz��Xʚm%M�5��.|B�+W��񤖂b�{|hdH��@ ��������j�PI
%��g�V`n��0\�*���y�̓_n^��J�l7��3�뗯���4~��{��:%$V��[�ར�t� ӬQa�ꊻ�
�zbx$�0'�.KEc4�#���8uધ!�}y^�Ah�g��r�L�� 5�$��IK��Co��T��DT����%�����*��ơ�S%�JcCnݯ�߾����_��<l��z�E����~�6�R[Y�ض��Ë�J��
ٵN�EŒaHȢ���lh�YW�u*؆���8!4Z�RWt��`O��`
[z���t��l@(3��'z��D������C�s f�����M��+����S���'���~/J��/<���8����-\��S��%��F��?�#�Af���RJ�.����<U#�9?&*G�H�a)��z¸��`����9r�%t�"��M�c��18�U��*�O��]@6���Yݓ͝&u���,�t�=�!ۂ J,3 ��llm3��;>��X@S�R�F슩�t!��ok�G� �HF(�f��Q&2D!uS׼���x���T̨���D�P�Eҍ�P��Ӂ6�Z�?cP���˖����2Ǵѽ�� 1]�P�!D�1eIt:�������V��1�qZlV��y�߻����|=�[��ySu� �F���L�4$n��5�'���!w�GY�篏�ǧ/��I\em[�����UIX��h�B���?�P#�h�؜2��9�����9�DJTk����|��{��rq~�M}vvLt�u�Q�hu��R����44��Xc��;5��������R3�#��<����]�@:l�R٪O�V �hpV��!x~v"-5X�# �́>. �wHA"���RM�T_F$�woސ�ϞJC���7d����g�5a]ˤ�.u��X()Z��w�^Σ=|E���?�����di=f�Ϳ?̢��N�;�ߎ�e��|�w�e�F�l�&i����I���p��+g?z��tzLB��\^BZ�{�b�s���8�Hź&NWr���T����m@TTҵ�V{���H.5���F��b�*+u޳NIߡ���y�44�Au\v�x���ܼ�o�:��pB�V��՚Ӌs�0�f��Ɍ���k��t�^E��VQ�d�>ObGA�6ij��������@��b�`9���0��/��g�4԰X�s}a��>Fq6&kN�@U�g�46����-A�����ya�pC�Q� �?VG|~��H=�� ��ºƄ�fU�@5�j����Ơ(5��y���*U�;�����rr~e����bU��+G&&�+�o��lc��<b�:���\P�G���_p	��ɑWmu]}�P�A�}ecW1��X�)9M��Ǯ
`��R�0�^T�+J��:����r@VI�a]6�w���=e�р%�<ǹ�l��wYr��#"�,�I�r��5�r�?]{�����=o���ܧ6O�h�@�iP��Ҷyb	,�q��9��,W�Im��+��í<�`$@��
�����2C��>Ea��M��:��>���F(��S��0��l�Q�$�ӀB,����.���p%�˂X�&�R�Onߺ/��-ݗ3��#�hv�c�O-�y	c# ���ꀩ���Оgo`b1NB�\����h��`�#W���?ڕM�����T�t�� ޔ�P�.Z��^\(�|��n��^��ǣ�x/�a�s��}_F�	Y�E %6L�J��
`X!��B��c�vJ�����<y�%�;���r(n܌��ԕ�B��ِ���9@�o Vq~�0ㆢ��w d'Xp#�c^�!�Lq�uE���RW��t�<�8A�
mʪ�ӎ�-A2��~�2P�N��Ŝ���C��R3:
�-$��D��)���������
���Oi(q��#�-�((����y �7�˥ݓ^K����S�tlh����Kg�2�Ө�_��Z�;�)]��n�aN��1.ZP �r(pYޘ�^�vtQ=��n�D�vw���?��Mhl�L8A�y@G�1�R/�笑���X�Oޖ��O��8����e�b~u�:.G36��ӭ�Ȝ�!Cv��ܖ;�O���WG���K��H4�lpE�> �E(WX棣g  ���k��ں�U*� �
����k���\��u ��u���j����wem�������.�9"4.t�#Y@֎�XR}`Jd�AS97��0�.ˉ��z4�g��|�R�s���]ť��8&"��3�}��<�81z���u	J�$��b9����޵�� �:'G�2�dws��t$�qB'��u����y�xT�w���t���5��-K��1�b	f��e��;�/��RS�Jc�hX��0\��52�Bd���I��S@ ���EV�� ����l�����vOS&�XJ�eH������_R��պ`e������ۥ�=>?��1��ǣ3!H;>�Е��շ�P�bmc�A?lxM0T�zd>y�D��0��~��IpE��BU�a�"Zh��9d�M��
�iԱ)X��u��:��ᠢv��A�i\�����UR'��̩�L��*���z)�M��YY^\�����ww6ȇ���C�X�����\���Ņ�]q4	�D_u�@>�M���㾜M&F-r��,�3�W�О���`�R�����9��G���77)43���w�,uq���B��2�9]�'��A��4�(h49�D}
���Q�'Aq-[5�M�l�v��ӳ'u�dV��ѿ Ť�duq�3�n�p��c���-6��s��O��#���ڼ�F\�z�9j��?N:7����(�����ª%Pp^O4i��J1��d+U�p_7�~ͤ���p�v���	�8���&i@��S�=[�t �࿳I�TrS�#��R��~25���r#�k��������4)����P2±O�FRҠ��{$l�F�$$5�K�5��Pq����ɥ���u�d��7W�>xqؗ^�,���54�Z������!G���.:�f�,P���O�|<���z�.��w� ���<Mi�7G����Z@`U05FcKJ�|���?a��c@�2���g���lf���B2���t &��F��1��x���%ޮ[춬�sb��I��9��рN����G�2ʧ阓�����E����ì�>�Ō�$�DQP��� �WS:6��I�Kٽ1�)�k[��餎��B� �a�S5lhȸq�j��]�i �wP}0q��L��YbrRIj��8����"��"	ͱ3�0ٜpF�QHB��#D�0�D�Yƀ+=�Wo9d F����l���7��T�.萗��Ba �f����F�i����Nb�$�7��#�� �1�����Y\�ڒ��,��'� S7ָ���ֽr��{��z���<z�Z..ۤ��M^�@|7<�d8�60x�S+�]V~��$NFr^�JX�0�Ն�L�MO���n�3�j@�P=�v�#����Q��{tt(�κ���B2j��H���}���8�c"�;�MO=�$k���d��E��,#���V���ﻹ�+;�[&���"���:&���*+#I��{�	W���[g�m�t��T�,D5L���e0��z��'g�H���G�<rN{��W�� 'o�_�����_ǭ5�]��%�dk��,�ebWR��"[�0D���U"#6<Bo�,_��I8�˳���i��?+AF��~GuM�������� ���99�D������Dۯ^gh(a@�Pa������
v�j3��;���:�VD��##.�_3}u"�N�:��ke��B��e }�zJa{cbh�Y8a�<�0�V����/��<:+8�<6�:WL�na\y�Uo�f+��z�j�-�bS?b`
�x�����SO��{�e�Ihr���B�+���'�v�=a�C̽���׬���!�
��h>F���B���p�YIV��Minճ��{ŭҔ�P�\n�W�1�m�n:��V|�`op�����g�;�ݴ�'��#�G!�-럳������ q�ҹ]g�<�o��p Q&V%ƞ��P���7����f
��s<�5�=ƾKm��?o_�]P��E{a��{�����]�X�p.�<C���-O��x�'Q��B��1�|�"�w������a���lD�E2�'�������&FCEc$L�[�j��jy�����\^�y������ʋ%S�����O�`�~���'����&.nA�7K"�1`+&�c4*@[�|����9$
S�G��F��b��#�ih�� *}mc���j]�`0��oE��u�H���:��w?`�����5���٢��c4� �T=��^���m9�q�� `���#9o��&�>N8`
H|�j��+�W�6ܮ��D�U?�W�j�~��9%9MAK*��s����I��w����5ϱd��5
d�V�%��������#��$��֤�-d&�
c�r�<͠r�r8ڜ�V��ʚ:�
�4�aS�w��7� �� ,6�/ڀ s#��l�4���B�����y��`�&6z~{g�\5"�(��8�扐()�Q��D����������?�Q:�0�A&<#0�(��'�z^|v�š=nSX�qL�9���Ґ��;��k�-pC�]�،�nw�@��ݽʢ��s
�KdJW_��ic�'4 A��k��[=���wXք�ѻʗy�P�Ќ�a$t������t�ޖ�>���lL}��Sy����P���Tl���A0I8�D?R�(fT��	���E쇘�D�3�X�@��A-�擏?��|���im4d[�,G��rttJ�퉮�qb	�očY:��=Nr����@�2��V�����H���?�ZE���ɹ<?=�.�= c����W�i��5פQ?�� �l*#ѥ<�k���9;oy�6'-bB��J�,<�-;�kj@��>�(!�Ze+����p ����E�K����K���s��,� =H��P����:�J\��m�)c�_��PV=�&U�P�K��C4h��锊��,"�,�\���v4D�]��0�P���tc{G~���"���2��HK����;����6��T�ʚ��*�C[WP�B���c����맲�����DuP���|�yU���RC �YŠ̲3������G��c`b�L ��44�R�����S9z�����б� dJ��ľ��{���Qq
F P��n� ,�&��FP�Rb��`�ѓ��_[ۛ�?�@��$��[{���ǂ2?��?J�ȕƱ�|�N��������<�J�0~4*H@�4���$����*V�20��woM#��{���|��sJ��ܔY���ˉU��b ����ݙIDN�,�xaa�I��N&I6���/>P$\�!�Yp����O���B=�?��K�.����O�� �@�[��~�����Շl&@=������Rd@�-y��i������.A������u�>:��_*����U��D2�$�9mT����<E@0���J����٬Rʄ�4������ q���7t�L��� (�#���i�������c���d!ű��%��<`����4Z76Vu��M�0Ю����=9<:�M({�n��;�t�����ͦ��ѿ�����G��~���M^��xF�T+F�]^^��(���z����="'�#A ��=B���~q%����,R��"|����In��_`+u�˜.��-H��d!�ʒ��A�d�
�nv�v�9@����y���8�W��c����%Y��.-P��(c���#B04`� $)�x-���ԥ�(��]�NѸ1%e����IX��Ǥ���W�!�=���=Gz#.�栻:q�`�2�kZ��:�|Q*T��F��l�g 4�-x�204gb��H��&��8>���qQ��x��|lDaf?�fG��{w��p�5sr����r��	�ؚs�S�oc���4�����P���FT�F{�ˢ���P���r`Vp����P|��f��g��4�a��&[�`n��Ͳ&'���xu$�'g��&���Ј�C&�P��k��f(�:��$�ȪF�CA��Hį������CpLl���ޗU��Ɍ��䵠��������	Q]��td��^��q�8�Q��d���@����cY<�%��Dp*�q$O���/��^^�>� }C��b@���i ��;�8W4��<;�۷nP��U���6�ˎ<z��|��7ҽ�@}m�J���4�d|%�R {������3������H�Y��;\�Po�m��y%�Os]G.�v�1������*�S����ޡ�)�;����թ%�샠fw�(6��01�L���9$���n�/�膦h�5��&� ��9���^�ξ��0���m��{�$K,�yx���d&�UWuwu�zF�k�߫��$-�%�h�K꒺�L:�!�$o��F�wĹ�$+�� 	��{ω�c��_�
����z'�������O	�
�~����?�$�������J__�.��]�X��Cq��C��C:%���ci7�Iv�(J��������O�Xc��-���|�{"��]9���d��}Ҷ���!�7�Ug��Y�_�du�d�<��x��]��V/$��/���	%#_��+uv�Izb?:�n��z��%^x9�;7�����5.�{��g'70K���3	|���J�q�����^��}�������X��Vo��0Kr�F� �n�
5�F����"&m����Np�����H%'[%�>?�'�u�54/]62uO�t��bq�)���Ff���
�P8�6|���6}��f�Ƈ!��G鋅?/h��G���X��r��ha�:h��7fs-��ԁ�p#��J�4w�04�O�	��+������u�5F�V�$���&��wt�8���|�p�n�K6O��`���a�k+�� Ӑ�J�M���9s7�C��$s쀉�Y���� E�r�:g^$��e> �GF�{O��M=k�^|'���<�tZZ��zk�V��<Y^Y"������U��CYL
POO4Y?>������	��HҮ�%��3�P��&�c�������8�%]��]�̳�Eeq�f������>�/s9��]	|:㯛|���H���7wy��VQקִ��RL+xI�ϰ O�.ذ����\j�� �+Mw�����S`�y���tbRcTEHmJ�4�[��ZZ��M�1�}VI�BXM��Fb��ᔭ��:̻w�ӕ�	����I*�0Qw_x��{�O1�{��s�#5	2�zMq�I�Jt �U� N����ӱ#L,���%Q�о��7�5zcog�@�]}�?^kr{$�ޑ����Ǐe�����&�G�X�8���Pँ�ȡ]�ľ��ڟ�*x/��_Z��M��E	-?�dpp� ��޹'��JOXB���y��H����(�䴿�D��Vq!�K�#W�q�Xiն)�X����2iB�	�u���-M}�����	D�|d:x�I�A����$���Y1��\_B��6�F��r�@-��O?q�w{s�]$�+���$m9<=���c�^�/�W�J�!������R~��>���#&-@���
W�ˋky/a\1����׌v--�2���t�։"ɷBo�D'��Eԑ��%t�tCZ������C}�,�~I�_��h/���8$^�}.�נ��u�4+촨�����~��@d��$�+�(6U�����pp�(��2)"j@U�SH��G�9����h�k:9=�o��NN�Ϥ��!��M\l�䥽���,�x��b#-�����^Oڦ�'f�O0X�z)ٗ��3 Hز�CfO�ќ�^��T!������+9�����%��AuZ%�������"�����EG��U�0R��W�/���2��9{�`_�q�^
m�	�ᨨn�s9hyH��<�N�x.�7&�QS$�/^��!��sӭ�ba0�������:�8ǒϠ4��̝��V[r=�T.�,����Z�/�.���Գ5�}1���QMi�D.)5nT�s&�5������թk�{����h��H`C�ԛ��M��Ԉf� X��8��H�P��,��?��F�k��%������Qn�������/�UE�\����ӣ����B��Y���rC���c���>:�%g�N'傛}tS�>J�D"���*����+���;�S[�O�~��t��Ё��y�4t��ƯW�Jh�	]wUΘ��f`G�	�3^�c�y�_���ٕ����kF�T��RҸ��W�X\^@'5fE��2ɛ?��Ő�B�D�ؓ�`*k+}J$w:#�᥾͘�SH�dRW�`�WϤ�����P�* D:�+�	��ٓ��28���+(��,��]��$q��s���A  3�X~Q���EeT�ԙ�x�fQ��]H�?���E(	B��)R�'�AyjUk�f7��?�	]he�m-�ņEK
?�D�D��k;TA@����7�� ]��Ħ:�$���C���$�jo����F�yD�}�I�` �	me$�����D1�� !�`ӊހ	"�H�s���Ã6"� ǶjA;�f))@b����R2EX�Q��mR%��rXv�c�E�֙�#�ҜOKos�Z��f��9��!��	�IU��?����=�D��^ y3v��L4Ac+73Ī�b$��ՠWh�.~��rsM����o]G�ß�������ܽ#�0��{���X�ׇ/5y?�i��&�%8�yl�EH'0|c��yR��ZQwCj��=�6�݇ȋ#��v��2�z�c�:1��k���$����M��z*3]�p�$�F�h�H���;���8َ`���� ��4�L�&J'�,��n���2�k����)����i��Oj�~g2�p	�H�G@�>��þ3��5�÷����kR��Vg��|yv*o~~)Ǉl���N�Wruq���&yƆ�P
~xyA�X�?�XW@���5�_+�U�AZ�!nY����Y��������^������h~A�!3.	�%�O�ً��#n��7���rŬ��YZ�C	���B-sC�K���^l�~Ċs�~��n��9k������Khz1v�ꄅJMN����b�wHޡ�N�.�a1�YN
ՁN�?|M���4n Nbߠ@`�?���t�\I�|pAi:��; I�8���#�$:��c�ba��I_��C�0YsC=tN��O<�5شj����a.Gީ��M�8�9�T4�6>��19�ا�� 2��ͭmr�OO��r�y���}#��	mv:�v����t��`X��[YnC���x�`�1��J��k��D�~#�e�_�(c?������� _[��xya:������'��463����qCN�0 �qڨPs�ZX	X��!X1�b��`������e��mZI&��guTZ��F�ʢ�;�6��p�����L���JG3f&��{�]H�;�a��!���$r ��}�| �y�x�a8�Wa�YT]�5�0[w��}r���1]��ԓe�t�RP"s�aE�+�j@D @��=��FY�y�p&s�+%�8���,�B��:�Eцp�°CYq��N���=W뒅�,J�F����~-�N���s�{�B~�Q�|����LϪKYֽ�C ����f�Ї�����L�� 
�����ݸ5��rVF���vGsՉ����8����	ܲ�4�,h�r?o�����s�	����Hp�����]{Q���~9��+��Q5p�O��I�5~P�S�;gI�m�҃�L/ڑ.Pf���<��[]ےg�~!Z����I�Z0(Z�Z�df��&�	,�,wX�&��Gù4FS��WhC�$ �hl�8�p�	�Q�\�0�:�S��J�.��'��J�ۑ�;w����<�.&8���t�{HDM�#f�$�
+_���K��.|�W�(%X_���
C#���$�"G���['1Ld��Ɓ�k�3��y5lJ'm"r0�y�I�GOɝ;�r���l'4������1y�%�U�C�ea����$�&�Q���]9Rzލ�E�:�v{�+���A پ�H�4y���!w���~%G��rz9� 1��>�͟��B�	R\�h��=x9=@�1$�u0C&�6��IGȁ�ｦ4Ԑ�L�Q�AO���7��L�E�Mζ):C�gg0R���'�A���������A>���V�@s��<ʘ`��-�ٳg���'� ��^��{�+D�`������%�N.ɋw]��] 8�n���=�=Dg�����QE���������5�բE�����^����+��0�1A�9��D�1r��=�,K��k��b���:���1��ntqc��	~��#���w�+%Q��F3�WGV�G>���	]�V��Cތ4:�ޔas�R�-� gz����Z�WM��D���"G�K�&&�3��`��H��e��⊾U䷗>��.���(��Ijە$Z&w7��	@��@�/G{�G<-J?��;�!^g�&P���Fr���k� �G�Qn��@�18M�m��P����\")o&0K�L 	AH�	� F2�=tMA�J�Àˈb�T����K�	�!�8�q��>�w��?et||(���F���ӏt�te�V�rps��"���mR��	i(�^ѽ��)qT��� ��A�����	�e����I�k��Ô�ɔ��L�4���J���#٥�9���;�}��5⚦&.��Y!v�b?�C��ޓać���ɲ+�xAP�����@/��5A85ů�cni�f�|��!�XX����>�9uG��bS.�+@�#�俻�x�����'^�sا�)_Ǣ�cl*b1\U�h�i��q�D'�O ��C�t���ݑ'P���DNUs^�{� ��܄*��Y�mM�5�#A��*h��Bu��N�:D���
J� ���Fu�*��΢��!7�A��G�|���\'�F�4�j��f�rqeW,2f��Q�"s�LJ�JN <��Qz�7��Z���S�S$k˲u�|��s9z{�������uoNz�/�JԼ��`lFw(���^8�K�"^�x�c�{��нU���{K�,$�\8����3��wxɔz�����2���`��fl��b��S�0dν.52�[Y�_tbE?#�A�k���MY$��k��O܈��ds´�ȯ�񡨰y�
\on�Tf_/��O~-'��r~2�M`�4��|y��3Y^^�Bb,W��.���܆�g�Z.&����ݻ}��p���̝RKW�o�������L?@��Ԥ�ǚDMtcm=�+�h2��������x��8W���̠lZL)��	��@	��]p*��@�u����s�Ibɩ�`�@D���غ�@��n�����6i���B[��������X*}gry!k�Łs��`�����@>z��ڪ�X^ݐ��&uH21���_���<_�7;
�X�t�+���6�ِ/T�̢��!�&o�hH�g�Z���P���.����H�������@�QL���յ���J��Ȼ�MW*2`�N,��XMRx�j��3��aV�� $�����-͏�ِ�II���Ց��w!�z>�-��	Х�t�$�5�>ۗ���k��ʹ&E��>��0���ŕ&?"+�Kw�Z aC"=��x��%��'��R�$��g_R�>Wz�_�5�k[?���&��9�������:���5w���eD�,�Ѵ ���M�&W��O���ҁ�R�w{x��n��>�����EA������q�Clz�ޯ"�3����~س�1�߮B�FS��ŋY�m,~,��V?���Q�&ז=cnCX��PvM?1��G�S,-ޅ?�):��O��eu��嘉�f\/D�}-��=Ǩ)?���h$:�k`��N�0B��I�w
�		�q��0G��Ҕ*X4$��$�yN��c&�Ƣs�٩ދ��{>g�v计hFW���*Kw�X�$�&5h ��D/���&�@���1�o���ֶ�}�B���@~��3��	�Ņu�F�I�>�i�X��@���ܸ�֒i�#��(��p��Zy���q��k�V>����p���~�����=sK_߯~��68d;[�k���V[c�%�E�S붍��gv�`�f/���Y������n�/����.�N��L<�s0P)��)�!Ɣ]8��$�B��8ۺ�-�g�3=\AH���Б�ǈ-96�}d�����QH�K���1�P:m&�D�:Q��Q�(Ft6
�{�SG,RK�.��p�$�5Ŝ	���	1;���H0dP����憦3��S�3�������f �B��)dԉl5� &)*�x0Ҏ���*����{s�s��#��&��CXS��3wx����^�K���k���>8�#�j��F��ѩ�]�(��^�3���&�?�C�}��;��Py��*2��8PL-7����@��GПR���i����9����\���lC.��sZ��)ꉫ�������!�5�;"�xmȩ�38�ۿ������ g��e6����'SS��\���U���s�\\3�4/��3��+���5׉���H�����\^�x�����}����J��I����UY��@��N>=$���솋b`�@��.��>��z]0��%��VֽQ�8�����tqom�j �e"7�C��2�L��7���"�	3��VJH��t2d9v
��T�r��t��Ҏ<��99:��~�/D�!+��'��펧7NZ $pDg����֧���&-8��YS?q�z��m���Z/�4�7���ѵ޼s�?:��@��u��7#[�����1`aZ�xW�)_y�i-mHs�i�d9Z��pTÂܢ�nl��x�D�b��70ɐ�,(DP�I�iwJ�M��h� e����b�_�w���,/ɮ&˛�벬�������m�~1^��J��h�*A4��b��ô�W�HidF	! bcf>��Cdc|D��4�a�f}c��Pk���F����F*��ԣfqEt�ŀ�Ih�jU���6λ�L���2Jj��$��x�<6
xc��D�����k�����҂���JX�߿�+���w6���ԐgͶPa�C�v͚��z�rg�z�+�ʷ�~� ���������A���?����4u�5������}-ħ���/e�fJ����>���C]4�h�L�	��"D)5�P��Z������������'y��9��Z�Ӣ��Ik�ר�@1��4MZVVx�p�?y���<����w*�z!oOϜ�e�Ȝ�R�J6Xl{(��B�!9W��孻ǜ��}�����@Ґ9��Ԛf��t�#Z�w��mSR��� aZF.6�Zx�h��耢�^NM��'���C�����|���[�fCցsb��bpL�J{��i�z������8W�ޢ�ǣD�~�e��h<�؉��5�0:�H�]ڐ3���i��3h�7����5��^_H���ڀ[���b�����Ԩ��	��2+��n�u�����j5%��.��K���PDj`f`njh8����{>��l�˸ak�� 1E#|�؅�}-�(���-K����bf
P� z�+��h:���G�Ov����k�����C�
�'�g>@	�����xg\�vn3"�sAը�|:H�{! �Mj47P�"w�%�!}�憁C ��#ۃ|_�����~G��9gn��	��%�,2���?#Z�2���0؝9x'������&q�y&��|p.9�gK��A�j�n�z�/6�vH��y�8�0�������m��01���d����b�BY�T����p=�Xz9�2���v���貿*���4�&����5j�_A%��	V����WJ���	Ip�:1!��T��NJ簶��bCc�/��,fG\ʤ�(�G`,+����=��Q$B�F�$����V�Z����)���\���[�Ӣ��L��چ����rvy�}׊6@_�|�O�&�==+��w�w����\���U�O���#W�e��=Y���� ���-a�1�� ,}̊�kQx�T�E-~0��Oi�� �7v4(8�F��x��������D+˚�q��R_��zM�>|���D�g��OԤ��)Z�76֘���ڦ��5����v66uq.3�6,��.gd��L����t���A�ι>ϥ&�H^�˫��g��O?���Mp`�k�s�7�b�Pq�|C��׃�e�n�����!id�U�V�R��c#Ǒ�z�}Ac�<e������pp�z�6�i�"x��6����ǂ�~O�ecu��P�@���ں�1�9CX�˂� L�8��ĵa2����jD�+o���,(;dC�Æ�5���'9��.�4s!��2x1�7�f a'j�Fq=�ŀ��F׍���k��B�c�}��v{��l�}�-~T�3=}��vl��X�yu(�?=���S�)�Zԓ��|��^,9��	�����-`��D��Z�H����yL쟞��G�ӕ���H0D��i��G�hS��P	p�w$J@ɇ�Lf��C�(F�!��?(TY�M�ד|�D�4���U&���M8��ڶ8o�pķb��D���4$Ғlb?�#w��C��Hǐ���p%�9p�=��?��	gp�0]�5�k]��d �o��Qa	��..�[��b^���r��WP���J\+`�X���Gd� ����ә)��o/1q��FSf/�񁃞.�\�y���+�Э�/���jθ�1el(lP]���ed�	M4��]�hz�I[l�(�)XJ��jo߼���a�-M����g�C=��,�#��ߗC�?J�ݽ˛^�xJ�+��'/O����dm���9��](��2�dp����ե4��v����vb�f%�q�'���	��(D�w?l`���[��!.Z������.��x��xPL��1$랸7�`��GN!�S��45n��u� !���Z)�����'�o��tz${o�\��F������Y�Y�SyH̠��J/Z����!`l41(0	ד�C��Qa1�7�����*+}�I�P�h;��L��������
~�����i3��>p_�d�rԅ�7��m�l�K����Ut���,�l�k	(�j[����;�X�pӵ=�L��v�LYm�*J����3b�!gOb����������
�'�|$�Ԍ�"3b\\��H�g¯�%��r6�T��Yl�� �Ƀ;;��Oe|}&o�^��ה���`��nʽ�_})��[rxx(_���J��(Qf����iGN��d����v@}�}�n�z��~_#��RW�?�+[��/k�4���tj�=�Y��ܟ�6���DIcR �k4�2A[{���|��:.(�n4*���$�X��S\��E��r�j��f�3����d>2=v"q��<J��*���ɯ���_��(+�l,P�=�!#�jFlGc��g�_��m�l�j��4n�)7���c�ݧ����\{${pP����|񛿕�ڦ�-M�f�6(�p ��=p�� L=�+C��;�ơm����}D�����򒴆�)3w;qWк"��(�Fϒ�:$�#����S�FH@[�.�*�����>��Dҵ��H�ݔ�5��@���"A��1���@Z���IYE�	�%�Y�I�䖆3�{@�۽.��u �7� r��@N�/I�`�r�Q�	C���1�-�ؓj0��.R��kPnղ���"����ɪ�c�X����Ҡ�	k�D,��2����������2w�m$/�^Ù_N����:ϸ�8��sT����P��&���Z�Ӆ�l�1y�F;���(|��DOp��@��J��O�^Sm)$\#�G��?H�Ӡ���ŜC�;[�,0̺��Q]���=988"��hT9�%4\��:���q���?b�+i��&�{觟~��o� �W@E�f3��D�Si�!Vy�n�	�-�wA����:��������hN�����L�`�ݒ��QM�c����)�ɊՄ��T$���4�J������јн�Dn(�*��rP��[YiFם��ڀ$��kp�t��ĕx3$a��v��(� ���ĭ6[�((��a�oj$D79�V�!�k��uE��˲N���s@u�8�m�%���{�{��,~11���k$*>�W�7ϡ� ~ݠ���3��8��ޖ����AV��(;�p������A~�&ڦ�nT��11(|� �9�ńT�-�6��"B
1�kM�Hu֟FP`F�����?���jV l�zD��0���Q���o��q��+(���"�t������(�#����8���Rd�´�r�78�c����&���ʧ��tp%Ǐ��۽ךȿ%(��{H��ܡ;�X oZN	x��33��)�����82�+e��b~�Nє�M��T� =5I�Hl삱;��e�yG��̓���6r�1g��u.BO��ٝ:�%y"N"�Al��F��C�zovZ4�B��t��n�`A��5��'��������Z`5C��1ٚA�q#^ ^*@�צy��?O�E����คs�nKt�U����{DFS4:����{w���d<����6�#R��ڶ�������� �����"ח���k��@�Au͡��Н���NIɵ�m���Z�Eh��h��i��=��rch�U�9 �{�4$�lřR��-7/�x^�,	��8��z>��L��%�3w���'-�������/<�^31���cM��ک|�寴r�%����r�EtN�ZXloonP��$,�!�w���5��\w:��F0�L�f[f֤�W�s0-9ћ���]�}�+y���z������C��<$ˬ0#���T���hR�7x��/9 �ɗf�;��B��Er�xp.�r���X�l�߆�|뗦At��iax��0ȩ�=Y"��զ�M�6n�4�"��ꚃY8(O�O�����6`?�%M��[�s�^O���O[t�āen�)" ð,d=IgҤ���\������r�p�Pa��_5�����KB9M�r"�j����Հ�w�Q�Rޫd�&��SIkr�_3jѤ�
D�Ee2�v�W�A���m�#���ū�j�����_����_L���K՜1������H�Ձ�"F������0{�{{��l��ڌm�	?��LE��N{���8�˳�&N���������<�V�ٹ�!�HL]}�Fb�%���^{p>��n�2Od��cюv埾�Ff�&ƽ%�)��6�i���'��bߡUk�ƹ,}�8���)��GQ'7���T���z�>mY��G����j����{y��eT%*u����0�Wf^4��GB�@�L6"^�	��Ӱ�H�_���m��ꂐ@�Ƭ�?�<e�V/�PĊwۊ�z���iz�Am���Da�Y�=��|\wO�����/�ZB ͋P�K)*��(1�P�T�ޟ�Qr|4=���ؽ���?�0�K���2�[\��3�?��b�7�(�g_�~%�^��%���u�k ��| �<81��|ܐ�@����K��A@�AM���o֥���@{�!ႊ�Hvi��d�0���I<��$Jv�,�B܍=R:�ٿ�~��˺�Q5���-���n#���!&M��a����R�\q�E�~��'��|4�)Χb���]�^{�P��ccmS�[��ٳ�h"�a�������C�\�EN����Q���T�qZ��]��e\W�aܧ���]-���n�D�1)�=�1`a:������ �R�#�� "HN{'�D;J�m�o7���>M0���Je���8�8o�6<@r s(S:ʼK���>u� ��T]]��6���Xka�`��P���NR��[���Y<Ln��/��X�y�z%�:x�`�+��lş�e
�����_7�my��'�E��w_�Q�Wgz�:2�����\�S	��>��{���)=���~��ǲ�g1d��kZȯiQ���K��)���˲���B�+�����6�J�#=�@�½����`�a�ja�^��5�{�,��X����-.(Z��Ol�(���y��5Jnb@�$�,���ݰ���&+�k����K;����>��w�ˏϿ���=����]��i�����g������D.�Sɠxp=��6G��dx=��g�r>˛�M�JN�n���Ǐ5��R�7�d
i5 �l��0n�S�)e��ASY� �o�p]s�P��ȝ�	���L�5BT�Q��*�����縮�aA��/+���a\51 ���6�c��O��F�AP�{�3���q�:m������HJz�bX�+~oc}U�߹+�n��̯��~��[����տ�ۿ����)Ϧ�]p9���8��-��;D3�CEA�y���]m��u�H�\�8�sl@�=��$��k<X<u�w��]S=�ĵ;�a�s]��"Pi�I *s�
e �����H>�z=��72]���V�;"�i)N_����h+��3Y]�k2ܔW�^�A��6�p�)���]qn9D+4����;��_ʛ7o���qy5d���u��qYR�;��ɲ��t�Nb�^mk��3�g�l�=C{W��+Z�]M�{��.[lW���i�e8+)��Z�I~𮁀bh0
]��v�]�w�kr�3��?c��x�~�B�#&�ej4� �5c'��L.�84AV���!�<ȋ�mtP-8���b m�~C^����*���qe�p���8���3�i2@��ș^u"@���u��@kG�3	��AbϮ��%���-n��D�vZ�T6�\�ˆ`� EN�e�lD-�_S������#�G�k}l�@�g���mI��X4�E%�i.̦�n��&��w��e1��DT���[G��߹��\�	;}=����\N�pp���R6�6��g5e1�X�DE2���ä��Sv�WQ���թ;^Ĵ�~#C|��ǆ��SC�Wܐ�$ʒ��B�H��}s�����N8lx������)D�3�*� �T�.�O��:�Ëk�������1���� ��Q��-��B����>y&��;���GL�������0�ʬ�º�9�� �לf̡���k�,L��	Hy.�XZ���A8�S&n�f R��y��qf��0����b�rH�1��do��_�$�p��X�ѳ�����jO�}�y�i���� J*#����t�����A�^�T��2)Ӡ������W����Z#�ӷ���Ӫx���4sgB-�Z��(�L���V��l+�:�E6���KD���8���|�ŗ�x�p}���Wr�9`��o��	�1��3}?z^-�oA'R�Lz�r��@��������b��ڡ��E��������D�O�=�l�����6c�3*�e�M]��%���(��e���3�z�hY�oj�W����8���:[u�`��b�N4-C+��.u�ܾ(6-�t�u��_Ot#����/d���)���_���	��㳁\i��N��-�D_�X/�S��A5�	 l,�n�=�$�t4q�����sW?<қ�I��,�#a���hx{Ih7��T��}��s�^>���C/��KC�㱛	Ka�Di�������+P3����D=^(�-r3�
�e�U�� ����tK����tP��Q�ٮ6%mgt�.�����w&#�1���=���ʿ��j�����_~|�B��xq�T��p5�����n���c�U�T��8���0�E�1˪�)�хX�u@���`$xx��&^�������kgӑ����i��<Xj�e�Ŧ����Qy����뱘��4�����I�2�0�
	+ׁ@=h֊ݧ3=̰z���{K����Ho�{φvVV��{}9֟ˊ��������L��~�������}��i&��|d���8%u�7��dM���Ӯ\���F_�z�0m�⥫I8`��,�5��Zmw�dmcCή�Fe]��e��}yyp"�Z��O�:�A~����0�"8@�N޹���{��4�Go2�B�a�9�X43��ĩ��ƅ6��n1'�D��e���v��4��t��\1;{�M���[Y=����qQ &yj�&�	�������	J9%�<L�(��0�p�8��C��uq(��fZl�����Y��2)��1�y��9C�ScH�'3]����i�7@w�M�R���>�D�-���0�뗹�^W[ 8�P�	����5X���+��\� !����?��C2s���-�@��Q�e\�Ѹ��)��pGb$0��J��f�I1v�(@���QZl�}Ё�a�P'FN�*u  fu�]:��O쥖�FN�p�vX\L�o�%�n��-ỷ�r�`o��� ��JH�"Ь@����^��&>��벱������Jx���Ͳ�Dz!d�ل�����l�%}��RO�>zbF����C
 d���<��޾=0
�&�i�e��}p:hg��hҝ���$���ǸDڙܚ�r�j���m�y}-#��^�Q���d��Aj����<z�Hv�7e}����$��ɱ�+x��;w����)M�ٽ��l/Q�gB�g��g�Ba��e�x,�r��VҦ�h]�f�y�^�Nw,|.�iG�X8�a�8�4#DN8���;�VDFVF��Q�k9 ZQM���NS�=�K�WxF`�(�����}�LV���ΓG��� i��6hzP��=wqx$�tM4�k����d}L��+[w��osP�Nt�3nuu�Ժ��M�U�2�Ҝ�@#Ѡpn5l�K\n�0e0_
���$%�m�(֊�ivk�_��=XI7R�����T�w��F�˼F���ɍ/�����,��XT�fвE�LIC � It#�9�I��ր����&���A<�H������
�D�Mlt_bPí�O�\�ۿpb�e�y���.xqґ��[�n��+����w:B�rEe�ȕ/*�w�8���_5��� �HI�.��^�Q��y+p�j%�?�ZN1�?�ÎuY���s?|��Akx4��p�Oq�؆�sw�M`�<`k��> �f�4�Wn�a�0��lb�1���4o#Ut>`v �O\�aDS��pX�VP��Pn+6=jRL@����bZZ�S�
�KI��Qp�[��$�ز������{Ĵc�����5y I��&�#�u~��Z}��	����e9}A�38��~�1'�//O�Z���F#k-&E��ȃ?���F]�pl;��N�Wr������{��o��J�1ђ�t�H�-w%�3f�x&'z���0q�ӏ��q�
��{��>dO�6kptQpB%���o�aK�J<�,�qZs�Y҃�L��@qx���G����J����Z�o�e}���n�H����3��UF�r|~%�篩uwV"���Ǐ˗�[I��^��#��)r��lY���FI���*����V	�'0�p��~�M�P�b���@��H�=�D��S>(��?�%���/錈N;��,h/e!����*��!c������5�|�P�f��D�۪v�"���!K��D63�:�Pd)̤�t5*�Q���l��{91��]8iVv���!��H@���#&��.���c�3h�H8Ȉ�j����y�7<�L�Z����s�aiӳ���uU���ɻQ��ّ�Kp����YEk�d=�2v�l�:�L�*"���OK"䈑Pp�/5	T�j`�J����Hc0�B�
�܎i��P h"��dU�����'�M0D�5�ȱӮ"�ꫵZS�z�=��w����~,���&�@�1,��	v��`ǯ����v!����)��	#�6�Q��٨1��SV��6~��_�9XR��⹇����E�Ğ�O�:<m�f��}���7���)�e�� �cd�8�$��%����2���v�����3���`|��y�j=�6�P����/ ���;����j,;Q��uk<^YY������\>���-v������(ƥ��rtzI�+N=�P�ٽ��A����]t]��8��~q���;��m�s�=[�z��R��#(#��Q�ZO�n�P���]�߮Wθd3!k,)=	P���F�%i�p5:��j���e�뛾���6���YG�����DJ-�� ��l���J�ﵮ��%���#h�0y��ٖ��E#4��Z�w�H��k��x �g1�ґ��X��Ynt,�<�="5PLM��d�n�>����;��i�����~R�m��g�<Kܓ��:PZ*s��/�����vFh��@�v�7��f�`\9�琏~���M��ib�n�v���sE6��������C���mX�c�
��-�WSG�;T�X���佭��R�/m���t�j��f��EF����?Z�LB��C��� T���+r��k�Z@Y4o(���T7ʌn�%�gp0�F̸%p�����T��L!LI��!����6�x�e�.ZV�ǃrᨮ�>�b?K�����-Q=�����61�F";tC�ׁ4	oY"���?\c�mC��C���gB�	]��L
-�^��Mw�&�@ۋ0��s�4���e��W�ns�]�5�P�)Z脆��F������f{����5!Aҍ�3-�����Xנ�և_n7i��I��"o/����f|��. d�gϴ8ɷϿ1����ăd{�/s�A�e������4��9O^��Rg��0�7�{�<�����_�l<d<������p�ZAA�P������'��7�������!vpv���#ٸs_�v�8�Zz��҂:�-B��d0��B��;Z�l�I�������CFn�i,�NT�����������j燽��ŀX�!���[�.�稢�z�S�˶�zFI0��EH���0�Tt�P��G�F�e���8�G��u@�(QS��T��^キ�g%�f5�Կ2F�	����-�����L��;
��9�XG|�X�AMj����;h�H��_Z���,A:���[@;��*��y�<M��N�)e��358�Q��m3��ƚBh����'b��SX�J֋���eQ���� �w��I[D�3�HD~��-���L<�X�"a�yĠ�ٔ������jEeC�M�O�a���e��}����>����j�^{y� �5�}�,t�y���
>���	H��$�XX���DTu��%55̾Z<�1cv�4z%8��܆��(t@���&�`]T�|"��� �e^�"6Z�� �I3i��A��ɔ]O8���)}����T��N5�mt�AE�ꣳsy�w�_/���a:���6
4�Hq����cB,������� ��(�&x�C�]�~�
�b�P�"' h�b	�E�{�9~��s>��o�w<C�w��@ri^����1�6� �rp�G��� D�s��0-;�܊\l��6��h\���}���s��ٿD*_�J������A";I~&s��,t���7����%�Sl݉� *g%�w��t؋r$�i�#�}5Ҹ6/X4"�j.m���`ǥM7�T��G�|
~%�2ԗ�K<w[ݎ1 ��u]�T;�L3�Kf���}�v�w&�����F�%a��B�C�L�V�SQ����x\<�p�b�U�6�5��g����sGFp���I6�|J�y��g��i����/��-r�nF�����d4�+賴�MՐ��m�xe�����Wz�&l�a�);*�>m5�S"P6�0X���4SJ�Hޱ��2���M}Zo�TY�]�����~���E���8�&�5�yi�i�Ϛr��,AN2Ӗ�X^�����E���r
T�N%�#�M'1)����b��Q���Cc����W�Q!@� 'H`��Tx�<Z0�I=���bᇤ������M��qC�,yK9��dG ��p9��*�r4��Y��/H�+��҇��V����|���������w�,nJk����x��`qeV�0����e��Aype۔)�C�㏟Ise$����Ŭ���]�3щ���s�/��u���d}sCNt�{�	��2A��%����ך�!�#��\1@r���C�O5ٿ�����յ���&�nK�>y$˽�.���_���ZO����L^�=$�� �~0qO�*��4	0R�"h')��G3rEiÕl�a����$��q�fK�p�}Ɓ��S޾7�I�o��ͨ��bP܁:�?-�
BQ_�ϗ�������yl��9�e�[$�L�%iޖ��Μ2d�AQ�Y�ϥᒾ8Pq�a䲢���{�z�6eC��д�-�� tY�ӂ/�[�%�W��L��;2�ʜi��y��<�w��`�ݍ@�AB�5Z�(l�x�B�9��.	�Q5Ȇ�A���^�#Α�@f���J�9��@��0��/>��NH/�C��E�(1$�a�R�9#�Ž��Jo.�ur%ޡ̲����w��,��YY"����׆���̦=��^��jL�>f��x���m�(tؐ�q0��{��.�'��Q���������~%�|�q9Z�������V��N�A�q��.��b�&n1���I0�	E@���N�hij"��%��rn�	�Q�<�f�D4CB��1����&ฎ��f�7b�<�[j��,�
K�..e��+]�{�¤� �a�$C�ܡH˅�j�?A��5\P��;]X
�z-T ��jK��|Y�(�pb�)���q�?S��
A'(����3�y ��3��?`�ƞ�9O ������7�!r50 �غxl{��4��j<����-�2�Y�HF�+"��eZ8�v��/o��1c.A�iFW�I�����*õ)%����P,h�{�Ü��Ԙv��!��~��&�	.��x4�\�p	]������G���%-]8'���x���$(���* �<��� -\���<�x��|�\�~�p�J.R	�H%1�^~�Y4�,���(#�'a��۠S
e��TRƣ)��b"SK(\�-0r
���&DMo�тTPh������NC�0�^nƊ�E��&��{O?��@�	�H�Ƶ��@82����*�����YѬ��+�!*&&�5�J�pa�\��[f�\�%K
YL+���������!U��R�&�J���qGV��&���'$h8�S6��#�(�M�p�f���H~p��9�h���H��"$�'�m9i��W�1����H_ɶ/���`5�{\���	p��q	�<���d�����
M~ �߿|#ӓs&qA>+��ϣ�)�"���|FXl�hS��:���Ж b6W\�-��5�Їk���C�C��	�SJΫdS��J��5�C3�9�--/��sB�k�� �u�*eu���Ͻ��)O?z(�K=N�C-h<?������_'�g�P+�dQ�˖�����l���m��V�
pܣ�Τ�s�E�~����vK��2D�����P6�q����������h$�����P�&��UZq�C��:.bC�c�	T`H8�m���[?Z�f�е��W[�/��QH�G��x��u�a�� ��ݻ�_?0Cq�ϒ��g�{h�D�#H���ktm�9L�b���}������O���|+�3K��p\Z�b����9���/��<��;[k��tI�&���V�o~�k�����t��P��"T�P���q(�:�W���7�~+����<Ľ�� @��<(U� 7����*�� Wڭ.]G	]o�-����j�&��nIoe�?{y=�ze,r�U8<s����w�#��!���\8{�7���w/�p�T����+��̿������\YY��r�A�sFsB�w@� ~���0Wb��
˅�����{� �a���ZEy�j�w#7]�Y���
�>����g��r��H��:����`@��$gꅗ@�e��{"��`B�U�?��皀���EE��`i�nl�9B�yxb�s�#���5& �p<��G�n1{�1)9bg�"	N!�Oq]�Q�9҆3!��j:Rb���u]��R)&2�o~�:��iʛ6ȝO�pp�9�w�p=Aa�yHjЙ\�5�gc���d{k��*8�ΰPG�O9������nP&1��)�ʔ�&s��k)�o̳�K2�j�V�oǮG��KKE	O�6��  ;�n��D�A��G�3&��S<w*���1���L���� �&z6��0�j�R�#}M�W���� ]E6��`4�:W��Q)-/�l&C�:6V4D>,� �w��?�E�(\�Q�w�`�9�Ɗl~R���<.���7(�f�ju����_ڢ���F�4���N�E[\�L�/ Ŝ�P�Z�(8H7�����1�C 0=��<i7�����Z�-D�/l@�D��o,ŜR㊷��]�-k#!�����-~THG ��I���7+�g���5�<ޓA���,P���4*�5e�0�٠��	<��i��qc�y�΃�)1��8Р���~<��~6]@���F=�ZVEHTq7!��a��UvH��m�L�/w�g�3a��>9�Pc���|���%;=�ClA�N�?����7q����"z�?�b&CXm�>��h(J�:�����ށ��{�➀v԰��(yn뒽�Դ��EI8���@�i�:M��H���;I���A�$����W�^qv���T���8��l���"kfP�X�Z�bx0�Umz�V ���z�ZQL)2��F5��"
6��;�{���O�n�>Ϙ�ar��he���LC�&������W:^�͝�hM�����Uʊ�a9{��=��o�������?P�9_;�#"i6�
GI��� �@���Q�_C��~�[��Aqiʝm=Dw�49���~$���4^�$R����B��5����??��?_��ƪ���z!!��+璴�\�ʛ�?�� (����k� ��u���#�>���<��x$�|��[�A����#�&G����[�O>y���T�7��Uw@�C�i�'���#��یo𩠂��JV~Fa�u��p�Y��~�S�8x ,t}X�����9ML����N�	:���/��ٸ��Զ�i��ZR"S.!q�h������u&�NW���I�,�.��v��ҕǌ+k�;3�Z�XZdI��E���n�\L�+��V�ZF�{��̠9g��?��̽����h>���Vn�����̲u�����Cj�k��m������r8�e�$���� b1���Pc�\��;H
s*D���M8�s�XH�2��^%�v��,t�KO.��݌h��8��DR��!(̣,C����L� �4����\ e����<T4����4�sxN и�>,��ݏu�b0vt})?�~��kT�Jq�Aぜ������~�P�=���U*���e��� M�s��N��$.����P��\HL��R����,�9�(�o���:O�>X��3F~��u�|%v��;3D���/d�0�T�g<�J��h��Y3yG1��,PÒx-D�k�-�6�M�)�)��X��qpܕ��3��!ܖ6�g�6�6"�4��{?,�ү~�tm�x��e
M�GEF{99<���ܿ�H6׶i-����7�8�=e�ې�����kBڪ't���]%�
	70.e��鉷7���Jl��x�C�𐛵�E�1��P�R,��<�z�X!��~��Uxʂb�M����<�q8u� h��D��cij��nĺ)&r��J�b")��u3p��M-8=��)0\*��&�H|����Xz]�h;��ʠ!m�s���\[��e�h�"j�R&6� ��q�����-�z���t\m2����*PO�?|*�P&��5I���p��By~�FHB+�ۑ���U�1�n>nb�lI\��u
�t�fWN��姗o���m�o�,�4<�Eԗ�}ys|)É#,�ЂðM��Z�Jd�кK41Ga}qv�븶��@nH�A凯�L�����t@4�)p��{�lH��n��׾����$}������jU���WV��\�;�>�E�S��.Z��O�������i��Rz�������܃��X_��S���+ѱ�{T% э��Z9��+��[?j	ϭ�o��ґMf$�ep���C*m�=�=ph��b'�������!cR�6>�k�����k9J}�÷{�������c��߁�hf�?�P��ۤ��󛿑���_�������;}=SCa�\����{���?���yHy!(w��Sy���S�����O�r"��hv@����X��
$�6vvx��9 ���С�9�C1h{��%��.�,��EH�;��^���QTTB�:��u7�v�gI|YS,%� ��z�Ox��1���__�8�u�ک��۲�1��D+�BP����Fd(@AE,h�[/tZ-v�MX���%��Y��o<%-Պ;�Jx�Я��I�P�euR�}^��N΍$r``j�TnEF}&���af�e���Q�ae��i3F��h�H:Sd�����By��#x��S��WS�E�h�Q�7~(�u{s(�u��q�po<!��c���6=�0��v�|~�5�Y�����,���?�:�Y�@±8���ӧ�>�L�|���Ѓ^�>�w����fS�\[r�U���NUx~���o4�^�|c��}:Θc�t-��Y��7������yȹ.PN:Kk�b�`�-�N*Nˤ���	�x6��7���]��Y�J��p�9s��������&c��^f/�<aD���b :�� #�鹋%�o� }���5���_�F'6D��3tf{�`T��I���;��9&;ג('�6�KH��\+=^���ce��&�E5�p?�Ñ�$MV ��2�@y�r(�˫��b��4�� ��=��è��5
�� �GHB��X�7y�!���������gC���YV��X�6]��	�m��s\1n��=��q-�z��~��Q,��n�8�wͤ�Z�H�/�C��J��a;)Ƀ/X���o�y�@i�'�!�L*:P��|]^��`�n���W��]G� �I4�<=�sA7�����Y1.�S��X�I��ǫЁ��tN�E�n��B��|
3�28O����>ܦǔA�/~�D�N�?���Cel�C�&�U)��T�5Y��"��*� 2xS&۸N���ĸ���k�?���Il(4�S
hL�A�\X&Y�u�P�����IE��Å�����l��.O9����2�x���5Δ�PT:��̮\^���TOp�lnoʧ�!w�7�����fb��q��E"���sK����f��:�4�C��.wߣ湯[��@I^��+���G�O�������I}-����iA��j�O��ڎrw7V�ʊ$<_���%9>ؗ��@��c��ڪ<z�ĸ�>*�Ȝj5��i]_�ޛײ���{��TZ
�CH�y0�\����r[��n��řl�,�ϐ�E�f<��^#�.�����c
J���|q~�k`��(o������&�a�A?�?��	�6]��-	}8v;����@�����5��W�|��H�{�����q���ȋ<�:��=����搾V?[��w8��;q��m�{�;�<0�2�:��E�
�8?������+,Q�x��ܺąw���*��4R�AY(�(��u�Ȇ�S�L9�b�C�l���:�{�qQ�j#>���jfǶ�`��g�wAf������c\��9���	��/|��%�?I촃�h����B�^=_4i�н�J�'*���"4!��n�RG2Ʀ�I&f��4���BRr�����Z�?���n�X�?e���u
�{��^��d��M�6IHt�Q �|���*C��-���A���sF3���}"[���|��Ϛ��a���xG ���%/	\��>_���w#=�4G�<�3hU�Zx"/�\�J�w8�Iu����Ī�}׃!;��¨�BRs���z��<J8�)w�K޺(L%,0���������ld���! �&���9��c�L�q�)��B)�B
�ǌ$]�S�|2�\�M(��)��2X9�ʵ3�9.
5�R�.���|�\c��w���;K'�W�x4�8�O[��3����sNtcyi����u�oﶻ2���u��F�;V����*s���CF�r��-bS;�)��T&��8멙�8"���l21��]�'�
SUѥ��3oE��j#Q5�Vo$�
�6Mh��mY�Y��:.k��j�����P�����-i�y3ͤQ�m8�Wv� ����h��gЫƝUvI�p%|x���np�g��P��=��������#�ZN����&��1�D���l$�9�;��8���-]-7Tؤ�RC�Хp=m�3�TCYL�l���y�?����]�_���kX_�(L5�ڤ���=O��z��U!k��ܻے��3�ß�������F��v)9Bl���0��#�_]]�����ڐݻw���@و��h���+kr�����_���#�eN���}wsC�}�T��Wee��I]��T�G���@���7򧯾�7o��l����8�(��i(�B�O��OٶI�A�����R��`��uf�pd2{�{�c4�� �R!��ź���Ȇ����߽��_�j=�G1Dђ=���>J;���l�_�|�pWz�����\����W?˟��G����de�'���G��~šf�2�}���L�^l�m#6k�*��J�L�����s������8���{2���N=y��ܻ�͟m�J���{9��G��g�$9@�Mq�2��sJ�+sSp���(�Z� ��hcm�h2�w|&m��ņ�@����n[<@<I�j��{y�I>{k���=�}�Z���2�J�
[��u"7�)O⫄�B�E��(S9L�7�T07���K-��y�b���(j��Xߖ�;���m�1SSnc{�j��*=A�<9�=b����Ph]j%
�E��'$	�q�:n���U`�z�6��x��o��9T�B����ǹAӡ?A���%��'�T.B� @��qoa�9=N����Y�(����$�!oA`�3�ù�f�Xcq�8���yTq����&��-�rC��A8]�ғ���{�U��y]4EFo�p=�<.�B��f�:0�,���/��d�@�޿'>�u�L��Xs���E�5S'�F����%��<~��]�٥ɗ���KK����)�wFr�)�d ��:�s�r���s��]���>_Wu��p-��T�<~W�"�[�Sc������p^��k�t�$o��M���z��������i��?GùU�.D$���Zm`�|L�{�K�+�g�0�� 99�QR�oUܷ�+��[a��X��z����
�&/��m4>-��B�������Z���tV��p}�
_lڹ��O��.�\���DN����+J���X��u=x�e�����ۜ2{�DG~8�4�Ho��gp`�x�69�\�ث*>NY��f�b��(�\�L��+s��+Թp�'�����v�4	��(�b��U�1}��y$nTf��Y��ņ(F�Ҏ�����h0@�0�6����!��4��X���ν-�D{,2��N�o!�ܲ`_+�4SY��THH�R@����W�I��s}u���2�����фeww�w�@~��ɬ�|�Fp���2��m��	U/<\s��G���gz���qe"/��w�G��A��n�i��^T8�M�X�
A��'��'�Ƚ�]��\���ɩ���48.�l�4��c�駟���3���)k}�����!Y��B��wY����B?}B5���Ꚛ1�`݁���ԗ�I[�D�PG���]�Bpl�{�jv94�ׄpC��&�ZP�fH�"�e�.�4,��脯��m-Z�:]�	����Pɳ)_?�m3������
:j@��u�c\+��a����P��p�2�qT�k� �^�������0���B�w�·�"FI�y�u�\R�s�so�z}jW����=�>��C�.�����뿒e����@���?���4p�\���"����K���F��]y������#��ߓ���ٻZ h����{�i�:�.����[J�޽�C��u������஢����>�F���s��J�@��ۮ�9�[����u��ҁ� ���yx������Hwat�:�&A#v9��5d�^�+��T��螞^��T2��ez3m0��h\'��}�:H�&;��WL�1"�Um�{\�D�2������C�p��GDH/�de�ZV7w��O���H�-�u[���_!�tzy�	%f��I�e�/3�P/ģ:}	�ka�.+����e3Gc>��3bq���2$����b�Ă�Yh&g0��Hj�j� �CA��5EEYq�鉀 bf��8q�|$��+bױ��g3?cq~�4W��t8�scj��M[��7ya.�zFL���k��A��Hlf��������-/)�Ⱎ��=T	~Y���O��1�cs-�glT�g����l�{�I����ã}9>>!�{��<}�TFñ�6� ��CD�Ν�WKO��gz&=~����:)�Е���`!u��g��	;V8X�& �;����sv��K^������C��ٜ���(mn��H��+�z�}قl�܌��������M�J~�XH�+�èQ��>�Vk����W5V�r�������a���G�,�rΩ`�dISw��Mx���X7L�����I�4��H]ZWWk5�3;b��b���Ҍ��@�/�iw�3`wq�ѣ[w��"ufD��s�"�jzfA2�j�D��O�������Եh���,2Y�Rn{˘)���cMWa���5��i&��tmy��6f^|E��#��g <RYd��-���t���R�m(������d��9�ٔͷ��~,w�?��n���)ͨ�>9%'
� #�rO�E쮖F��%.Ҡ侱-v���j���K�����1Y�4��'������q<������sl���Sw����P6<(���p�G�d#�^��� %�Ϋ�Y���A0����p]�(��23��pV��z��]=����W:��ߋ�=9�ߒfb)�
�a��[� s |HA�[d���4� a� ��(�b|"��2����ԵX1$)�x�����h��}S~�񇺉�&&p�&k	8h�������g�,E��jt��<t {�$����*���P��x�k�#Q w����������IԎѱ�&�olޱw�d5)������~ڠ;`ó;�o���ܱ����yo����h��9x��z���i�����:�!Z��>�����mr�sG�Ut��3:0�8LQ����s:T�,%���A�~]�s��ّ�����O>�X��M�<CA��ϟ})�������:Cj��)W�f�t�0�~x&��O���q��d�W�O�֔���H�B�Z�F{��4�f��G�u��U��n�ˈ�+�;c�N��񯃖s�;����ە��l_4Q�r���@LpJ���D{?P?�ь�Z5�;i�p���_�X��E�k����A<�#����TM�n���|�FԧԦ��������Q1�/�0���r��M�{��:�̓q0�B68}]��ɓ'T�1�qZ�a}h����0pn޸M�����}}��-��xТ��� n��"�4�E8+��S���2��H�Zj��T�"���;������1��r��3�4�RښEq�B��Z�a�z����류����i��3�ޕ<�ƈ�
�2�8�X���8�+��Ĉl���Ҙ��s��g}����Y{:��yv�� :�� V33T�t�T�ۧ,�ЁD�q�B.��٪�Ǐ��1���b���/!�wčh�A���;-�?��<�A�CS5�GE!��O��!Wz�~�\�hh�ܲ�I��DP�|`W�+(4�=E�v��������V��*)_�{T�j�I��Ίπ�E�83ՉK��:V��C�y�w�\�/(x��]T�z�I�f��Y�MT�. �l]��v�e̲�bͫ�`1B"(�X��� \�8����B��D|g["���y����ɾ�N�'�ɱ|�����M@Pt�a��{�m!]Kg��숵8Șn�yE�d��n=�8��a�xZ35�QvJV8V���;��A3��m�<�e�j�1m���Y���tC�D�G��c�?�T����lA����(��5:�����E�6���UCV&��o��� +KU���g�V%P�bMLT</�aR]�hޕ�d���$Eĵ�A�F��3��}���n�`Ot{�Y0"���0=k2��"F"Vㅽ��w����h��J�;2_������m�����n�<}W�=<~6�KEMn>��c�ܣܪ��1Z�1%�����&�SQ�Pm�X'�1ZH78P�X�%�==�Ȋ
)Ez��:�4aP҈<ID�Ǟ.D��&�j�Ô�#l�&���̽t= ]��čL�;�J���N��6Y/�4���
��
sfI���4���f�b)s4U��t�@�ڿ5] U7�Zd�Z����������J��@��.؄�3R���}M7�J��&�=�g
�"�(��G{5:�3���,�E��DFcQ��o���ϱ]�xt��
�5��C���H�������wyJr�,�D�O:i�͢S!6G����h�$J��:e��nTP�$p���o�02����(�k�ދ�Ӧ�����{��������UF��
п��[�;�s��p�3O0эV�`�����R�X�LC;g9(�X##����3������/�Ȝ`4J����ͨ�nu�|� ���W��4�����Ky��5*�`ܼ�QC���ɿ��O��?�űq�ӡ]>d�>�5 t����?	5���@�T�O��/:��E��h����ɓ��9_��
e��,p&7������[T$.��U*�%����#�b�"��b��h�~��ɞ�n�֛��>A����{��'�0b�y�j�p�d􆃎4�U�A47Z��e�l�v��mH��O���m,��$C/� '�M[�!\Y[f��8�X�3�$ �r~~&k�̠�������Oj@	|jD8���u=
���\'!���G�
�rg�F�Lb�7�����4�[�[�7	�0�\Ճ�RVQ�~�s#�i����d��G������A"��'��}��J�lﰓ%Z�j�P��3��uh�gŋεO-�P��H%:�9���չ�"Y��q�8{�@/*�'��(9v �sR�z.�gע6�l\ا��b,�(� 2�8��q^HE���=�������3�WV�X)������K��=t�Gj_��  T4;�yQ�m4YS*/�d"�[mJI����h��9��>��F\��GՔ4�5eP���F��������L������Dvٰ؉c�)�ř0�ɞ`���� �s+���D��\���V�p���zAft0����C��ܡ	�(��g�6�����ɉ��ݷ���Kʳ"�芰�8s���K�V<LE=�̲,Uv>�1���׬V�<q4��+x�{��^6�7o3(0���P�s����7���t��i�>%���4�9�����#�O��ĳ@�E����΀��`�2���pF��X����͓�G�T�(��Y��\ca��L*Uj������z�wݫ]]�j�G1;ǳ�!Pʑi(�˫:���,,�(>��$��4+ٿ\_��O�fן�x��g�E�'���¦��K�#���ƍ飛�N�O>��5R������SP� ���p��Cq&R��H��S<��S9<:����xHД�5ĴR�b7�s-�@���B��"��1Ba��}�D�%�{^0�A7���F�U��L!��h҃�DD�N/�2�*n�ں���i�����
�@uP�j^�.�řY�i�Np���O���gr���
���y b�h�fC+�K+b�b�B�� !��/��\�`ȯ>���.x�<�
��G	Q!�V����.�IF�� $ 3w_�����ekF�hD*�1NG��Ji���GP	ڳT
��;�%���̛��u�����?��L����Q>թf�dWҝ�91b�J�e�p`@�M3�-�4��d����;���f�*� X3,&,
a�?@h��l���)���I�[Z1S#xzr��o5������X�5;7�+5�u��ᇺw�ҹ8���u���>��� v��]����������"M;
�������14���b�`��ȢZ�:4ʨ6�-�jN���ÙBJ�k������x p��m\,�&/)�̫�=�r2���I�U<�]�{�c�k�NB���"������}�gf�@�E�P�������#谏7�_׃����`�*4��3��tM��Oz;���7D�ġ�=�H�c��� ��CV��f���+�B����������E�]( 8��Ef`Q�r�Ԓ�N<%#�%G�<������Y5w��c]2]��{�Y���&dV����>/�$��� \�m��>�G�0������Ğ�g� 2���#98:dGcvЎ͉Y��l��
��ž��U;O�pNx��j�
8��Ҥ%�KAR�X˓�C�T�N��i5�o1�A����<��bm��b8!d��:3f`'�@���&�Z��;ջF�b��ϽsgB�aN�����o FҨ�Ø9�)���I��'��e�?�������9�A����8�z;;SL
�k�r�tdq3�����EǛ�j�t���5��[|���I�E���ƮD��<�	`�d�m��c��E�@,�_k�ij5"���ɀݸP�g�*�qj�l�4�<�g���"�L��pX`>�H��'��<�B�g��A&=i�tM�ώ���9:�a��S�t�Q_��BpCd`���q�.{� ��EG�6��Q�"�Lb�B����d�&2Jn��˹�[NlR���������=nDz=����:nB�c��K���7�� �'���xĬ����Ag�}�T[<��|2��e����,�}���r�����F���2���vc5��_y�$�O���/�Npe�4M�^��#�ͷ_���!ӭ7��������:��u�L���G�giy�ag��Vn߹.7��ʝ7�`/^������ӗ,v�$XRmmyÃ��U+ny� ���?wQ�"7�ȼ��� �uӞe�J=��M{�݃5����5;ѐ��Q�ȼ~��"2X�؈:�}}]+�/d�Ք��;���a���[9y} g�O�t����Cn5�ꭝR��p��NOͻ�eC3f^�$Q���a����e�_�Y,���2(��VH*��b�C|�?F�t��ب�~����h��[�v��E��
�yFA9��E�S�l��bt���)^�Q`piV\5���G]���C�R�F�ȋ�9�o��B��}��ebҖ;@p/,�˃�1��*0�X�,2T�o��ܘ��S��;��Cګ(��P�����V���[��`h����w���m���RS%�^�b������o?���/)��'B2�v�t�#Y�֔���,	d�@���[,:8��g�_�J�)���F�AۣS��0b�HWӶ�R�M}���y��#I��q�Wv'dV�M*�v��\&5�&;�݈�ÛE%��0�����<�f�����6����ͤ�����@�re���s.��ڨ�3���&�nݒý�ӿ���8Qޗ����PV�M��|�oJMS]/7Ƀ��
�W�~�&i1��e�Ea�Y\�	�%==]�pX]]����x����@r��[��x/��������g9ݣ1�_�a"Y֌��K�>��b����6��b\��E�}��g/O��^�ܸ[`����%�#)hz�.�e�<��������������änQa�B�*��cl��K�DL�2ܳ9����T�. �6i��Q[b��G&��z�%�2�|M�SZX��}�??t����3o�8���F[�]B��wr[#5�9pN���k�#X]|�m�<'��c��%PC���T�A;��=)�7�Ú��[�(/f�l7��t�����dn�A�*Z�#�[+jUƌ*{m�A3�A���*�\s�����
�}����
r�iV��d[̷�+X�]�$�@(�Yv� ���@�
(dXQ?|3�@�=�q�\��-�jZ�?�Ad� k��9ʌJJts,*�t�L},����Y8����$=	�ScdH��;��3��|�_�VA���^�L�w*E��=jF&C.g/�O�!�~�R���eai���{�;�T�nߑ���Rɬ��;.��"��.�%�v����������4��d�#�8�� ��ӱ)������+9��<>ҽ��lr]f�&�׭ s-h��x��^���M�֒B��Oz0����V,�H�f겲P;����Q��Z�ڗ�����E�)��]�AN8�PH���i0�z��Ǉ�u�+�yz�Cp{խ�\(P��n�{���r����YY��끲 �[r��J�^�.7	-�bf`��I�m<���*jH�%~M5��ɱ �Y}�*a�fZ�/ �E�H'��Mt��ա�ߵ�u�����N�/�>�S�(H��ĺ�РH73$���BF)\��љ�?�+wW�rr�+��P~��,$���jM}M���Ѱ(�Y����f�JnF� ���}� �i@cŚ(��S^b���K�� �C��x�-2�(E��x;7�P�U�D���P ���-!�Q7�02�Q盗߇�|�8'o�1�8��Y#+S��-�A�H�VO���I&WW�l&�A2��/��~/R�6� �7�m�o~��ܹw��f|�iC_�?�[��j����c��AZʦ/��ew{��:��a�ح;X_�n��O =�B���ǖN�4�~o\Pr`�qo�ʷ�[�)�G��&�N��=�"W8�����O�	e�c�.�2*�h�y0P9�"
�t�9֨�`q��6�n������������D�Y�A$I1�($���/����&���B���L���E=/^RZk��o�#�Ӡ�Tp�=��W9�%��y�,++Z�=�x�..�3u����3r��_~)_����}��W,d�nz��]c�Y�2m��D�����bS�N�&"�S�-�����)v���ϲ��@����ܳw���^��$��ו�:ܠ�����(ƋL��y�u����I�&{( <�y�#��x�7�臋������V�2.�� ��d���f�F6�md�Q�k ���H-��E����8/�brg+�� 5�ljdZj���d��jƕM�*c�Q�S�`t1w�ui%�����(�=��<+���BAe���n���� �����fшj�k��97����_Sl ��57V���-뚋�B��ž�����7���q�l4rg"����du
��gqmIVVen~�T�X��0@iCt�m]�1�"��BC� ��$�֪s:� pvj���nw�u&5#��|�濶D<�a�k�g�s�,���9���F?��+Ij=#X`�g�@m&���-O���<�V�|�h�6�jmd<T�τ�U��,^�o��{P�Q��ŕ�S_]Q1�,|v{l�NGF���-��뙰�`�w8s(���Fq�Z4���_�s���������񹮟��q��GrnF�[q�hz��l*_S�c^�hO*蝑�; ����?}t0h�z0B,�x�O�Fل�tUFg벨���Y=�t,��d��4�{2�������Lb=ף�:�}�sE������r��u��`�2�t�F���Ҍ�Q��7���R��g?��.����\t(v�P�Vo*���͢�ȫ�oY�ƽ`�|������e=pzc��`������׽|�`����ή��k
8��[�'�ϭuyu�H�$< �h�c��	A���\<(��ZT������^l���=�̪Lo�����f����u-�[������Hd�z�����S�k�n�Gx&'�o�Ƭ�a��Nvdc~F6(�~t[^�_�����5 ���Ɂ�y�\��E�Qev�c�s5C�&ߥ�Q�ۏ���܆��$�^4�r����$���&J��%t|���j�ЋFzх��}�����E��8M�v8��-ә1Ó&F7��X�3�	��ŤZ&� �&V58#?7nE�0�H����z��8o�7�~�49 ���5YZYR�<���M�?>�aX�Cd��M��
�`8F�Í� ҽ�ƯެqmL={��#�֛o��/�ҿ�CЪ�Y�'5J��[D�zݾ���%�:����R����Y����ԍ*�]+���_	Kąpx�yin{�D��:*���x����C�WbK�߼�!���&�L�N#����	�Q����O�;}��0����̓�d�
ՋȨd�ְ���l��bfKS�<[����\����vV^+��?MU��<�<+�k�7��O�u!Dj����K(���=���/^����2'͆ePB�$:����
�ť����T�i��nfE�ԩã}~����^��4�-����ܽs��H���}fk��lB\dGqH㽪�~!��/�����YV��e\2�"9��RJ�x�%[��ru+�3&�3v�XR��yq��L�
��r�F�(�S^I���\��#�;�����"���/�cĺ/�����͆}��;��Qh`�̧���D�22,�(���� ��'���\�#�<�}�Y����������ݕO>�����/>��	=+�m���';[����Gr��V�����|���I�0=z���y��|���� �8#�R��.+7e6�bg�a'd��޻'�nݐ���E�umn��߽�uks��i�7�l�^"j
zɎ����1�y4?�� {Z޹A�U �3��g���N��O��p\Oy]��Qj��暑������;�&�;������j��}��ר?�q{.;�[rt� f��:,�F&V Cr�5SamIʵ�]�Ɇ=:E�l��
�_���8��1Ll?����I���h���j~���Q˧�I������޽7cm��T�'����c��I*�ȼ��;v~>/�΅\[��q�X2=�"��9V�x��-VPݗz��Α�ˁ�h��k�ƴ���9G��)h�]��vJ�|\�O:'(н�F<�Vb�����\S�P_t�'�zE���`��rb�j� �eK����:���B;>�eҬ��գ��v�i��û!��G�=�0�%aeѥ֨��*@nR� �#��|d�fl<�S���	D�`��s.o���0�f(��u�)8$�
���G���ģ|��籑ѐ* �JCh� ��Ŗ��R��fgQ�	#��Z6�V]u.ԋ�8�����!���D��(������r�b��\�J2�F�7'�L�H{W�B�����m,��L]f��:	���=U�5�Z�!��x�~��<��A9���\ܬE��{��sV:��̳���$��
Cy�L�B�O�p �	��6�A�ir��O���{�K#6=[<�1�?�%Md^tu(g������+�4`n�B!�f�����7���kv�[��X]�X�� ��"!�t�w�ؙ�T*H�^�h���ꂵ  ��IDAT����,����b��s5�����M��:~�!U�׃��˗t\�Ƙ=~�X_Z�;�����z�p�/:~.�� �w�ݔ�wn3:M�*9���9�*~ eDl�0 �§@A��Gt�������55~F���}v�!S3�|.��fp�~�f�������g3�y����55��끺�@��$�6�i���?���@�쒤���s{LZT{H�J� @�z1M$߅Ws?䓈{�;.�'Q*�k,���b}O�@R8��˘���
� R#�-K32`X��N����=y�@��E���enqEnݾ�(�����)P��Cz�o��9�k�o�����`A[��d�y���.(׬U�H@A3>`dJ�Αi�0�"���ߗ��u���ؙ0����K{�64��#\���ԣ�iV4�1Ŏ�v��2�8J���Ц�M�n�Ԕ"sR��f�.�0������X�͉!.	mń���k��e�C�>�p�U�N9c�GA�#d"�#�v��S,�l��c:�	�T\/yC���N,"���U�U.�/Ғ��O��ݶ���/���x�̗�7�;6�2֏�{Ľ�����/�+H��n���e���q�6<~�A��ڡ��1�f}�r�PZ�A��������{�7�(f��(4<��=�^U�[X�_��r��=�mw/d�����AJ=�T%�6�����c � 4�����*#C a���9�w���X_Q@��㾖P^[_�׵������	_93��yXw����=��޻��|M��i�G��� =soJY�9�uf�)!c�&��YE<�d��HB.����Qa���O��%k�\ l�Z�j�p_$ERQ$�4#:PtH�<<?��=k.ؾ���Y���=�0�T�#���@�Q$�#*d9 ���)
��o�3P
_C/v���C��q<T�^��h��4\�.��cf$��#���r��(o)��Qۋ��z�n�WP�1/�Ⱥ߶�u}��(�����O��M�u=�٦	P���!�JE���ʷ�>���C��](��Bn\[��/�̭j�&�g��D����I ��
�#4��@�]4V58�aJ��j�>���}����
6�!�����%��7׬%0�jaVOp ��Y ���@D��6&x�Q��BJ-F
�����@Ɉ��8296O�b>p��Ɓu(�`H�$���F�q�9dZp��i�^�H.��r��G�,�Ωz�:h�3S��E��4+2s폻��*x���{��Z� �`��H�gZ�toK�κx��v
!+�B�x¹�'���`���A���\�$3��W^n�߫���d�B�:�����}��huH ��(�.�� �S�8�&-,�ɭ 6t��{��J�T�m��L\��Z��8��gT[S�ڌ{�t�*��;����ڿ��a����c��_��T�t�%�u�ԹO���Q��������F�Y�e=t��C� ��O��ЄlH�MF��z��_��-,Q?� (DiBgXD�s��6uݍ�����.�9�F�<��Rj5b]F���}~�>�����<��Y�����(�3��%-����?���>5�B���9�A��������2|�E�I��لG�3��^RF.�/���#p�Y^�y��};=��@�$(Z?y�I=�wD���3Mc�����T1"Z��X��|#����9�V�-4��qSNԡ�?8�;w��ǟ������D=�����W�H*��f�\T�lnm�x<��e��Q�n,�x`P"�k�
_�\w�G�8��� *"�d x � NA���j�(,��{��.����y����d�5�sI��e�R����I^������'�b�N���{���Q���'?����%�^��`����E6�X�U`˩!c�;qGQ�$�`<jGE�������1��&E�7�l��:��s:���p����xO/���[O��^��6$����s��t���{�5�_L)g7�)���+t�f�6��aN�d��;�(��	�E�c#�ܽ�y�曯����o؇�(Uք�+�qm]nݼ!M]ǻ;���w?0�
<��Cj����--ʊ�驖���+9�ݕ���uϾ��CY]]�=ݷ����<�!�2���	�26���VJ��6{��/����}u�/�?d��:����Y4\S������X[�<�������A�fHeW�i�1!���U��'US��s��{qa�R�oR+�żo�E;(��-�5)�'5V?�`o����
������#s�paT��g��IU�>D�����X�� ��}�;5��P,��m���:cU����>�}}Cn\_%}��9Vg�P�O!ݫ�\��A��D��#�7��-��/dU0& ���׹����=�#6J���d�s���lWw�Bi�NO��^�yp�:��T�Xz�?�>?	�+�<W+��V�%N5k��c#�fq���w�s����9Ƚ#�����Qc+��Ы������Kf���ơ]�E\ǔ꺬YpR���CԠHY�m��`2)8t��;��&�o�2H���{BI2+Xaw9P�5Ɣ��M����V���:�j �T}HxB�dV��jrzv&��n�}e�^o�:b����וׯ_��k�� �<�C$r�S���$w71��S��4{[�I����}���{T;��'�H���ms�4�؀a����Y���+ȝOZ����]Q�+��@���`���Ź�"��\P�J�!��<�)�H��)��?����+���*S���č��0�~�H��E�S�j%Pq�4�N6��89���U��MU��0?Ϩ+d���?���G:=ͩ�J`�G�@�
����#O��JV�eY�fm}E^l�~j-�V���?��ꚬ����(�C��i3� G�Ͽ�^�u놼��#F����M677�f�s�2V����H����1���jfvQ��#̠�<��[f�H4?�lA�_\�G~"�Sz������c���3~8�AG!���}���g4���qB��c�܋��.�ג��V�0�a?� ��gDX�w�����-�g�.e*����H��U/��������鹼z�-��z�$��׵y|&��O�,���o���gm������B>����n4��8�Ͼ�L�w7�����Q㏈����<}��I�����+�	��`��b�]7?�C�l]Zy�	�?�2x��Q�yZ��յu�]�V��j
2HN긂��u	���,CjT��^1�u��d��[j�c���7#ږ<7��;s��g�hsP�	�=um�I?B���t��g�Y�z�����|��F.���(p���#�3�{��/H	��Io���@�����D��Bmu/>�.�f�C�pX�p�e��(���2��e�4+�Х8���"����n��EDE y߳Ȝ��BU�ԍY�(�5~@ ��]���)6 "�B�.P� nPS��S<垕�Ԧ�E1?h5��O?���ͧ,R����������y@c�Zm��'� n\�`�{��o��gϞ@c����PUk�L7e~n�
+8�ww�8Q��c|����7E�k� �z��%.ȼ��`�S�3��k��9Y��7o��a�Bϕ��zm^3��(S����ט}�ح�����.V��9��N����h�x�:E,7�ަέ�bF��N�ل���������Ŋq�^�S:�,-�I捼h��xA JA2hLi~Zd
�+NO��x
���;(tm���33Ͽ![8tIт@���Sf�1��'g:Ɩ����y&يJ�2��i�a��@�
D�[��y�Y%�/��Ֆ�uV���)������q�
�ss��@!�Z� ˦��g���x<D����#�y%�?� ����;��������7cW�kf�3�Il���U�#�@I��" &n���ֱ��=S�i%�y�|ې�E�y�`��.D51z
F����w��8�ª����$CY���4 ��<ב_KJ`���K�S�v��=�=����C�H�:_S-�F���(/F-�V����y\엹�+��L��HĔ#�y��;�E!�s	ܖ�ȕ}������W���MR�vm����hQc!���jt��rv،�����S�����ݼ.7n�@������!��*)E��0�������=��Ci��Sb*Ul�E	;*��Q��B�<���k��~-~�1��� �}�9iV��Ż�JTH��X��g&髯��'_~.7o]�����kk�m���V���{<|�X�֮��o����_�d	�7���-.P�鶮�o���҄��>���>��F*g���n�	��R�݄���q(s�� ��tMA�I&�!"Vt�sS\�T,�Y��1i	�`�!��U���E}@�M^0�u�,�X��k�5W1�ߠ'�a�7��tLL�H�C�����)jP�'4+�iOL��^������)�ᐇ�^���t����X�<6i�C�q���{��N��-���ug�Oz�P���޾\o8?�Gm�u��y@����P����1��u	�#8�hw��"bp"����%U�bK����T;�;��C��J���2G=g�i�{�x��{���9r��[͋�`&��	��hs�2��鹚ਃ�Y��X�9�L��ް	�D-#dM-����@y/[�f�W�Ǽ��ObKza���Ia���n��JT7/�˼t��;D�Уэ!���s�򸾠�T�_�(R�A\ҨY�JRe}����o���ۤ4�V��Zl�3��^�~��8�3�miMM����������5YY�F�h�z�Mi���k	��W�ްVcivF�|������k��ttۺ7 �F��U��έ./1#
����T�C�_=/�M1LG����jP��r��-YY��>%��)m9 �h�K�,�ȥm�c�E}W�t���:�~��䂳��V��$�8#�`"�g�U*?�1�I���D���:F�Q����i�#̰5�tX�'��j~��3��5&lWhχ��=�|�-�)�๠���c{�FG&~���8�#c��+�y6����s�N�~���5�>ECǾ�N�$Б�����Ջ�b���5�B���.�C䯏I�F�on���d~�Gԟ�L��X��؜v����٩���란�F��1��iH��Cv1�z��ju���{�� |�Y^3\[Tф���R��]<t���HP��բ	+�s3L��Ǩ��yf��D~�7�" �8�Q(����5�r�V2���)�i^t頜Avf�m�S�E�#�f��铇�E�'�"�B]�nn�d-S��Q���rmь�s��:�e�:��:��*�,����{e�d	���G���Hd������*�?��HM���͗���kϸ����_�@����\�.Od��
p�������c˔V=��]c���>e1�ǿx$w�?���=Q�d�el�ˍ�S�z;o�QT8���擃48�žqʀ��{`4�f0lh���?�^D}AMZZX��?��|�_H����E6�w�v ���"!��¾`�L������쌇Q�u��ѡ������ �B�	�5rKa"]}���<|��/,���9#�x-��=")cπYfز80�,�˄<͙�9��zj�(O�#���L�DH�B����׼ެ6��Ţ������oC� s ��O�]��~��i~�Q3L'x�NȦhQ��G��U����}�eEP��k�K��N�z�N�cd�N�,��H3�7$�����Cmg<2~�ۦ�k\kJ�?��7���g X�O��;F9ѵ��'l����:9M?�r��������H�֩U��Νe�,�6��bznE�
�9ǡ���.�򷺧��8�Y�psj^ߦ�`�
���wh4��8AEA����c��o߽#�S3��`$����	�N����\:WX�D��˞������H��'ء(� �{��q�4���(< 7i±�Y�i{��Y�1
r�0���m����P.ҹ�2����_�����\^on`:r^}��P8	^R��
M��'ۃ��2I��Y��y8��z���A�0
��t_?�}y��-R: A%B�>�˂Ƃ<�ˌ���~$��{DP
M����� b^Up�~��<R{�9:�̨8�x�v �q�����")-]�ׯ���*�e���|%/���A��/�ޡ_�@���\C�=kru?O^�@�Aݳ�$�����D��,,�i�#��,2��^	����y	8%w��p��J,;��T�h�6$e���yb�]qVH	�#�%y�If³�3	.:@3����:D�)�	�+gK�z(sT��~!!h;�p��S`]g� ��R����s���Jb�����	�k������X/�1H������6����5^�Y���P����������@h1��]])5� ๦S$�wH�6�AEvSxy~@ҷ;�����+�?=m���au%US!��g��k��{!�8����ÆѫU�M���������2-�*2�O�GD�eq�Q
����`,�Z�ё�%�=HWƒ��UH}Z�D��D��	��2?\����G!��JcA>��d\B�y:�k��0�3����_����&���t�?`������B�8Ac�i�,�u)j���U�)3�H���{�n&����%��;R���O%t
�y5�?�E!�I����+`�CN�Ul�q�����G����o�Ӓ�(B?�n��ԫ�8;'PD����U�S�_�dafJf]�l��2�\�aRYK9 �w�a��R4,�k�xM�UH�Bv!�F�ؤ�V�W�����C1�������_���4 ~5��%��Z��d��7��;w�0j
J>J����}�zP�5z�^kHf׎hw�s��Z����ˣG�;�k���?|`s�ׁH�	0zÑ�	2��� ����C=X_qN��T'�"xz6|��������|��|��T��'M�ᠷ���hĴ�����%D���K��10�M����Q�%h#N%l4?�%R�������<W�G�h�5=�٥C䑬��"�)�A(h�&v��ej�u�=�6�t9Ҵ?����/�z���H�:�z��]�Êe(-:��@�N��g'�Yz6����;�����$GG[��u:T��zc�(3N'�]�c�����g�GF3�?>��~_W����B�0��poEf�W�c?���K�~4f��l���"��q8P��|��t�^o�������� B�u|&1b����Z�{^}~���hbxI�BW9�3��d��L�b<k�D�Ƚ̝��`���33�\_�55w&��e�K��{r��J6&-�3J�P��Ӂωc?S�+� �������w:n��,@(Uq2�!DDqp6�'j�O�m���a�]J[iK�M,}��`�ͱ�%G�y�Ƭ�]��� ��
ur�E-Lݚ�u�a�S_�,���A6*"Ո|�U��Sz+��4�g��-�[[������34��9=����5�G�<ږ���C�4�򳾶!�n��� �㌪���A[T0z�����:OM�Y�`@�g��|��.�\�0^lM<aiز#<t�= �{%���c�¬UX�E�M��B<�}�Q�o�xB(�XW�N�
F4�2�X0#'��8��f�'��m����?oٞ��)J'�(��t�4qҡ0�g�Q�PM�9�N�AVuqaF��_��z�NU�*2��{2�y��h^�����3p���L��.��2�Mc�'�<������i�=��A�����-z�陞���Ũ2Gg��P�U�óy�rڠy�R�Ƚ��G��pX��	��x�|'V�R����I�_R��B���xT�/��J�=#�H����AН�D,8D9,e$����/�/CO
{��A�RTٮ?��
	��N0�6��DQ���+oJ��I�'X����4���, -�+���8Ǯd||lU��{D|��L�iS�j�`(�^J�6������uK�M���-�a#�s(KK�y����$��3 ��r
��O�qV�������݆<�GbQw �j��1�*�����;[%���4> B[�o�po�E�P���!3
X������6%,3�v@�׊f
E�M.u�+�u��yD"�\�D�3�-�("r0H�⫮@�ѣǲ�"S5j+K���Nƛͷ�Z��~ �_>�B�c�س��0���������jf���0��=ܿx�H?����)��sq�$M}����(=�3�B;�&]�+��ܽ{_~��Oeiu� o�h�EC����0����QC0���g^�f|���{ţ}��	S�z��ǹ�-�î��ț�]���odw��0����KG�A��	��^'����D3���5gV��T�^�x�'� �5.�z���!0��4���:�zbk��$	�?�mpm���g3Z�*�����1��!�[z����@���e�Ri֤�׃��|pfR��w=�f�x����(H g�9<:�u� ˫��`*��^=�5�g\?z`�A-ﻹ�%��_��W��P���ѧ�rpr!���4fd��*X�{��^74��S2E�_�hHuzv!��[����k+�n���3[m��uD�����VxqhȄ1�RzD�=�
N�%M	?G�۬��[���6yL�Pk��e1��'�p��qF�����W�vdt�ȑve?~ݕ��oO�
'#�&���[)�t'E���n/�`�g~�A	Qj�
=���e&WнB�[1����p�X��o�''�{���klX���H�XN�yz~Q�ڴ���쫭8<� ����'ǒ�������vp�[�y��&��u}�B��FDqdՠ��3D۟3���$}�,�3�v���3H���ޘֵ�B�����Ç]Vf�sF��;(q��l��+��}G�,��ʧ��r����;��p�T�x'/֧�bs+t��A7���i' }<��c�&Kh=OR+ %&6Y�C>HK/.s�DC	M�x�"�v	��C����-�l�]ӑ.J�;1��8n�$3��E�郦���oШIL��jbAX��ֽ�"%�5"���*ȕ����
�U�������C�*@m��P.�v������l,j������Nw@JV���Ә-���At�\�i�b]�ѱV5�ah�����-p�gR�-s��\_����^?�Y� <z��%����u�h"���P�����̫W�p���<~��5����#�9���|V�P{sxYd�r�s68���0؀�Ӑ�,x�|R O���H���%`��G����f�HF�.bxNd��l��~)�B?
�d��,e�_d��]�F��8�8����f�k���V�(/}fD�kp2ʏ2 /SYʿ+�M�]>\
J�H���8!�5�U��t91e>�y��6��`�E���޴t�9�&yhbzs�AKp��_��j�J�se� t�����BD�� W(�^ĂȪ9}W��Ǒ0�H�㠍� ��ٍ(8��Q��˗L�>x�H~��
��02��"����N(��|�����jh� ���bV�܊u-�zv~���~���P���[���������{ϨD��x����Z��A�5\��r�:?ssr����������7������[�zlomʓ'_�7O�%���֥�Y�E|vv�ءy��[Fn�e ���O���M9փ��>���3��*�l[/��}��G-��a\�,�b�g��tzcW�S�
� �l��kV���Yr�GzM��s�{ǧ�闵ЬL�I]�T1b��������>�
'k&�29ta�` �U-8/��3=h�l��`1�_&u�Q�W�,/ƓNgb �"hC�)���t���P�����N�C�>\(f\+5k�n���f�wx*�L�:&��҄�kk�@��9�"�2dd�T8�NWF�mi��O�� �{tz�u<*�W����hT����&o�@Ҕ�J4/+f9P��;���=]D��aᶍT���L0�[ó|俋���~!��p1H$�c��(�E��2�̓�_�ń��7+�?��⬔$!/m�h�Ltf� �C��d3h/ �p��Z���$���ĉ(����0l6eZ�FEQ[���ɩ�q�;2��"Ss�Қ=ձ�#��.�v��#���=���>��կ���Hsf^̖T� ���л���PK���0#����.�G�O��+�ktj�k:�fY��������Q��OA��%�-�Gg,ć"�O@�E`��h@{k5tAP�8���:�0GW�d���J�x-��&t��eՙ�PC�F�͋v���]��눀gG��:|���B5�ޓ�c�w�jOgb���SXg��	��B��_�!ͭ�Q�<1Iݸ��,�ӱ#�Z�Vӹh3K�0h7s?�
b�|�@��������#�K��l܉�� <W��@�P��E�
��ծg�Ϟ2������h���EF�TBH�F�r�t�(��5 d����"��:����о0�^Э��3�������<It�`���ؠL/���	��47ó(�1��4*��b��J�?���|Nt����\�A]$sn�ؼphֈ���؋بӞO$� �Q����q�c�ZʁONZ�Y��Ǌ��A��P˿]IGF��b<��G^К�q�au�]6+X����ش�'VvB���gE�&�U~PkݳD}J����0��6Ktx(��%�%�Q�*������,&3O��[�K��2�%�~|�F��<p�ý����3Bi��α�&4���*��3"HU���pQ��*����v�VL�����P4�h7@d�/x��.V���z �_��s�	�l���
4�pO���A�A��7ԗ�|�?��(8��d�N�O��{��:3LA¨m�퓓W�[j��T�ۡ�!"б*�O+:��AC~kg�RF����kYZ^���3F�1B�v�qx曛�4��Q�
��X���B-&�~�h���>�>h"rx�C�6���9�g��L+�r�QQ4#���R�bh�����l��	�9(ᴡ��m�-���<��ҲTI ��4gl:��C��k��{+vpd&��ƽ���#��A �5�����C�� *X���E�r�鵠�#�κdF����?���'�LD��)�=�~+��{�0ݔ��5i�A����8�4�8Ǟ����G�˔s,sD�O;�?��s������OT�l���Q})'��]%.&\2�3XC2���=cm�::�Kl�˧�^�0m��Q1���S�<��â#oP=B���S��a�M"x��U���=���	 �y�z�V29���'s/!L|QV x�%3ϴe&���@4��b�^�؋l��>#��Ix��Oˑk���~�f&%�
]�����-��P���+��ƥ�ty�*On��g�9ad�=(#h�c���C�w�P�Qf��T���ǥ� ������JbDS�q�������W�[���k��.�����t�-��l|1/�fF�L�: E�!;�3R��<{��T>��ܾ}WO	�@��=8���s֝ �s�@u>k�6����Յ=Z_��g�H�t�]�Ê}rpt"+g
4��o��oI�h�ͨ��V/�ً��2��9kF?�.���s9�>p�i�R�X�=$�w��2���t�ul�5��E���=X��y��^�����ƌZgY�2�Q�b �~t<"�웃�;�
���B��nŵ��8��=����)/�U'�Biɪ̪#�83'�(b�[�s�;W�}xP�`����X��uZ����io�����&)P3�9ڼ������p(k�Yݑ�g$��1�g�Q΅�� ��V�s�i3���EJ��{T���r�N+�zQW��:�`D)������G�<�1�:[�D�t�@���*����V3^oT�)���+��V�����|N�����.M� ;G�<�m�5�Sa
i�̊���%�G���/\o����Qh&3d�X����"rjCH�ą����5� ��#3!�^�I�5l���BJdx0.5|C4�ء������	 ���=L~��&�����Qm��vh"<QZ�Nd�����ţ��(s�/IB�(5e�<��n�/�ġ`�NH<���|��<E���v��c[��>@,hK)b�ν+x��[j�6�\�Nh2n���y`C$�Hw!j�Ѵ�so�n�g�WW"v![�{���N�Ls���	S٤O�G)F�J���36���������}�`Ȃ�`|�>b/�@PH�L��B���	�p+z���u�T ����{�����bt=ͨ�+ i�`��Z�"j��-&������&]��k�?P���k���g����:n�������+�~�[]]��������_���!��(
B4x��:��:}��'_����t&�����T�|����ZM9�C��p��tQu*���Mc������c��Z[]���Ey�N�t�8�8�5�f�T����*�*�@�fu6u~*c=0��J�^I��}�u{亿9:�ZO�#�h�9^��æ2��B���I��i�`�YA?����jI�%���v��� "q�]W�1�4�X| �FS��UJ+MET�8d,�B!R��Ѓ�KR��Ss�2����	)tp_���Nˀ#���5���Y�3h���fF�B��2��D�������۳P�nϐ@�1:�$*�.z��4c����^f� (�\
jd^ ]Rm�#�)y��6�����Y) |HD�lu���ċ�="	�5��oB셳�q">��2ϼ��P�߉�{5�u��c�4D�%s{X�b��%��ޣ�ꙺC�Jd�e�Q��wt$''엁H��鱼�٥Z�;�����ݑϿx"�K��XB�g	�+\��j�j���(�^2K��9�?�3J�w�#�J��"�U��lm�Jq��ʭB1c�v{���p0@C���YG�>�`�L�FfwAꭌ����Ky��5?TQ8.Rr��kΕ���bdq]dGd����[�X�A@��A� 2{�����u��<�w���\�!(}EQ��[�vg1V����Z�T&�Q)4�ǹ4�4�%�>Mwf�3:�_W����\:>ܧ��Tm4�07a�h��I���>)���V7�(j0��m#�ҧ�v!��`�f��u~���,�Ե��Y����X���Z���E]{Q��
�O��A�.�S��;�
7x���1�O�����?��<긆˦����_��vZ�H�s�&b�^E�S��#��ōZ2u�7N���v�<~:?4C���qfEU��RK "�0���`�	A
� ?5�Ġ	kȚ�*��h���a�sn��w�`���֍�،m����8U���(`+�>୉Gs��o�	��h-�T����&l,�'�������d�[o��I���p�y�X�*t���������vG'yZ�M��%T�P�^�u���g�t�o��v���Z��i��cZH�lԹ ^�Ǒ7��,����疔�syPF��4.pD ��0���L}����Q�
���V�A�� kn�[�Qg70Q���Q����HP���^�t���B�ok��)A��*����a�����E�9Rf�,��ql�����&c͔���F�PЯɌӈu��* :9<��J��������Sxrzvy����zPJbkB�5���������U޺y��ߌ�{������(�}��\[ې�/^ɗ_~���`�|GWD�͚<�O>zO6w�dw[�ɖ� \>|�ܺq��z�������]�ei�Y��� G�j����������� ||��3�`%:��� "��mU�dE>���W/�C]Y^����Mb�� �;���o���P���2��R.��L�;�T������W�Q�"&�l90fVg���v�ϫx c�-���:�(��u���kKҪ���f@[33� A���E�k{��C��Vq�6��=�����M�z4�Qy��X]��o�|�P���WLǙG�]�$B��zx����ࡪ3��d��Z:Ru���:�8rcz������Fi�ZF�����V��t�������r~�jQDp��	�S�%<��Ƹ���7�zV�����$�S�T�FrEӰtT�r�'ã���#GU���N@�?'�"]f#�{s��a�&�*LuN@[`�0�bD��v��b�$=�L))#P�*����"]�H.p�"t��]1	@��W�\��8Ig������~։����aA�9��f֔����bsS�;
����R+���峯���;6E,֔���Hz�{�ȧ���%�!�P�WF�P(��`i��7��տ}��Q( ��;���l(R�,��� >������R�B��C9�j9*����݀4)+z�g�6��i�ȀI""�r�,ʃ����<;�5�� -�#�On:���{14=��/*Z�gQs���^w���O6hyi��.�{���q�vz����#�aG5�#zP֫N~��&2��N�86;=�{:�qe���������3��zK�ՠm(2�Z���c�n�s]�+�>9;�� �KMdt�՟��2��/;����E�:�./-������\$�E���ݻ���f1��2�#�+B9KАX���.��ӳ���� ��`1���7��/>`C���_���8��z@����F��H�&%dKVdf��뱜^��D����T�~�����y�4��y���yA��a� R/�ܨ$}]���Sƌ�'�g�s{�����1���Z% ���!)��	�M�&D�i/	��"*�H\[_O�	�l�`��Ep�G���O���p��P��ʹ�WogYAPY r�D�Mā�� �Tm��E��
8�я&���މ�A�#<�k�$&~�xp��G��a�o�1W ��'D�&�ҷ�X���5:�$�M��W�*~���y��G�w�C݋3&&l81ʭ0��Vk��\��pk�,�ET�����eF_�N�<PY!*eaʏPa���8(�KO��ޕ�!vV�����$��;]�g�G�J�Q�ן��K�cщ:�%�2��d�rqr��i��1ދjT���e	F�N�y�f�
-]-8�}���}p��&p�Xs �aeiQ�49�3�Y����/���[g˚��p���#͎!	�k�-x� �il�PL�{vhL��,ca��ZB]h8r���H���<Cf��L
DONԡ�O�ļ���3�?<��s�#�P#�5���=2�ئ�;�3���"7`A�*�ɤI~�+�Z�:���	�i�vOzޓ�S��8���/�٣@����BwQs3�`g����ЬE�|v��L��z�
�O�п�#��u����ֆ��̬PA�}��i��4�`Dti=�[��^O��'"	.j ����8�yAu*jg@5�Ǚ �p��p(����l�9�B~FD�}�]
7w	a~���*�H���|Ϙt���@��F��������	��&����Ӆ�K�F��u�e���kfƖ�u��J�m�Z����%n���kY�c�����q�g�C��؝"�s��ѐkO(<9>�`�ӼN��J��m��W@���SF��b��� mt��)���;n����ME%�]�E���e�4�l�����;tp�=#U���h�x����mA��3x��0�e���t�S�!���<�����@O]��,�����c^:UW2��F��C�*�l�1$]A.���^��aHB��z||ȿ�S�}a���2�Na{C�;D�����{435���M(�zZ��X,h�����xw;�����̂�'rt���?����3�,d͔�,@v��ؠ��&u:Ī{�Ě�ϸ�>S�yG��a�����;��٘���e�)<�Y��b��f��GM*3)��j�l.���Qu��}:�����0gd�0$��I�}���G�������
,~���W�F�	���8Wԑª�Q�T>U���^Ʊ���g�X��ˑ $u���6n�,��H�����'��W�9��}�p�R���
&*�e��7ڡ�A�R���� G,�µ0�^�p0�S���#�kT�R��?ϛE�'�ha\/�_!���y�+�m����͛�������6��y��_�uD=�́7	�_�o,E�����G���+�IQS�[h�`�Ώ�*��es��B������;h�
 �mz�%���DP�=�H�g��������9�+��n4Ś����u�:��١&���_�Zn޺G�_|��D�%�%8��Ǥx���0�R*�����lPl|}� `-�Ҋ�p�
��+��8zV@��	J�Q� @��y�0�H��o脊ڂ����x~~Qfg��8"�Ř�a�G��sR�iɴ:;#����Z�w��F xD�����t	�� �(���y�������LG]���t�<\�M:e��A�-��t�XqT.�Zu��C[���-�=�`�
���fSiQ3�hІ����#�U�!���j�FRa��J�bdQ@�|{�%o��8����T�)���oυ���vO�iS�Ss� ��F��9�aH��Ҹx]��b=D�
��aB���~�����z.G���bI=���;ΝR��x]��Ԏ���gl����Q�����w^Z�7�o�����X�βB�,s�
��X���T������:A�DbR��Lx��+)��Et<��=q}��+�t�td��|���p}�`㉖�=!f�&P���R��H$v�j�~H^��L��]BV@yd�Y`:�9�Z8e�V�5�xC��x3���>S>�8r�9�6W�r�7 BԘj0Cf��51��N�{�_{��6�U�I] �:JL�w��~o� ��ةE��wG/;VC��V��A`7t���&�N�YMA�.��P�;e�Ta&of�����Y)�zHJ�\b)�9p��H�ߐ%���b͇o"�\�W�L2���N����̜e_̽žs+PW�x��g���Q�|�n���3�b�4c *�)dS���<mX�<X@��#��I� �E>/N�ɭ7U����l��eg��$Ŕ����5mg^��/����������q����Թ�jt,{`����i2�� U�ڐs��C^���>�|Nsz^j{q��n*/^o�\m+b�S2���*?�;9�.��R�ԑ<aa6�n6�Z�삝T�1�3=�W��9Z�CS�1�7h�c�7N��n�������.�_|a`�b�?4b�eB�N��I=�f �Ho!]GV�	�IP��!�}�u@�(��[��Հ�q����e��f��B��? �y~n��'��G�d�?����&lrG��yD�uU� !�)����1�=���o��^���[E�7���*+�_��<"�
�Z;��X����ws�gϞ��RQ��޸�HS]1�"͂l֞�h{��L7*o�/4ϕ3�Ru�j�W=-&ii滑/���$�8�9�nD������;��zW�ik�ƥ�����yE���z��.櫓X�FpN�2��_XQ��2�h�ɳ�rycC.m��nn�^��O����?L��=�גsx����믐�!�:�܃k7ȼ\P�+�w\հ�#���?���a���=/�}=��ݑ|��g,@]I�%�������t���|%��T�8�@�<yy@�����K��t�y�(���j2%*u�����9��Q]il@�~��������xN9ɓӣ<�����J�h'W�l��z`?���4������Ɉh;e!���@���� �Y��&�.���Z��멇<G����*��^�*ZA[1�ӝ9�ܜ����k ��8g���l}���%���S*h��$ jԚ�T����M�vYFؗj5��BL���؈4�ds7x"Mv0�4f+�z���ٴ~���g^
�%��DTQ+� 0���k��YͲY�,Y��§Haۖ�Sjgj����� |��/kR�����Ŕ��������V�Ih�j}�
�k���v{i�ep������ֈ>��D�0G��d�s�RЋ�$RbO<�^��w(�Y��a����0��%'��q�.\B�+��g��L�se�G�,��	�n�����ص��:�n_iO�x:`�UAa�T�*˶�v���˃V�;y�� N��	�斝?�ƪ�)����"X�݀�=�wb�P��ea�&u�P	����Ĭ�r�33N�{���{$�A���VJf�S���0��o���jz�:�͘���OYVF�+Ie�w���Hs��5�}�& 8��zs���Ί�9�`��%��.�
�٠E�ߘCpT�!�3�U)렣Jr�c�-�k�����F�f��r6kk��-4#��s�5{�@1>V�>9���'�b*0dg�S�;)-)�  �`=�"N%���jW�2?'�(�����z`�Y��V�@'~���w����:!�<�kf��L@��a��4||=�줝{c>�}p�����ϟy���Sy��v�ֹ����<9ɓ�y��Z���}Yvvv��섺Θ�8D��PS�P��kUs 7����ry�
S,Ϟ?WjIl�}+2�HԥV�<P���M�9P����r�[�Sh(�({�Y��-6a�_�mn^�_X
����,��a� �`�4���˂*ɦ,��Z5��ł�X�h!jo}\�����/����],\��������XfT���������XI�b��M%������Gl��~�� �.��dQ��y�8h�z�����/��vt��g�F�H2�5���7�P.`/\�@�m��v��Xsh{�Nej��vl?�v&D���`,x1�X�g��R�⎽9�N���%�>�����4������՗_�9�+��o�*O�>�F����F�ϱ�9�BH\����Ϳy�Db�?X�����P��)) (��=�3�tQ47�e$CU�d(ee���}����J��C�Z��D�Tz�x�(��Ҧ:45�S�Qjj]�Xm�T t�T,PN����%�ZiJ�Тg"�@&�ϏN�8SE�n4�
s]�.���傍Q`hQ0�u	R�o��� F�9p�af�����q$Zؕ�=l�MQ�����$K0Y���lE�.7�t�<or��L��S�f��e�kP#C�����~^RW�1�\��K\g5�Ƽ�e@!��U;_��"7?
a�=�]��B���oȤT���j�2'#+������X�)��)e3���~i�MM.4X&ĥ��sIWA-��AW�h���hs�X}͔���F��l���b���н�.��E�@A�C�!�G4�tTk���e̎�]rܥ��:AF�ҵQfr�c�X�k?���i�j�whh�e�؅7��^a�7�֠�����3R��ڴn���̞?Ls��=cS��)7VJA���S6�c�H
6�w��.�#X������ ��V�n`�8^��*�����R�f+*�"�e�0UR�;��qN>јNy���ث��Th��Րt�u��\�Z��|�Q����;���ؙ�**=G���m�>�Q�ҩ`g��� �� ��R�2��fȾ�w�����ʁҳ�	K ��S� u���u��A���<;�ʳ��a��}dm:��π�R�z�T��41[G,��t�OF�v4�;�?��`_W�5կ*[�v�̮�� ��e ��[`����6����fT̪46X�)(�����h*Sf�:\˳X]���g����J�_w�'z��v��T.v�MZ�r���?~��F)q8�ׅ2s���CC��1�͑'�0����5.�'Ϟ�2]U�v��K^WM�aL
��p�@@6	*x���i�����d*[�?���Ÿ�з�e�X�h�p�^��A��1e�XT�Wv���[��s��e�;wBl]����6r�rhzJ�}nG�/����57���� c��"k��rp2�<��e1�V�5%W��d2�w�^�����v���>�?h���8��;��^�J�G�Q\�7�4[�~e�sY��c^�����(<E�Q��/r�s̲]�3�Q�b�����~��W��'r�6+��'g�ZhT뺜�+\��&�R�K5|0�pn�Zz��'g�G��+iL�eN�|2�(y��&*�<4����6Y]��r�O����
�W<�Sts-z�(*�S%1�a��I{@��3D� m-�7�:��IG������;���/G��p�}���t�̗e�7>;���Qtc��|���)㓈�.�xT{Df7Պ�ksɢe�u��:��]D����7���"�ֺ�v�#�C_4�pSR���M΂v�����9j����:b�qş�C�U��p!�z�~�%���^��������?�K�kQ��Y%�q@�S���7|�k8���L�)������m�i�0�P��2 �#�-' V���\*d��/9(+�v�!@�g�Ҡjw���|������(�
�`յ�Nޥ�!8A3M��V�K���Q"JRYzt�p (���&Az�K�9�Ut�T��&�r�2d�Tw���e��>
H.3\�8Q��Q,B53������/�L4�$��鱿�L&�9�����ҷ���/O�>M�%;�!틂W��6����+��NR:���b�̢���
`�U�� ��V�\�rW:�L�f��x��ǜ�&`�,�lmnȻ��&?h�˰���`\V�1y��9�>6��s^iT�d�SC �T�jh>�h������3XB����r�k�`��,��vx �\��x���ҡ����y� ����Y��l+ӹO�L�}�x B�n��F^^��S��t�o:�/��Ui𼓛�f�mP��5L�F���zM���ْ�J�W₰�UL���U�Q�lS�W6em�ڢ���ow�����׷�����46�y����02����T�ͩJ�����٩��д"8T���{�a=<<VT���1G�(ba@PW���Ry��:���-�پ�3㫎�Ts��KS���ȋ_�mmi0}�&sɿ���jT֪A��Z��ϬL�(L.(�'E�<�e�̛6�et}ّ_����3K�m�ҘQ�^$��6-'�$K��M(���(�84�j�!��s�ژB]����ޜ�l��5h�dC��L��tK��"�7�a�B7�P���E�uv�З@��w��4�e�2w���Su�2���r�\���.<��~ѣ���e�{r$��99ܧ��� "xb�;��:��v��T��k2Px����"Ї�s�ӯ�ؚ�0:�����ʲ,�.]ʇ�Twn^�׮�6�믿������vsPJ�ٹJ�/=��M&�Z��֠>��� �^9Ę�hi� �1-r:�p���J�}�ϭ`�.]3)��FjME���u������j�7ի���Mr�B�5B�5�r�K�vP�v�/��^>�����,c�=�bۡ^�5��M���#Ŀz~�2F:�o	P�~�fխ�^p��7�D��a�u~��5�����[�%����aM�7�\��Y�G�~���fTQ�(pa��Tz^X�4���l��B0�U��z��I([Y�X�7l(K:=X�.ZL)���l�,ՠc�
����2�5�k�/tZE��$��t��I���Q��jB^����5��ƁB������-ȡ3�)� sP�k䰖�Hr*+�LB�S��؄ϡA���qyCu�J�S�P� Аjs�q���N��G#�+�vTecM6�ާ�����I[m��`#�ֹR�ut���R�Γ�Y#a{~͹_��7���P��?F,��-�w�p��Uh�k��+��^��VW�]���ճǤ&����C������W*횽H��OԈ88
�h9j'���Z3�=?���i��
m�`u��琀D�aT �		f�Jұ�?�z@W�sp��,���W�-�x��.��6�y�;�a/��  e!h��ٱ ����C�`T���rL<؈��;�������Z�ZY�Զ� ��.�@�Ne��1�vd�Z��u7lNO�6�祩t�����X�a�l�p�1��AɵۥA�"�P���#p��e�-΀�.�����{�! }G ��9�3����gY��f�H��Oβ�A74�mpY�2/.,�}�QTb���f�Z~`���ֿſ�/�N��� �V�"��u\���7"d0�½�'��]���&�\N�倣u8�~�E4��Yo�3~]0�����*��'�ܵ���G�m��pߺy�����av��rC�ӣzM
a��D�:&�7�h�T�K�yV�AܠL�lm��#�C�޴}u��2�Q��_<��}�V�v���6#t�_|��C]���S3<��Ε����<����Aw}��bt�"����j���W,������O�@�Ԏq'{�}��d>��Y��C"��WWtjpis�˿�K����tz��W��|"/_�����}�����?gG�޿�JN�����2@G7E�Kv^� ��V��`gD�h
���Pg�_�+��n�ϧ�:��r'�e|�FeoqGB���AE~��Vǹ�Q��-��*G�C�fD=�ج�mR���&��>u�2E�[�����yn��V����x����Q�W[Wd)<Ho�a�t�-mOh�����ߧ/Z���]ǆ߀hB�]:A�I�n}e ?|�����0����"{/_��5`g��NF�q~OL��c%U<��u�Œ`�e����3Ed9���6S@�/Ź8eC�Q�Y�f>���VM�:T�����Di4A�n10��P�tޕ�ishp�T�����L�W�4��y펥5@��.��N�4�a-�̝�%�9�i�E%�)�#�W�]6$���x���Z���5G�q�`�@K�Gɱ�[d�CuxΗ.o�y���g?#h�z�����,'hW�ݏ��ة�q����׆W۵�Yǽ�N���&�bt�3H������1����Ԧ��W���Z�)-RU�l�CiY��W���<�+�]u��쇅Q�)?��KiH9�z��t�i��z�u �aOk ���
��C �Ĺ���D�����UV�q� .X�ó28\���[����m����9�@۟q�3�66��JF2{0�X��v��{�]�U���w�"��y�`li���m�0�{�J8Tz�mN0�/_����W��ԝ���������O�]Y�΁'�SS��N6�m�r}bh�bc�pϨ��V�/4O3�N!`{q��ƹfg�����;tQ�u�-*�ȱ�L.�����{�$GakK6/mqbaa���T`��Лw,;�f�|�/غ�Ty�ѹ��Vh�`z����rJF�ݍ����k"	0�(,�ÿ��ICF�X�j���R)/�Q�W�MѥO��\�8���e
M{sik���\�՞�0d�xj^��;f������d�Ń���|�P�/���Woȓ�{���n3:�Ug�yN�|�Tu 8���=QחEIB*Doed���E��!��H�B�z/@d��ǟw�U��{+���!W�Ʊ�Ti3���,f��T���ra�b�"E��9&,b��YZG[[��O$������7�~%?���Xd�s���M���ﾗ_���|���i��hk0��� �?���ʻwo��o����_ȳG���h,��ca����
��Lez�) `�|З���HNR!����v$�	�?����ȟ���d��@��O$Y<Stם����y�<��.�;���k#z:�Zo�M���˚hP��g�}
5�;�9��Ҏv��%�Qm�˨a�7�R�J����j��� gS9��#f#TB�Z�����\�P�Ӟ;�%��aOS�h
�*啪��6<��э$��%٩�
���D�̳[�0�J7u4�.�\�X�s�~QП��lG�h1�;6�_(NCa"�@JW�k����_��G(�����O�W����4���Li��6��Ɗ���W�R� �ԫ�d&������ܶ���.�d��bW����BvӥH�`(�Ҵ����W������D:rr<R:@G�Ng�Г"q�o�/�K�S�_�p�_���~�F�1e"o��ζ߻m~3vE.Ii�$��YA[��,tia$�(�Y-�"x�ME��70���F�Խ��x_���A�/~�<x�.���/����}m����xJ���јv|��[�=熂�*�m.B~�l·���\VE�� �	�)��,W��(b�N�Z����
R�0�k�K-�����P�t*hģC)��j=�E��Y�6��:��������k�yS����1�2�ݻ0�֓���<��:�-'/vu՜Ϲ���\� s��������,���F��WIׂ���]�4�<�@(kf��S���2��[@��(!�0 �"D&xw�(v�*9���x<
'���N�u{2A2���	e�+�[����Q(�a��h %Ȃ�w�(���F�͔����v���@ȭ�M��x���A�'+ ������
bZ��Q�%���z�����R#���՚z�2�iD�9ܡ�b�Z��9@AGW�q~L ����=馁[{�ard���0mגZ��q�c��ZϪ�t_�o����7;��[H�0q^,4&	|�e^�w�E���1�'�\ٹ&k��P�WdecK^�q�F�O��4�����C\����sKI��Q$ӡ�cz� H�K�σ��N}{�&�{O�w��e8K׵?�>�����7�ޓ���!�/�˧ɑ�	:��n���=���:����FVT4��]6^�lI�����覷��S�NR0�����Y��m�A5 )�7uU�H�3�17�/����ƿ9�����Kr��=���k��'(��kz��7�Y�<pn�5�1���}�>��P�j:2�rR܅ˎ����cdP��r��_���f �G�-�^;JR�F����ưks(6)���|�Dӈ��8X������T��K��m�Y��$K��"��bǿ�̩
	T�Ptm������}3+Ϧ#P�6�I=R�[_�0꺐L������z�>��e��8�� �X�F�i��#�������%��G���~+�|�{V��R�UDh�Td�A� ����5���FաU5�Nvl5�Z�u]Z�:�'F�CZo�'��'Ɏ3�Fez�u�4C�#��K��Vx�M\f�<98}6�`ɛG0��v;�Q�fE}y:iZ������`��9�cņ]��R]'VJHm �N�q�u��f�$������ʬ�����
k�*!��$�j3��߂�J�d��|��'�q�s�q������Iec	4lF����K�<Z�t���|�<wD�IE�>k�k�UѺ��A�'R4}F�?�?NVp_e{�-����t�Sj�A=�sf#d��?1'�r32�0p?t��|�>�La� -S�m�u���@.�Y50�]({�<]5�Y�9���bz��ϰ�/�(�s��1�m���F���Cs΂�xD����d��x�j�w֮�zA�ܬ��`�9Zߙ!����l��� �s1@*M�AV0���_k����yTj�%��8��'�d���l�0.oG�}ڠT֔�=�OU������Ρ�39�/�8�u�㕳���.��E"��Z[�K5�h���h���xz�`��jף�[*%��7s`��BiO{ٸ0��d�����q�(4�C�dT�]�����mH�Aeww_������C��+W_��/^WZܬ��jCiu�-�fى��X����j߿!ˈ��y�)=�e)�t�P�A3��Q�����iQ"͋/6�)�8(���t�،L�fX�$D�(�ن<Vˑy,��D�a�}i;����s֔�����K�Y�È
��y�}���լ��s�.�|v}�[x�Fg��ȍ۷����˓'O����2mZW�F��뗻r��;��j�֎qͱ�tkx���@*�L��q���S��gr����G?��E'mt�~�FP�J��k��dt��ʣ���J���o�;�d�}�JR��:�����Y���L�&��k���?�����w*G���S�Κ��k�r:�s�>4\g5A�"���YA�_+�pX��1� �#� Ŷ=-��$Y5I���w`gT�R�F��˦Fu�Ϭi�g���ײڵ��P�ë�!�P�4���Hfgc>�`<�\�UU��|u��tO��韝�I�{Y{S��$k��*�(Ue޲M����1�F:{J�R߷P�N���p�h�����ύ�$F+���!N�_O6��>�P�mo�������]�.��p�)��,fCѼ�4��&C��h����v��Rg��#�nf���7SitL�˧���j����aF�:�%�?��\�G���*����5���Sf �Y��@�ur&Yъǹ����h:���t0TA��Vqnh��`r��0�=�LN{eE�� ���GmU>v�,u���z����(�]I�w��+��g��Zr��\�&7��ȫW/L�gJ�M�������=	�}ȳ�M��������X��7
���.��W��b��`�l�;�J	SIS(~�ٕ�͈k��s�6������&4w�ךv}�����F����_����5R���=�-5��Wɯ�6r��t-���Ь3���5����� Pk�����K&'�^\�w�K�8͕9R��}��|���t۫u�
D�;�DF�=�.4+{j�����/y/o~E�?Ʃ�^`���J��q�띭��_TJ������Ŵ�ŏKO�r�K����(+PKZ��=נ��Sm�nN���юVlΰh��N���e����2��fsS	�B�Kk���d7��V�@�����y;��Rdȟ�\e��z��W"��w޹Gg��Ǐ��d$�+���w ����d�U�z;m6��p�����O?rA�&�oC��c���NUq3+ۼ�%��\s��ׁ�'�ﾓ�/_R�N&[y�����a�҆o��^���>�V��d?�kkZ�/\[l�%:!�0Ss�M��H�'/B����j��ρP{l��z[�x�X^�������UpvQxzrz&ϒ���?��?�ҥM���;k Nh�dT��)���+��\�Lɠ+�[�r#�˘6�Qr�VS ��{d���a/=���e�0�+BZe��|i�]�/��gi�|����ݻ��Ïh������6ҵ�~�\�?IkcON�QV��lh��:a��RR��@Σ�G�n��V�k�74���ե�ߚ᫈6�ӵK5�~4�]��������!\�cii�j����:9Q��ğ�+!����֍�4�	ԕ̤*�T+����dဲ��hu����&�Y_��1hc�Q��̜u�y��NG�PlV���������=H�lv��ar�gl�C�B�!�;�ܙ�Ҟ�G����h�kuί(}X0���3~�h��~zW.oȭkW9�P������nS���l@&ȳ��Zu�]e�h=�p�k���˄L�W��+�h�G
N��W؞���4ŌnU�T�^:e�N�Q��fn�ϱր��S�t���]����ۘi��'��mؔ���:��e
�}�c����Q�̻�.�~��Sm�G��s���[3-z��D��R��,��!��Ʌ�*�I�X�?�YWY@{�e��{i?B�r5y��6���$��?�4+V�G�1��Z�L�*b�5����l��=:�)#S�h�EH��I�	i"����a���5�K��J��{E�n8�(���6n>�b�C%�J�C��늢�i<����h_�_�\�``~�u�P�`X1vm���,�-:��e0��ݰZ��~��Eߛ��dC����D��#�.�ϝ���pD�:���B�3�O��·jb�=��k��Q�a��.��4���$XF{��^CZ���Uh���S�G��^)5��jm4��{x�#ڙ�.�E6�W��l�,Z�:d��Rn�{,���c�&����=�k�z�!R5�u��*+2��0�km��Q��V��t�]⒍@ju��FP��V�ܸ.w��#��j�ur�^��"2�jwO^��R~��ϵs\Z�(q���Ҹ&i��4�ۓf���ga��7����>GN3;Z�F��c��H�������,"8�����r��=Y߸�{���{N�y�<���X�B���C���q�]����u��!9�d=*�����<���Җ��.�V���i���ؓADvo�����̡L�g���~���m�E�:D��]AU	V�����{�ӟ�9�,v2M��@���X��[���v}纬���N�Af�vӦ���>��d�G䏦��@�����&��,�47n��v]6S����<��+:Z������u�ӿ��㌔v'L�_vsC����Ύb}vLt�(!2P<H�4F�Lж��l�����kr�Һ��iO��_��C�}��Dq���mL���dH����tf�����9�a�j�*��)WV�Z,�����ξq��~����[ٽIV���tD�X��d$7�_��W�5������/�H�oĹ��d" ���P��zS.ݽ.��+�3�u�r����}M��j!s]T:-�]r��a�x殱�������9���ۯm��Um�0�p�S�Zr�6�s���39;M�����󮬯9�Z4*C�H��3տ�-"-������Z��"�!(ͫ��3P��6o1�n��n�(p�
+��s�C%��~�h3@�ĩ���8Ǥ�OZ�E-l3����d Q���D�{t��+Z���і��[6X���`�k�;e�M#攕F/�e�j��l��\�R���j���Zk�إ����w�s)y�A���ZWp`������M�񐙚��ƏҺ=�� =3���|af�y6?&g.5}�p�/V!V\]��¦b�A�grr��eDU$p�;��%�qq��Q�S�[U�<F��C��0Kk   ��'���%pM@|�������P��`���k�%��O�Y��R�<H��ǘte�bݙ�J�
3K�����-/�ױ�8c��r��b�l���~R4�H�49A&�������\Agu$^E��gj����z��!����Ľ�Ӣ !�]Ȗe]ܾ��9�~(����с7�ݏ���fcDu6�-�ϯ�qcE���������!j���S�����=���(����T���9=�!�0Qk����]ϩ�FkH%���VdG�����*dr�2ד��h�A��Ï����`��r����A��ʟZ���>LiҶuluQmm���Bn��EǴ9ܰ.·� ����{�	M&,V�f�5�߯^�J����%�پ��6T�hj�[i47�o��3)�Vd�Ǡ��m�s\��t35�K��4UC���:�W�\�kix�6?�3Z�EU���I:�t�w��S x ��+�c���s��ܼy��ӧ�_�9Y���у�>�Hd��+�������rzrD�:�*E�^��a�s�0���Snn��RC:��0m��k��O�]���)ǇG�<9U7�ߒ[wnS!�k���=�3ln��E��ՙ��(B���A��WQi1V��(��i6Ϻ��ޮZS�u5fC�ڜ�^Z���!=����������u�ɷ_�˯>��`��p�<�Y�~���\v�z��G��`}K^��=b���96�*2p`'W��{�ʚ�������^-G��ɜ�"�VM�<����<����?OA\_~��_���K9����Y��Hze%��=9x%�s�|��{�u���}��{98<�=�|��踈 ����b ���<��lȂ�x�f%���Щ݋T�Y�����}%�c[C����tc�����������hQ���]�Du��}�=�إ�*M-Ċ:�Yg�Zl�<(�����%kQ�:s�(-��ư6�dO�7�su�Y��etudP��g����/��b�0�r0�5J:�χ������+���U�l?����,-LpOu��YY�յ�]ǻ�z�]f멷�U�KW%�fP�cmGcZ�6��1���f���.��P���k�^Z�����Ɲ��Pr3V�x# ��QtPi��9��=0�4�G�P3=9���	P&)��p��/T~����:*R8���Z��B��:*G�w�v\&&��AQW��u�bN᝭��I:?�6��>��k��
+�5�c�Kua�w��hs��M��v�V���J^z-��Z��MN�]�sk�����:��#�#���[����G����(�[h��،�$�JٝW���ٷ�K�s�&�N�)�o�E��׫uiPR<�����|��b\��M��6�!� |r�-��t���&���<�F��tIs4�a�X�wT-B�k�5~#�Z��x�O/m	mTQ)4@�u����h��y@E���d<���0�x �lm���}���\�!��
�pf���~�]2g:��)���cZ�q����i��>'u�4�$xɽ���"'��/��jM�����3lp�(^��Ǒ�R����潙��6tv��j�ئ���l�񀅅J�֬6�f�ir>���"�ZMq�\����c�wD�M�9Ot�ś��� $�όW��2?�[�����gϞ˧�~&�޻-׮ސW���kW(���o?��?����l�Ʊi��iv��Q%����
�t�7�W���{2=9���F����-#�?�;��Cub����/����䣏>�k׮�J�����!Gi�|�h30�pB����?�&��W_�l��iZ��Im��Y���P��9���.H��TJ��B)Tq�lJ�9O�?>�n�_�i]�<�||���t�L������"+� O��ׇ�����\�ܢ~>�x��JeTqݐ��J��֓+7�������ׄ��
Ȕ�X��3�NHNr
�6��ҳ�\�u�`M�ܲs�<�]]�I� Lǂb��r�ۗ�Ƶ�Ķѕ�ar�7S@�
�W���(�@�����;��00[��)D��D�4�z�0�����v
|��,xӑ7񼗴�;&"D�z��z<�I
6t���1h�c �7�U�fEG�4��d�n���S��bi�4<p��6��I�+��kyj7�t��RyD�O��)ҟ��D��sO���� (��uRd���ص�!Q��Q0ϔ�:�>�e�F��K��gi�ɀ?i�V�n�:?K��U��2 �2K��'R%	���7u0����8�*T���dh���rz/�+�J'v-�Q�����M��#+1J�c���xB׺î� *6��ȷj���=�璕Ƥ-bQٜ�˸y����T�>�fѼg��^G����)�Xa0�{B!Js1]�r�D�:�NI�Bh�Q^�?7��a ��E�S��z�n�&��������S/�m�����ܟ�h�[���a��qi�ݞp��;
Pi�B����E�!s��l����EaH��Jz���F�1�9��P�3U�֌�˅�:�R��6�����с��R�aݫ�ުb�V>Mθ�|�"��BŻ7V�\0[��MrUְ&yR�b��!4W4K]QY���6)�E���b�Kﭹ�<JFtB:�!����)j:�T���?D���i�;�������3��K9�d�v�c*�� U��ɘ쥈��_~#���\���k�"8��0�`�r0�i@2�FT0 pXgP[
2.u@��(����Nm�;����.r+=�ֿ=����r>�~�G�8T��C��ٳls��'�@����H�|��ͼ��@������~��lq�莱n�Y3F�d�$pg�735X��s�A�#�:��8Vo�F��ȋ�[y�r��� j�O>��<=�������8nɣ����O䷿���z�J��L�??��(ԋ�=�#��\�n�@�`W�z|tvB���A�83/�� 
��n�3�; %�y���֦����Ç��@*X���?�c�����'���JӃ����*	�b04\W�4_�ܐ�>�k7�3UL�c��Ѵ�s�r����Oψ�c�~��Z�|�H�z�X^'��v|ε*(��P�:Mk��ֺܽu'B�duu�3Ji���z����J=���%2jg����a.�o^1�qz<"P��ۭ�&Õ��j�SR0�v�V�)��,Z�B<��	u�&�v��U�����w��*��D��@>H�y?38'��^	��(=����I���S���w�\Y��@P����'�4gC$�Z4�i�(�.���nv��Cxp��$6=Cڎ�ӑ��`s��y�䕂F���٦A��0	T)Ȧ ���E��������DGs"F�i�0d~:Z ��dGu9�_M���wGHQ�5w�f�u3��;�H��Q&s��Q2�p��]k��n��4;�.�ǻ��ĝ=��P9��u�ѷ,���ڶ9˪f �)�T ���*� �g�{�V �^/�O��Be�i]M�z*(�� P\_X���+t��Ѕzb�۸�i�g�L���ͬ~ڃ{l�U��ԅ�XO��k2-4��j�&!�b��w�i�	�8k��I
$�err$��^��Ds$dvF)@v�9�(�:Wն3 @俪j9�S�T��d��S�������,j(o^W����3f�2����A��V��1�i���A+��ur��VG��?�s5�m��|]����X�Z$�6C�o>�6��6���Zb�A����a}kn�>���,eY��	���Z蘭�Ѐ�>g*�ДA�����J鬱�4���%I�TQ�?́O�:��n��WQ.
Ʊg��H�wj�'/�W)�A׆�:Ջ��i+��=U�Y�3�/-��Tk�Rg0,�І�Jk�� t�õ����X��Q|����?���O�d�Ъɜ_�Z���r
ɹ&��^���g �����K?����4�4��_Y�绯���1
x�t���`��䀠�X{ol<�4��Q2$�D���h*@>I�Sq�f�_D�l3).@�E�M���t����(˺(A��]��u����F"�!7Qm(2�Ѹ���~zf'T�@�����e�q�vr6d��dp'�|���RW����Ms$���!G��� ������;�FC5R֖�L}Վx����5Oc^u9�>΍qꃏ�������Ypf�_������w��M9�^{� ?��/�����g����U��!�̢|��<���&U
Nڨ�����]�y��l^ڐ����r��|��w���K����Qr�?�_~�7M^5
��� ����䋯���?��ݾy�Ůϟ<�_�������in�ө����A
6<3�Y����t����c�̏ev|$%��Pl8C��GИ����d
\g?�k4�`��!n\�,��{�l�.��"�����k�=9�ѧa��^��J'�v�C1h�6�A~��)?9�ݧ!.��L�fkm5�i
�M�N��Ɂ��$�
:V�����荛r٨wx���6x�F�)n,	^��Y�SV��'(>m%�sym�JD�I���iflm��l�$=���z�H��y�c2L�"XN���xL򲮍J���V��Q���Pi^m�܎�1�OS�Z����.juAb0�"z�̦[@��t��Φl���Y
D���PI������!G�t�~�M��8���_t�5��O2"�E��9�sk!d���$�����L=�/�*ԕ�EȋI�?k}�s����F�)�Ә�(0Ӵ��fJ�@�G��u�37� �LjF�_�|\�b:A��D�uM�bE�V@T�L�_��1��M��@J�餹R�vZ#!͵�/_�5�.�TA\�̏�H���5�s�,�`<10`}@U5\g��E�'gG����k+}>����u�N�Dv:�S}���f5��4�,��9�x:7�{롚�y{���e;B�@!�s,�?<`��f�_�Z3AP�;M�
;�j�� @G���	.R�����l��"��p���	�X�^�ǰOC������ۍ��^)[
��x笾�naA�ΒS�PnZϪE)m�YE��?w� ��H�`.�j�n�zn1�T��k����̝v��\F�j��RҾ^/҂�)�:J�3���t6��﯃�. �ҏMQn���#[P��!��a[(E/��4:�)�7ot�gs�M���e�D#��b�Z�pp��9�C�6�M�)#��ᐱh��H�,bA�'�Ty�ٚkD�	#g:�t"�a��I5�L
T��^�;=$a#��V�0��t:zQ	�c�k+;��a�c��8zZ1��=J誚DkS,��I#A�E;z(]�}G�\�&k���g#�V��҇@��?���D�x��8+��u�߬�A��U�C���# ���T]�������{mOF��j8r7]#���B8��V�ב�1��/9������Ƽg#b}=Px6A@�*�>Q�"�'����>��:L8&ݠ�v����r�t��U=���B��S
,a3E)��N��8����j"L�5��a^6����Q��h���׶�?�V��D�Vl,g�"���j.J6/�%x�0T��b�C���m��Gˏ���r��ӊ���wSnݽ'��O�D���@�Ͽ�y��m�ve��u�tu[���;���0�]�d$���/�W���tƵYP���~!Ʌ�f3�x8y������y���|"/�?���-��a��OW�|0��jЯt���H-m��޽/w�{��֞��q�� Y���&�3��f0#H�Q/������
[�9>9��v�֭6(�ITf��&hp��
��@ ���Cz˴�edhlu�-���{>_��^ެMc��^����#k0K�v���ӹ�P�99S� �ڢ�0k�K��49�G{�Z`g=ͫ�ѱ�NFT<Q�R٧��\�N�m���87��p����ij�a}˷�6b.����J_�[�A�bȧ��7�%�]+�AǺ�
lw����i�_�\(2�y�fz��heEl�*��ߊ�Bk ^��v4����� � 
`O��<�Z�X��)������wqm&��K��!��j���ע��l_߅�j��EL'F��W��9i��ə��<�6�`�A�[6-��}��E��ϼ���;Ժ=����]�]V�>�]����ݗ K��W��*�XS�ŐA���[����*m���^ �cH4� ��u
\0� @�ú��D-���,QYX��׸:����6���`�eɦ�����؛�6H��+;���Jlı��%��*��Pv���km��2��|z���7�έ�p�:=O��l�V'�
�5�_��M�{.��צ��x�A��S���K�\��k�2\�T�q4
s���4XnԶ�Jh���}�ЮI��'dQ�^�� `Р�c`�����V����,�Yk�E���4��_w�;�.N[���r*A�!�֭M�h&Gǆ�����"h��"�hu��b��xb�!��[�Wdd#�^N]`BB����+����B�{��ņ��OQvm5E�i���Vd��k�TG�ä&����P�$*D�
c�y>P��e��#"B� ����}ǔݰ�e'58�����@#�N���jrj���>/S�@T)=Wh�!w����k�`���f�M
��x>�����~^i-�� M�����.J۴�@T��r�m��{��8n����:��]Ғ�*_�N>���$�QW�4^ ���Ixup �����'�R@3�E+��"�NYX�R�]6h��JOu��S(�q��u�� K[���X�=ї�6x%�۵��Kl��~����_9���_$/��zX�J�dԈ'1�U���r��:�(A����Koe(<�P�&|u�����7�ɳ����z�+���@��'?�{��ɕO������EO���g�u����4��X��H���Ѯ�L)0(^%]�T:���I�G��������-�n�	r�<�&J%T��fքLࠞs)��Qaj)~W��=�Y�,aC���fu\Kj唯⇺|�b���p����ғp�akz]�bƹv���n���SQp�#�4�����1OQG��/�AN|�^F|pM��a�i�{7R���pM�5p��=NA�����G�Q]�����������"��*�؂�]K���,g��<vIÂ�Om�F:�3UJ�a�j�"Ք�+<S��E����+n�FD�o�ͩr�FγB�1M��3���T����h'p�_�y-���v�#�HU&g�����4Ku6K(���\g6���}E�v4�[b
���.���3M�����5N����顜,���̚����qa9�I��2�� ���<�6�Q�X�&���֪�"��)#�׹W�DтJ]U�o��=dy�jQ�ܲ�A��i��lT�4wz>+�m�)��4�H�`��=�Jp�k+�-�4�@?��N?@�QaE� %1^GgG�"n�[td�����>뮷�N��޺߄����(�ᴢ���)��Q���w�����2f�}����lR��jKG���,�yQ�՜�e�����_���ύ\w�t����YFՓ&��8n�f���r�с�td��#;:')�
|����"z�����	�*T!����A1vIS�G�hw��6���Dn\�,��ܐ��̾x��<]l�PZs�|qP)�>���D����ɏ����+�1���Lyw�Nqg%�JX�[���Db�0��$ʴ#�M3бg��C��wjCG�ȡV4ho�@~��O�	T<�u���;>�4���ݒU�=D]��D��ģ�ũ"�J��t)Vhe��]���3����R�=�h�]�j	�$�I-�^b��1��y"Dؿ{�D?}EN!�f���	�27V�t�RP��R���W������h�C�}u}#_g�㛿6����^T6b9��m�S��64�	J��pc4��A�uʹ9؍�c�����d%� y�x/,ty3»nϙ��2��==�PgH���;F��z��ܠN<�����o~-���.��GLu��[Yې�K[|߷�~+���_����x,7n�aa�`u�����ã}��>Pft��5N1mhИG��MX:r�6-mD�}l��ɽ��y�{�) O�z_V���@��7$W�;��yR�����^��P�i5]�q�<�[���ϟ��3r�4��
��q�?��y���<�z�m��ٴ ���k�6�����mʌe�C�e��
��pj��68�i��,����Y8A��zց;pp�]fu�PT~	�΀�<�Git��^(��hx������_�סm���Z:�E?Я����4��	B��S �V�:�@�u�������:'��hL;>d'lm����P��M:%��3�ٴ��\d/���C�^]:�w�]Ht7�?���U���0����1g�6Y@f���Ը>�����`�6˪[���v���f���]R�M�j�;*����>��'�n�(�Q�I�8����Cƌ�S:���!3H���M-r��捻��Z�����v�k�g�W
���(-�!HԅbMo��J)��	;PՁ����`7�jT~�G�83�_Z�-o�*V�d�U>жLS�A �:��,�A``�%=�Ǐ�oƷ�~�����$�}���xa�Zj��G�	,�/��=�-jƐ�v���e'|ym�m�9��7�]~��k��U;����i����[κHK��-������m���4��/�n;_�yT>O_����n΋�Ot�i�k�&��ZW!��6�@��3>õ�My'm�X h�����y"�N\jO�>u��Uu >�'�?�Zn^�N����_���3:�Q��f�"�V1��-�W�����S00;I�9���&7��

#�t������j`C꠨JG2���H<���j��`0�*����e`��(w�8Ӏ����
a���B��6O�	�d�Z
pG��lґ&����)V;�U1�oB�ZQ��&�SiD�]H�ԋ�2m��t�E���WI
J4U�b�N�d�3;����<PaO�fl��s�y&�3�w4��*ص�q )op$je^��}[��F8��k���5�	�x���ah��ˊ�X�,J5-y���"VG ڡ}�ɽ�8�ǿ}x*N,��i�S
�}D�X�P�.щ �-"����([�X�=!�{��$.on*�#m��;W��(�o�#wn��s���{֙�b�i2q���y�:5i?:=����ɩ����J�&��1]K7y�k��A����;����۲p �}��\����(}�ֿ��JT2埮�48N{{2��皂� >�j��^)�}���\3Z�a���	]���Z�j�,�Zr
�V6��zmF����|͊q���'e����-4�ō��u.T_�"���jQq]tw��4�<<� ���!�~^� �����y�kO�ЬjMz��h����ԏ��Ӂ�9y���x*����le,����[/�N���Է���A�qC�fTs/* ��@�i!�j�=���0�C���<u�j%������ʮР����T�2�lՊ��́G}�σ�f7h�3�4��4�i;�<ʢ5'�;�M{�J.���	E�R3pE4��Z);4 '=���{d\�hc>�(���3hn�.�n/�"�c�H$_3�&w�k����ڰ�lv�ˠ
gF���]aK:���:���5Tg:z��ᐁќ��ڀ*�c4�� �m���e���� °�#p@$����@iz��Ri�sِ��P�y"#"�Z���^e��9�l����峛^8t�b���X\%�"����}�u�/
le_�/OX�Y���?�kׯ����<{��N�^Z��i
B�]���v��'+�}�l��u����TϦ��ŵ�25-g�"��Z?ǘ������\�Yk�������ZqNUwyO��y�?�����7ܓg=�����A==_���/�^�kEX\�
���h�^���M;e����F~lߧ�	A���(<��ߍ��ú�6Pt�C�Υ��K� '�`���NxD�L��D��6��&���K��i�ޒwn]���w���'�zz�|�H4�)�޵S
M;������or�'�{ric���oݺ!�w�LF��Zӕ8���"�MUn�t�ŚQYv\%���'j*��j#J�-�acC2���F��mNL!���}�&�HvD�o�^gA��uo�_Zd�M�]�e�|�py=�ܪ5������L�im8�#��(��SG;��Qr-P0�!4�@��rV9��&TxM���r��ӿ���+"d]�jy�(��ق1L���%���.�Q�m��h�j�P�̜���m��3�t䬠�2V�s��t���s�V�`N��؇�o��?�5�qN1�a4��
�X3�K:̕����[F�4���A1�RH�T�ش���89�hȅ��[�nɍ+W���gp�W�t|��n�o�Q�����=����ӉBP���g�e��ݗ����"Rz�ʦ����M�3ONT��v_�_��� 9Ɠm�Ay*9��q�CO�/����L��G&��p|����7���'<�X����M���J'9���>U���cX�y6FR�]�$��Ԛ�P�
�?֢2m����˙�	ք�YK��Պ�/�ujͳ�6��b��7�Y�ؙ0����&�A� āf5m����uB�7d_^���� ]�0Р�V~�ˣ�kY���߿�ڝ��A 7��[��m��[?��=�F�*�U'�1P�d!*9h�XI��u���d��6�bp����u�);K�,̦���s����.���)��k�|����I��;��ym��2s�����.��Af({�f�,��Z!�A���(��ep
�@x�1_#34�^�,.�湙mI�\��1����|hJ����|�n�G5���f�pıO�5���b��	T���+��+�L�8?�f�J�]�i��v�<؉q:�hRɵ�����@�G���3�B
>��gT�x��yԛ�Ok��XH���y�+S#�u
���xlm��rp�'W�]��?��>�P�޹���2�) *n\��A�E�{���T]� �4��u[��XY �Z���܋�e�}ى� �
6�˜>&T�"u��!�����1;���:ƥ�X�ܢ���p�x?a������1��g'z�k��5�x>�a�Gj�,���ۮ�|H�Y:Q��Dj29V]�sA�hmHE́��h�==����߾.er�OӤ��+A��/pW�Y�&�?M�8�g���*MH8P�{��rX��t4%�j��P�N�C�]��J�ʤ�J��ɵ�y����dܑ/��ViaBVJ��)��-R�#�����p$}/�צ�㈔g�'Za �@�Q+ǫ���|C�u�v,�ț�"��Qd�k��wn�n�X��e�ƈ����ę��\4��g�*~�о(
C��tچ�[n���;	����7NCٱ&#�� g�
���ա3_�=k�a�c(4�4�&^ױ�?�J/Qw��P���@���C�a��^�R�U�1(���vbD��ֵ֊�m��q��}�{�aW�ߛ� 6�����V�ѩ;9�1T�H�d��WlvP��xwڅM�uB���/���H3R]k��=Ө�#�����˟����Nr�;@�J-�-g��2j�9�3�g�C���&�f��cs֩�n+tŜ��j
��޽/[���Ƥ`��}�q����%x���|��a���Sp=�ޚ�׷�Sї��8٩�����`^�&'�����
!�ʃ��	\�ʔz|��ׯ9�Va��n!�:�������oz�kN<6[:���}�r���g �/�J�ωF�s��r�Fk�*�zن�>_VM1'���v�$hV��Թ]� LFg�wt"/wO�@�^ ^*���������@h��C�c�T�X�$��B��-� �>��h�M(��$�s���>�28Ǡ���s�2�(/�+���8��ϠZ�܇Z�4��zƃ�j�p���^��Y���@�YD�G��Ӭ�u΀��Vqg���*�;������
���4�43�8���u�<�~8k$"�B�0
���yU��� #�L���03;O�0��X�/Թ� �=��ECM�=*�}��b���{To����*_�I'��{�{ɟ���R��ɓ�1�%�=})��m`��8�!�v� �Ke=�X���w�Vm�����̋QDtN#�f� ]�F9����z����̘����Ɠf1ᬟ��������:�n����̮�-�Om�n�@�%�9��k�"�=�����K��o���?uP>�hm
G�m���u�j�ѫc�ʥ�����J��C��h �Bn�$����_���#���#��ߩ��B{�7uU�i����o�&-�����]�fH?�N��uB٣UC.�޹!?���l�AE�BϹ�[!m���d$� ��Z^�h�ڵ��{�e#9}w��N�-9 �5:әJ�t�(�k�d/��������Ε��u���������[�{x$��XQ�w�Y3"�Y���<��D2EʹYW�Zy�Zt�FlJޜ�/�q�܊��Ȩ�=W�<��A�,���0���Eti��4�@���M�w���t}��,Tnآѽ=��Ī��r�Ƣ��iג��jK�1T�i��M+�7���q��Tk�5Fc��������&�L%�h��E)�q�Y�2�Euܼ�����|��'���|��]��J�)E��Ô�刦�ISٚ�t���K�;.��MǠ���%�\�1]�����Ed ,����FS��躽gn��#OҢV�C
ym����W��<��l���K���$������[���۷�N���Ƭj�1�m�9�Τ��}��[D����W����Uy��a�/+D�����l���0Lk��~MզTm�i
�6euc[�>��餖��)�x�D��si�n�������ȟ�[[�:<�p�Њ tg�wa��=��7�hӐ�`lQ:�n�N!��>)q��z�=3|N���^�<��TΑ9�9˧E+�����s>���xz3G��9����?����iܢ�v_��ёU�0��:�t|��_��e�Ε}-�]����.Xmߔ��۬Iu����`���K�����ka3�؂g���Կ0�Q%����Ki�m�j�����M��A�Z�d� Tm0�F'��ٌ리)@4#�=צ�,:V�9V������0�;�n(+�㘠���3)LYY�ᚵh\s(�8bԙY��=�~��3g~���t���N��;B�����Ӽ��U�S��hB��'����F^�Zؤ;G�S`#Ag�o�:r��R��Z��a�8 ���^��M*Ki�-B?��LP�4���9͵@@|� �#�����X�#6�uH!��� �!d�/_ڔ�W��F�-��_�]=y"ǧg����/YWP���J+5e�C��Yh�$�3�L�n�`m}�k���?�J~����<}��l�4ۗo˓G��|�L�O8/a���5u4��,��+լ�qPd�{@��;����㏢����r�A͟�ڴ,sZ7 #זS^��'��2��(ZJ{����A��Nk���A�sܜ�-G�����ϭ�`L�4���n��;�i�&v�Cn^ۖ�|���zr����}��lj�e(l�L؉����\��R�}K�!�G����
e��GGr���bTp�����o@_�Ք��^r�3�D��P��������~�\Q�����a�p� ���~�6��	��:u�)9�(�5%�N)�Fг"Xl0����ͼ.4�_Y� ����E��>0PDȣM?���Vĭ�T���tza 4����C��
�����X�Qq�1���c,@�F��'z�HLu�'�"NDSJ��u�6k\M�
U��z>�4VȥՉ�	���8=+|a���(-;�����=F��ih
��X����*=���ׯ�8͍�_��O����JdE����\xPi���Xq��t`T!��-�gS3�ċc�D��^��X��/��E��|q��<�wFa:Ay̞]�F��"f�Ee5<��c<���`C>i�۷o3;Ӻx��X����y������^
���<��9Ik����Zd��4״�I�!���gO��~rt@�Y_�Vr�х��dk��R�Jȧ�u���M�@�d�ä�3@�Z�N�5[�c�����ƺ\�u�2[��+wyQn�������i_�fx��kմzg�ւ������Fu�n:&7��"�Bu�ڂ�#)G�V`�S#ʬI�r�u�gy��XkG@r�Mł1Alc�i���\_��:{x ��?����HlV�h!��Óј]��>u�Q�<_��+�p	zq�k�_��B�<Q��*�]����g׾'�[�4��?�I���rmF��L{�ͫ�J��*�ª�c�=�\i+��>VO��(
�E�60;��B�ϊ��h(�`ς�j_�$v	h8�œ����GI�=��e���L!Ҳ�fd������]���
:��̅����t�`瓘�Iֲ�,���룸� M���f_ؘ)m�6R=xv
�sU��ݚ�8�	����Je8M��	�/�o ;Rk�/����+��ek[�Q�x����# 	�v<_f9�3���L~�!��E��s��g1L����ﱣ�o���������m0G~p2b]�ܸ�9�M%G�~��czVD�k��0@{�{�|��C���)��ٹrY���(�s99�WetzHz1��B�+ u@��b�ǜϷ�F���)kJ��7������j�/��m�3"KhvS�����G��A�������P����ͷ�>�۸NK�[4�P~	}$���ua�lT�2��)0����^^�-�Eއ���$پ���U��"da���yEQTe��U����U���ɐ�î*��*O�%m��~��|����>�M�V��ㄅ-uv�0��V��7]OhC����:�a����wԓS(�L�=ͩL�h[݈B�4чɰ 5ʀ ȹHFQ�ɠ@�.c wZS�Ч�� ��+�CTE7�9x�4�K.C�Ho`D�"���=��-�k�5�I0�	���᪬�;���V�㺰�kK��P�o�e!��2b��uϤ�ȫ�뎥N,3�&kYGw$�B�F��A�$IJZ9�%�	&8")JuE�%"ǭ�xg�ʚt��2�68|Ƈ~(����,׸�t������y�t����t����Z�Bt -�Iƨf�D�I��?P�q�Q�HVO�����G�Q�S��������k�+��O*#����2x�i<��9/��7����r3m*���q~��}:%O�?���=���tL̨aL!�z��/���Fs����y6����I��œWЉ((㇍P7@43��9QJlvx^��9:>&�Gax���'�:���yڙ)y4i��,.��� ٝvM�5��%
!�U�i�a�'��D�b<XΩSQ�?h�6`R��-����(<���Dny�1��8`S�C���yxp0˴v+J�N����T��$��������󰋪����:mck�=���.�GO#�kCݚߵ1^�f��I�y�z��8EC�z!o�ÞvZ�����ŕ������G���
�˼Ɋ�8�}p~X���[Zl �7o:�{9��D�a����q�3���:j�t�h4F�/`�B�0|>��cE��ll�֐�3����e�(l�ɦ�����G�{vYrׂ��򦽃!#� H���ӗ�Z�f�_�e(i�@��m�������̜�wDd�̺�0��X��&�9qvD�ر����?`��q�χ2�ՁC悟��=+��� D4B^�S�P*S���0Ј拖s�멪��UV�'z���Fe� k�w3F�V�2F�	���	c����~��1�D�X]w� ůy_�fdpR�Կz���}������{*�u"J�(�dK�HO�A�l�ma �p�Ν[쥳��1;<��|#����T��x�7�_H=����+p��͂��B3������y[�e"������v*n�&��c��d]��wf=Y�֣�`�j��Ѹ&�Q�w0��cxFJi�y�/�)��6f�����}d־�;�V�Ϲ��Zt߃&��
i:���3
"9�  ��Ӣ?�a�$�ˬ
&n6����j��2=;�/?�X����E��{R�&McT��[8�/�ȭ���J$��^����v<c_��Di�Ȥ�Z�a�L�^J�ڠx7ce��p�g.��;a�d,���B�4���[iӀ'�O��n|Ue�f��{4�uY��2�v |��*&3V����*8���E7mb���z�xn.
�M��\TM�� ��� ��)�x�IR{���T�np��5���~��CQ[v��4rS_��|�N&wx=�{��bS�/��O�"�0��{Yv.���W��`uE�/_��JV�&��y��9�h<k�t)�Ǌ�n�C�4~9b}G�S���60Ij�n��>I-}zn�W���}V�7��ekO�(��-�ǹ�{$�1��%*�=�?~��$LĝK�d��(ܖ��5��'���3�{�\>8�=����k��ޖ��������駟�'�q �Hs��W�&�al�q�����U�{��6�(�����_%�qiq�F3����h�³��0�$ �G�<$ow<�ȥ�7dsk��л��,�!W� @}���`����(�M8�&����>���"HE[D�Բn��3z�	Q���ӘTqE���ڕ�#l������0GO�p�&�����^���J�j��FG��@��J�q܌b~�˼��]�66!v�Z�������)��.UC��o��U՚IN�Ds,yb�%ةŤ����l���\*���|f�:#�F���G��TH��`�l8v��L�Y�2���y�3��@Vp�z�^z�agÚ*[�_t���b�_�~qm��^Y�1����tVv]>&c�YՁ���p�ku3P�]�D��Z&�.r�S�Z6DUU�;nQ;(*�#����~s��I4���5��=k�� <u\hL�J/�G�kv�2�z��Fs^*����uj�l�QM��TJz�a��e=�{!��}E�0  ����v|���j4R�4���ϑ���y��u�I��ln��3�|$�j�[����d���4�'2
�8� �L�B}u�e �ee.p��=�G�)RY�у8�;��X�0��������y}�Y_���j48�{}��:�6Ih�1�]�?(ޥڝT�>�:4��g���^���̀��Z�>wbձ�֬0)^��R����#V�]�1�C U,���bkv���	]��٢��`S��G����!�n|
�h� �ۥJ��aD���+�R&J=�Q�>�I�E��Je�Ȏ��г;��� |��čO��a8θ�&	��P�O��)��&��i�^�k�F�atR�9��������k �+Kc�J ��u��!���ra\>@���k`��2U5�:
n�����~p�Qlf8M�_���nh�(����뫽s#&V�g�д��D���wh�/1]�p���#��q��.�V�B"��G��B�(hR����?�mhz�2���|�=JNV�!�0�&�H������	��ʠ�A<�q ����f+.�X���,�&ˍ[w���͋�����fV����}�{y� �W����6�����������g��ûw嫷ސ��[�����7�|C����h,*�ME�YAË��`�\󙂚q���w_�@��$}���*W��kF��x��F\}�f2���B�lp�U^��_Q�����J-m��">�zYCv]D�#@�f�n���e��Jkl W C��`=���Ô���_j#��e�s�M��S-U�HV������Qֲd�Sp�lB��/GG��2b�l(C'��8t�
;w�8'�̶��d<3��ξ5�I��X<n�Tg{,��Z��Ѻ���W=�����D��<k,[�u]' �9>e����kA6��Nt�4���SR��N�oƱ�B��|o�9�u �8�.��@�x�3%݅��.W�>N��!��,�=��{fD��J�p�)�\�&s���פ)dM(�g��̮G�{i}|������{�h�u阞��GJ	(iQ-��?\���n�i]�
iH�y� -��f�8 �5�6zo4И�>{T����p���Uy������7{{���a�T7��	Us
ˎ��s�h��2פڐ�c8Zc�*���G�&k�#RQt�iD�9�B��+2el={�'�j*�.]�|X�R�x3�W^TR�o�g������d���ϒ�n�3��XfU�Fs���n3�x�֙׊��Gc"и�[3��h��20����-��AĽ�>�wm�)<Q-^c۬�:qۡ'�YUZSK���=��}w�eX׊���jU�`\�{=��`�����{r���<���<��^X�5����n�t2�(rYG/�/�;M'u��E�sUH���F�+�1�|=x�k�|�y �gP��A�6U0*��VT�Qni�P ���0@
+8C@��Ry�D��v���=8ˤ����SM�V�S4�������au6�2(�u�q�n�I°�@4+���}������ҵy0���2�\-C�U)�2��4�I;Iq~d��X�^d֌����;e�� 0�����	x<
��"�gd3K�::�5�y�}��'~(�v�	�a�}Rk�%+
�_hca�V�ٺJ�JVz�F�Q-dr\*l���FaY���L��ۭ�fT��n"ޭg_O�6ŭ�j�wڒ:�d�"�b�o��eꄄ�xq"�'�J��=Y�� n��3�i�*�`.�O��?}!_��=��CK�4�	���̩��ڗ��z厼���ȹ���C�noo�"�������H%#=��S�S�����{�j-�e��r|t��?;����p�C�DY�Z���V���k�/+a1�!j0f�PCiܣ����ȥ����x�2����t<Vv��'��Nl�/��)1��|�Hu���N`&�%�񴹶.'��\(A�¼�u異߫���ȋ�}���K�ݸ!(���W�_���'���&�X��%�㱬�"���,UR���.(�gTD#��'�x����6�A�����[n� ��!�Y4�z4p��,,�X���e���YP �yVG���6�hX�������+R�m�x�/�D�)�~��Vg\��#�.ݠ1��6�C��pM6�E��cs�G�S��	�#�0xv�|h�hr��wꦴ����RS��0sc�����XK�G��Q'�oE�X�� �hM��̋t��>o�0��Bf�<��N�H\.
� '�_\W� %�N�5?~�|��=9:����<����J�W;��;�)x��5��uA5"��"؁�鋽���p�(��� �W.]&���O��f�� ީ*��K)��y�������3�ߔ���& ]�rY~���l���+�;&UR��h��fҜ�Ć0{��Rc
&�K��:�D��'�;�+	As66J뿑��@�;G�ҁa��Q||��"S
�g�'���H6tA+Z�D{Uj �-.R�氁xU����" �4I�<�J���pN����#�.�F}9>���@�i�b����(��Q� o�'�#b�&R��QO��Z�� �*�3�n�)E�Qz�!2\j4��D�V ;���\#}i�]`�y��k�U;��UGF)���~�q�C��b�Ĩ5Jiw\@�D!Ń��$�����֍��
��
�,m��9M%jL=9G}16@_ya�<�=7�ۤ$�qB�@� @��a���Q���(�
�I�i��v�K��[���+���ó8Ϣ�:B�@]B�i1� ��b%x��A�g��F��E��]�༼��c�ݫ���ꄑ�`��^֨� U�RO}�-��V4V�K�Wm�/��ɷ}/�dŭ�ۜFK�z�����P�?��@�$��j�F8V�6i����#e���0���D$����������c6��S��mk{W3 x^Y/�_���XS��Ɯ�����XѨ(O�bi���3�@��J9`��ƽ OkwG67�ih�&Tz�E�lY/��``P��X ��<y\5�[(!M�@E)\���E��19�^XL �x4��<;QkJM��	BK�k�u�
:D�,���^K�M��{mj�S���`��b�cG��k���#��7�j6��?�b��;8�?����M��l>Oke�%[*^��o�߫M\���2��ntJ����I��L!e:	 �bL�G �(is�BK�p���)XyD���=��N�?�~��Rd�b�ElE�}�'k�w�"*���wi�L��lE��ι�h7N�v��LZ� ��~���Al��$y����<����躈��&�N��;?w��Dfc��;o����uBF��S�5������ʋ��w��q�*(d��Np�/_ڑ�����,��8q�i���3T�=�~#^��d" ���}��%"Ú�+jq�ss����tJ{�b������v�( w�t�GO6���RKp^�������D������zw�J�^��fe	v�g���n߼%�(�{��g��=
׈{���QDҩPfc�)�1 �qm�y�& W�45��SϦD��ƪ��� �u�:��5a�����:�s��\ӎ�C�9E9�ճ�xᎼ����B �_�]]�pU �0����9-�&�|<��h!��R�%MM�/\8tdS�U��ri)]�@�%UA�0�5b j�P$���h��C��%��b�E�TӃ[(����Fa�fV�*���F���.,R�\�E�3�g-�h^ yS����M��5�ElѮ����5S����<PT�P�mT&�E`[����5�(/i;r�t�+�K�j�h&!5pL���l�Ԝ!���뽅zh���{M|�aN���q1�r��"�)X�2f�Y��(��=�NX86���U� ؕy���Z$�-i�&�#����P�6��1�e�*+,�/��>�$���K[F�V��3���s��.��O��_b�ΨY݌�B���^턙x�Wf�g�{��` w��ln��9y�k� ��΍��CqrQL8��'�l�]w�|��x.����&O�y��\~��ɛo�Hn޾C����Sy��P�~�HΎ�����p �0��W���� �7/_���)#.sk2���v��|�\�q3,�W�|q�¢zU�/A�Y��}�`l�GZ5�Ok>�ܢ��-EGV�5*ӷ�H2��|�������dK5⧎6����-}ܖ兩��&Q�&iL������(�x>�Հ1� �/����W��U���EmO߀*�k��$��k<�G]Aq�>�5����)8�8�4E��yM�|�w���j3<2
@���� �y�ݶ�]�tV@�o��jϮ�ާj'������YjY��]>J-���.�Z4
O���dnT�:C4o9
 :��b`� ���ܟG�D�I���GM����U�XT2i�ߥ��V;i�zoH�6�u� c��\aO�;7b�H��� q}i�Q\�����/�����ر�7(�$R;ސ͝#<M�:�	0suQ�8���E��7�+��V��<�-l�S
2mt󱶮���Ɂ�é=�ojD�`����]�sUn�y�$t�F��O�Dp�ɣ�|Z~��������Q7(��M��sFY!2��+�������W���~�S98<$8�]e�������׉&�_��<z�H�r@���j{>�{u1+�EQ�;�zn0��:w:�΀x��X��I�lR��)��^g�����h�,��+�l6x)8�p��ș�NE�~ ���V��l
���A�ONe6E����H��J�"I�_�Ŋ͗� �f{��nũ�r;t@�U�1Ҫ�jM��/ΊRh4`,�5��*
\��<ri �+U��+�����9O�<��SZ�L�>�<�T9�^��c���	ӨY�F��iƶ��gW����2�����: L~-�ĳ%x��MP�gEv�%R�����L�c�#H�,(�=�zvЫ�ں�@��٘� Q8�F?�L�&a��lz��6 �3 ',������#�f�P��6� �ǵ����Ex-l�)z�0$VHdE,����kL�C�v�HUV��O,1`qzq����j6-ioq^��$��<�Os�1�;��3��ꚜ@���"e$3믆��+D���PN&Od��(�=�LQ#_0�>��`�O�I�jdO��پ�@"������A6�������7e=|E�ۻW���ӏ?�'���7e�ceI4�A��2k�]�uKnGq\���(>�v�ܢ���掬�n��C�Ѐ�^I$��4��3�|Y�����dm}�ꓳ�;�ex(r
esq����Hm�'p&!}�����$��U:2�n�p Xk9�*c�q�%Y��Γ6�*��Iw�t0���@pDm�[���4c�l*�2h��V�F���b� spc{�Q�!�7gsv�T0�Q_,X�e�MM��R�2�]���ݫlW�wPc��c���`�X� �\j���ܖ�~����Y��ʂ���ؔ~�`����j�N�	��Q�#����l�M�{�����g	X2����}�����w
6f�c�`]D�ƣ�*&�.^�����R�2ĝ>� ���"��hS�h�q_��76̣�^��@K�z�6��86����0SZ�9�X��Aqݩ<
<o��Q�B�cQ�3��in�����_�Q� ��fZ<��}��$ꄪInN��vga^j�����S9+ ���P�n#ˈn�8���M�v�
�*"��.��+�*99�-�x�R����]�_�9φP��I��ϨT�%��pi ���;���B���A��>嵾�ګ��oȣǏ	�q@�(h���3U<6�Ǎ;��ØӎH��l`K�9�P�j�B[�ʷ&�9��٩,�{t����l��õ��q��}{�]�L�}j����iU&?���,	�O�fY�!�Od���qP��jx�=&��o��T�v��-hЩU�L�v^#Ж��+�lZQV���9�Ra�f�� r&�$�Pm���6���l�H���ϐ�Nv�eS�9'��EU?P��yp�nU�RoJ{�Y�w�Y��r��P�*˔�⃣��+���Z�TV�\Y�U�Pؽ#(Ϛɯ�_<�V�͠�<���-K����mV�Xqje�V��R��WU� A;�x�b*>� �a.�lH�z����U�~4ݬhJp
���=/Uz��d4��px��ɔQ�)��l��[9n ")�Pݢ@��d�b�IRG=1�:��xaaR�ikڂINVjĖuZ���
���Hw �N�����ǖs�}?i��Cb��ީη��5�B�	ҩY����
$	�js6Iu��l0bqi����k4�}���
�4PJ���T�x�O� !�ț��)�7�CVz*5
����|����x�M�{����������H�6w!�W*��d �t|���D��S���G�Up���fEƳLΞ��x�!�;/��eggW.]�I��'�lB7�!:��6�AM��rŋ��79eq'�0����R�J�������k����u��W�0�9���1z�]��}��ٙֆ�6���u���E��2WP�����b�9U������p�[Q�����*��ت�H#�D��}]
�V��xu}E^�+��p�Hx��{Jg����.�$� `2�Q�_ZӲP��\A"�4��(u>�ؕ&��jb=6�ks������{E���Vi�Ku�����G���;�j��wϙ�L
�da��Y=A��R�iS���mm��>� �R�REӴ���1�QR̵��#�vh����X4�A��蚦�>� �h��-��bbry(�%m��걂�#� ��
��Q�����5��������rWUJ��ˎ��
5Y۲ȡl$VǠ΁�G��P�� 2\�'������G����H�;C����T��ߝ-��`YwRĵ� 
%��"�
%#�{�š���)�j�55��3��u� ���4�;�oʓp~�G���P^�}G�/��措� �>~��� d17[���g��Sp�+R��`lt^�sMlSw�N[����Q��+�q_I�ϗ�K|�q8��;�:��Fӆϭ� =���:�g�.1�����E��XY���-y�WU.�kJ��EЋ����0��c��={�c��3�����`Ȩ9��?/T`�YZQ��W�+B�V��/Ue$��督�a��i<ӱ�b��p�5�}��"�4p�i��,M�����d��}B�|V�iM�Ђ��
>�y�ȣM�,
I���.�r����m�� ��3(�`�捨�W����x��[ʦ.R)��/�6��Fԓ�w�dƳְ�DJ������@� �4ky�g�RD� ���)`��RZ�_��kM�¢��dq���5�j�E�|��V��	�^��]�o�8��u��VvSݡ��� ������cQ�}4�r��`أ�#iJaw��''�h�
���� �Fm��u���N�CTG�3)e��)$�)AX�P�8(Pn�G.��]O{t���P_�2��(��ٜ&����.r�ِ��܌QvD=V��36��*2^C�H��*��-&g� �o	�: �p����Q�y�F��|4M@�)It˄�;z�/��Ͽ�����J��ڏ���V�����g��{��t*��=_����a-8�h>3D㢕U9y�������b2d=�`�N���û^�+���%J�X�Z�{�:Z3��1�o��Ր*X��*O;�0�3Z�s�����S�ʧ��W�\#���
��sΗF���Q� M�*E`c-�k��FȆ��H����Z��pr�],V�h#"D1g���#O��!��9��;����,��e�ΏGl5��j�UQ�!�`,%�~��j��+ !D����Uk�p/�5
'�w ���G�mU�Fq���1�<Ť}�����͌��*1���E�q'�,��1v*<����@5>��;U����MƱ{^�ke���:�}���1�+�t�FUI����'��9�8��r��ܗ�MѺ�6�s.�R*��Aa+��_7���r�XJ�kK�zq:���n�Wsu�*��Ͽb�������l����I	<�9�ml��x��6�c��E1!�O�S�-�%�7�Rw̾������6ς'��n�Yo-��r�?WE�g�kF�m�#�G�v	�͕+W��	�%e��e����GQ}��D���!#ㇴÙQ#}��3��f�9�5$*�g�5
&�?#��<θ��	k�{s:pH�]����z^(�����ɬ(6~X+8�D�ԐF��V�Sn�@T<3Кh�Qi�Z�����"Q	&��4|��@���4�i���YȨ(QY��xt"rq+�84��(kDr-�o���T]��`�-�#�;b�(2�*=���a�ui���N�	T�9(�m|�R)���L,z"�.��ɟ�8���m�⭻xņ26��/ٍ��#Y1�~LF*J"����=ַT����r��&��P�:|���}Nrވ{���{�t ��u�I��8%��<��^f�R[v.�S5h�<jRY���9ŕ�A�Т����8Z�>���u����v��L)N� g�<E<_! ��=��U˝�y�o�{}m�E)���Ʀ��2/���7��8��cf=M����l8�� ��οU��������F>��9:=a����$m�B���_�i �Ϟ��I-ǝC_f�VC�OWI#�L���)id�o�-��_AQ�E�T��<��g�2M��4�^fI�l�/@�'���F6ibR}�b
1�0WNOe��v ���Y��H��Dq2�5��q���;��KW6�Z���o ���6@�ؼ�(���|ݹ�O㌔s�!�[6����i�S#�֐�0� �Kv-�#�A	�Z��ش��ү�ld�`;���y��RR���ж�M�e��o����Q������k�wv%4� ;~ͯ)����(ڎ����{/�4��\��8NZ|zY���|4Ke$���mwH�a���%qR��+m�[��<:8�� N����_����g�{�uԋ$�� <��\F�����U�snMɊ������~6�gdY�N�M������;���d��,Y�O�u�(�O���|�LH� ��Ukv6��>|��������� E�ޢ�6t�eǩ6FCA��w��>�$0 }>��3լ�{��"p4������Rب/���c�����ҹP�pK�$|�p}��.��p{y>)���\q���X_��=��2@uq�z/�ב�'�>2��v��D�������s�5�ϝ+�<1=�T�;�(v�+��ʢ�/�XQւi�Z%��`�M����t{W��68�<��{M��O��,��
{U��,�W~_}�u'�����]��c��﮳�91���<c;0�V��)����gg�TyC_D��	>#F9AK9���NI�F�m��u,��)h��K�N\ھ��?m�ė��뎄rވzzu>� ?{�
�v��:葋� �ղ�s]��ľKҬ������緿��|�����t�X���񦳍��h�gyzt���gW2Z���.J�
ゞ�8�����֎vU�x�������?@oh�P����6$�d)Qz�dV�Ծy�B%�Ñ���R� �"��2�o��M�O��t)͢��xDoa!Jؚ�����X
� uL΂A�աL)���	�J�:�,Q}��@.6��6f/�E���+���b��� �;�����	RF��ʄ��9�LK���>!VYD6�3�Ú����E[7w�Q�4���v�
P��:����t�򺨥*5s�}0JұT���Q`��v�KB�Of�:���xNu�z�D�@��H��/���E��o$I ����u>z����������u|���m�u���:�]ob � ��t��]k���f�M���;!1�'��6�����-�Y�*��nLe\� &�:����z���^ke���t���{���+�2Ԭ���;�Π�?N>�f����[���������׮c^��E[����I_�~�@ײ��W?�D�Z�Ej[�R�`p�e�c��P���̤˦���
����ժ[ �^ǃL�o�!?}�g������e �����q��ڰ�g�|ɣ��S�Mp�q���))U���z�a�1p�2����ʪ�/j���H#�*��S�����+(r�8�'��,NDJ�/OAP�%�P��<��4��J|q*/8����S�y�A�a�n��*�3�E�Zi�K=�B��x����J.�E ��<����ԯ�iϢ��1U~z��3%��
��a�!��J����ʏ��vyuq)��M���d-
FӤ���Y5���Ɯ�c��Q��}p]���!�E��0��o(C����˳�F`)�����!r`�Z�<7(a�)�=s@d�$/=���B�虔�y�I#,�*S�q.
�$/y��9#��bE���r�(�O���[�"�c�(�S�a� ���#5/U5��XL��U��()hN����1c�1a�P����zC��<xx�O��������(RH/ �s^ϤP@��Z�����0��w���ѐ6�L繶/j=g�~�N�(�M!C��+�h�6$�I-��l��~�i&ǧ��3f7
,���1x��o�#��h���R�4퍬X�����cO'���C��
@�jN��U�V@C�8�<�g���:�8��hW�\�NВ2��K�#2�%�	������e2f��e��c���}���/�>f��װ9�s�+�A��4�u����E]࿨��MC�#ŏ�Äc��X�Gwى|WbV�.�o��,OJ�;s�'n+�Ko�oq�%���}�� 2�2c<���=*ݍP� 3��w7�~v?ۍ<�v��_��xMq �������񱪪\z޾��Y�A�E���Ġ}�kq�Ï�]�z;��}v�TΘ2�c���$���$y������k�w`�`Wӄ=(=z���F � � �t�+��DF�I���ɞ���w�w�z�|]�>
Mv��a�����+�g]���ڟmd�SU;���L�� ���u䪜�:� ɠe�Y�J��.e�����5z����v|���:�}���d@ܻ'Ϟ�����o�޵�L]�rY�678�7 O�O?��A����I�
��Fdv��"�fu�m�t2k�ӡϼ�3<+۫!E-��{�Y���@1�z�f���J+��'�Դ<0I�n}>��zb5��(����p|N�D�̥�y�F�r�����dT�!�Fk��I������T��Y�'0)��T�N�i5mͩA��5��9� ��T�e�5�����<V\���<62�4��|�||�y4%�.��ǯ�ѩT�<:h�E
<4�q�[�n_4x��� x�C�0���jto��*i��=�s��"毨.���b�Dw)'���Pw[�����y�O@�D�E͘=���]"��Hk_����/�9
v` jc8�������gZ(�
Q,@
b*�`�	deA��$�@��ق�_b�:ed���?(7��p����\88�ޥ����.A!gu�4H�N�Pz��Oaf!��UV,΢Aa�%j~�f��,�އ���@;O�Ⱥ8���S�|�u���,�����)���c)��Z'����L�oD�vK���x��c@�a`�_乧T��,<�S�0�9�<,8��o�&�+v�����<b�sw��2z赀L�*U�>��98R�x�X�`Ò�n`v����4V>�ż�9�'�T[%ڛ��f7�����8]K3j�l�R�<M��fe4��_�o(s$��z-Rퟳ�yv;H^4ϻv�k+y��1��8B���H{����S-'����}�@�|��o�,�2��N|-
v�z]�f �]K����˜��y�·���͜����ApG�kiJ����@��Q��ҷ�h�NiBJ(�_�>g���,�k(�*5��Q}��7O(��j���o�E��h�?8y~(kl�S�xri��X:��󯬖�a��n��\�,��e�g��J�R��R��P�13��hVa8o�����~c]����<hF�[��E`ŋX�I�
��K(|���>��ڔ�z�'2>E�Ck���+����;o�%��կ�<x�@���3���gg�+dm=���J�>"��pF�L��58��a���v��R �tF��Ɍb��o��+�O	-��,5"F�Zh�`���@�KV��t%��"-��8Vm4Rr��x�]LsJ%	�=TO��W��\5��T]A��
��s\,L��"�`�V*��G�D;��Ou�K��Rh4��x^�&9�5�� �R#i�����e�C ��ZF'u�����k�ړ���������J��	�}��#&�h��S^�a :�Y���	�!�$���<'-��J>&z��魻�&��3����t6��{��>�]��k���_1α`�W��"��_`�#�ik�tj��p/4�:���PiD6,�Eū���XAA�v���F�E�ch��T
��0� �x��mY�@�d ?T�_�rK����V�z�m�_��0>)|�5]g���|A9�D8��?~�N���_Y�8�;p����/~!��[�&���Q������c5�q�g�X��O�`���>{��e)Ogr@+ԝ��a�R2�Y]�FII+ ~qt ���x���^��)��9�#�1�k[\@����Xö��,���쪨,�KH���H�yN<�?�P9�zt���3��_Y��h_>���po2��w��8����G��ڣ#ID��(t*ޗ�T%��+6��s��Z�J������nôҌ+:�<Y�#��(� h�.5=��q8���QL�LD�D:�a��6$�څy����SfR)@��-��]��ݢG��*2�(�~�<����So`�@�q��埋�	� NL��:!1-ŷe��.(�~>�����ZkJ��8�̹��D���nv!>�8�����hyb@�36�\f�1g�JL�Y,b(�yU�D��I'��Ee�O�M�V7�egwW^{�x�1m+������^��M���u�z���_Y��Ϋ^S����c��d9w���u#�������?iޫ���Ī���c����5�w ��|m>``����Y/�F����� ���cލ��>�8�%�?p,j:ޡ&��ų�n�c۟�xrJ����~-{�}J'������Č�By��n�"���O*����?�M���fB�b] i�J=���N��)q{��e���[0�/�^ډk{?�+\h���!�\�YsA-ݬ�ˌ�v���SlˌD�WZd�EOF��5pS6��I)_�P/Λ���l8^�3�|��b�����6���q�Fֽ��|d��s�5N��<ʦ�5~��%�Z��2i�մi�4iw��^7-�f����q ��c�y�s�|"y��l��� ��9Y��Y(��%��4;&&�0��ƣ�T�e��÷k��(Nk
���|}�M=�4B��[�XG\VT��W�ɫ��a$as}��6�p#��/�dc%8٨�߾�+���0�'�����F�Cy��-��{�ӡǂ�����7���������LG޽{W�i(�P���
�����4쓑��Y�S�Ǭ�y�;2���<	NCD��g�NO�E��>��#�=�-���+���Z!�oܐK�oʳ'��p�p&�j=�;з��"ܫ�C>��T._�f�9��Bs�V���b�ͳ#Ss8-�482�p�j,՝/TQ�	r���ǾW���\��#C�5Ǩ���YYQ�ѥ�0� }�]�����[q�c��|yW���`Ɠ����/���E�k'���g,r��:��:� 6���-�'I�ij���)=5 ��V�q=_������hiŃ
�Sk��!�ҢR�b�{�F�>�d.�r�� �br��^c�,�T�X}UUKAm���z�׋e���D�^y���S�_�(Ņ���ݡ�t�?�w����2	]� �n|��9�1c����,�w�y�kZ�~�}t����;>��fr�x��}mǼ@J�4xl�rb]���J,;�K�M���hц"TP��"�Oek��V�=x@�~���̦M������.����� *�Y�C4��B���_�,n�ך��}mY��qR��V��De�*S��
������>�%?���Q]�;Z���cb!kX{�0Xf�ߨ=`WT@��,d�GJ��������&lnn+E�T�^ڽ,�n�ue{���k׮��Ǐ����MŔ9fA�A&8���1�͘�|섛�f�6���<�� �C�Nc �~F]L����,�b%<�N�5��k����'��x+0.�u�m�m�6Pdz��F-����h-L�@�X�a��FQ��4��c����	'=��9�U%.�H���juЕ�6j-n�I�N݀��D�c#�}Yt��s�B���j���<[Liҝ�H�I+2:�\l�ccO�,*s��� �a< ���	)4�|P�f� ����C�h�G	�4m�hɊm>�J�:,N�����9�lg?Y�<�Hi��D�d�ڔQuq+��y�V��N�5�K�����׋h鋪�a瑾���!Z`�6o߾)�����K�9g&��sono��ƚ�F���/%`���׬ևAz��R�&�zL׾��7�׿���@|/U*
��������p� ���WF�Fcr}+��Cv��Eؿ63� �5���?zM~����z�������3'c���ʣw9�򴡂h1t?8|Z�"��ʺ��-��W���f`���F+,��ោ�j6���A�&N�����*u	�\� 7U'��J)2��"���_��x.D�SD��iӴ���{�|�Z!p�1O�b*o�yE~���r�ʎ�aQ[��Q����7��B*��������g\�&Z�3R�S�!{��7����KX��G#�s���������5}��
��fI󃥬��TD�JLc�G�d������2O*pl�zb]8E�⥇��>PY�s�`D�d�5��LK��҆[��e=a�˗���� 8���yP��d8Xe����H.[lXUN5���i�Nbs � �>�.�qD�5�;�?N�Ϙ�,���ϲ���(�2�y|M1н(����7e��n�>vb]�.P����ق8�,����M{b`�NC�9�͝���rږYJ����(j^h��:clΪ��t�:ؖj@6ׂ��Wõ�"M��`�5s�@
�1G�ww��@�?| Ž�?�<�5��n��ЫǦ�	i'�49MD)�U����������n��\ߒ�bȱ���T������y������nk�d(B�>~\9��'����V���}��� �3Z륌���@��^S K�8��Qv�����I�l�z�
k=�ܻwO�QA�+�o2�3����l!F�s��p
 W�}x����6��۶�핆��b���9�a ~�(48Re�`e��.�s`F�W0�K��M�����8k��� H= ��+�yږ:��J�"$P>����9v�y:,a��m�ډ<��bý��'G�Z��N��w?�,=ȳ�s�.��̀/
�����_̊Z�16p/ˊċ'H�tt�J���HkՆҼa.�E#��&n��J���ׄ�`�� /�uq$��X"˟�ڨ��t?\��ۛ߯�����?:	��j>���_~!_~�'>������z�lno�O�siW�~��`,�:>�
�@}	?�[���+���������>���7oޔw�����׿�3\	��������,��B�������}!BP!h�?y�n����u�Bg�����v����uvh��2����F�5J��z�� 2�G��V7�ꜞ����	���G�/�,k�$8�34�
�c8��Cl/��B�y&K�"I�	����rg��tbşE��3^��ܒ��_ʭW���2�ч��h�N�n�Ep������*_�w����9�z��Ȯ�;�4.���pݷn�Z �pB����tv6ϵ2YJ�)U%�2����f���n�3��I/�Ϥ��H�d�_�ɴ+t��r^��|6-��S�ae�=�?��l�:���9;��#�9�auj֌;@�\�M��˝���b�,3�,�Sn|?]��Ɯ�?�81�{N���Q�c�bt��/�]�ߏ��
_����:#����W�{�w}�ks�n����߽�&�|����Ѩ�h�,�,�$gyh�Y]�*m�� #3H��#�K8�E
({�u=?!��`���>�W�oC����F\W�"����-�g��ءA�~��n�RG�w�B�y\u>yn�Vd)<>��\��i��t�jt��tG�qo�����~����ˋ�}\�b����L�N*���q�@�< ���Qk���,I�t�������Ʃ�{��3)�O ���t�y�04�V.87Nړ��AJ�nn-�K�4 N���F�LӡV��(P�D�X����D9�"a�91��e�'?4id���(�������,��z��|q� ��]��A|$:] �4���g��z�tv�����ǋJ�@t'M�9���ʎ��6x�he	"�ڍ�/KUf�!g�҂>*�! ���3�x���A
�/�(<҇���sl;^�P � @�oo�)l�I��N�c�S�K������П��%�׭���n�,#�U����^�-�lP��c��������]?>=����SVWG���ѡ�=y,W/_�y � �
W�qAu��B>���ͣ���G�����r��M����`ޮC62�ޝ�-v�(�݀ћLNI�qeW��av:�D4^쇱��Jx����d6�:���!���+W����,�	�L��U5�iLPi�s��"L):� ,�������K���\D��'��*���Lr�Ёw��k�r�h̆Se��l�*ޕ2���y�}ƾ�d�I�������
+
^��N���E-�7$=g�~E:��R�&[] v�������q>dj���K�M�l��<�X��73�� d�H%�l#�l�U�\7�G�;rU�Z�煪��9͐�Y��h���ʇ˨������M���hT�R�/��<�\�+CF��Q����bC��eԖ̔�ܾz��)-��;(�W�?������F��E����rĭ��G����۲�Ll�[���:��]�E�ߗe�M7r߬C���ҽ�q#.�ғbQUu$��I|����o����W��%�P�vH�	r���ڮ �	�yfM㬆v���ќ�mP5�}�'RNM����/	�x<��nud=1��y�MT\߿8�׬v^���|.�/lI���SϠ�< ��К̩]�g�p�(Y��Na�;Ǧ�=��D�ܟ%���o�G����	Y<ў�ӎaC�*� `�"[D�BL�ԩS�I�R��%iV�jKҨ�s�peX����],�/ߦ_e��sh9��Q���..�)�&�ɰǓ�(UA&Ir�f��dm�+�޲�
���t_I}L��vL���L�/ ����r�����wg��F�c��b�{ՊH�w�a�Ĳ�7 ����G�����p=-��P_�b��Y��a���>�iG_ �|D�����'�a�����QK{4��W�l�V��v�&1z�>[��&H����_��o��q�Kn<�$1M����`A�#X���98|QW��x&7_}��}���� m�o�(, +#*1�b���|,�}��QPj���D1�YX���{t|�H��~�y�7i(�￐���S���Ύܹs+ �U9��� 8�w(4�s�Z�ca�@����ٻ?��|���V砿 �h͕�p �e ����)Dè^��(Բ B ��Q�ft8����0��g�+ܷ:���x�7OKk���ap:��H�"k4�Zha6ǣS4,Z�s���Sy���p�e������E����S�����z�K�ə��dF}{]�j������x̿O¼G�YobR7�}0�sl�	�2��Ʈ�߸7I6P��ԋ�
��wѶq�T`}NU2R��4�,t��c��]P'bQ��$(�T��(��N�?�pLo3K~w�� �X�7-*�3����m����� ۖ���i@��NEϱu��qD��c[��M��A�p��yP�x��e���.�k��6k����ڻ����}��c|��Z�Ǌ�������׺Y��|��w�3��Ɵ(x���>�K����m�׵GI�b������@ �Xin���Aek��Vz�0�L�������E��vD}�`��ן�szy���w�q[��,y}�f�aS�����٩���֯����2�^kbQ�^�q���a#��;2a9�����PF
��<���֤��m�F��<QT#*C��9�|�NT���܂�ެ�	�R�u��䩠�w��w�SZ^$4OIn���v!�?�5��e1 W�R�`�8oV��ND���
9S=����`I���WH�*Rsy�J���h�.s ��sD�/-t�c{6m&�{��P�gRZJ��Wz�s�/6p D��E㧽V  ��IDATV�w��/f5����9g��;�����)��&��}��8@DjB6o.��b܆.�5�N���� >N]���&#��5Pg0Y�	��ln`��_��,�e|^����{��?Ƌ�@
MwX����<D�^d4��9���]�%9�J?���O%��#�k�s��S��u�]{��)�s�G���X�+�T�����JkBz>�� *ǯ�&���
��` 7��Xlt�$� �WWW��wߕ���/�W}:Ϟ>�o�z��AO^{����������������[7e��ݰM�loZ��ȋ @������D�~0��+C*7M�y�we��e�'p\8 ��:��]��x"}(��q37&���41 _jt��4��L{���^�#�����EM��'� D��Kx	@������/��k��M9K��d4��D���(�Es�q1��9�+���q�I��d���[8	 u�þ�,�);=>
@�DA��l8A󰀝iTs�yp+kL�O���s�STr��f5H��͕zT&�s�l����֧`��7�E��i&VЇ{�@
�V!*��j�Q�)���S	�Y�}�����q%����}�L��q��HX��#\�AE�8�O�z������ҝ����k]�, p�t �tmQc�b޸����(���cYd�k���-���[X�������[�.]tN]�M,1��Ý�.�>����1�����%q� ^'Y''�z��Q�j�y⠦�R���~o����1� �NNec���chN��j� "&�?�$x��[����B)r~+m}�@���JW�S�;�Zg0�����[�k�$���c�e�7�;P\_ɉ����r:�Vi�v��#��}gp&,nkw`U�_*!���\c�wǳ)���8s�������������o5xw1���tj+ǃ� �ډ�$��[�o����J�1���?�~b�5�9u��@_��2�Ks��@z�D��:2Wؗe3��/���[�)#ME����*	S�i����E�.�IS��>і���i}S�ż�%m����.]�֠nGc�I���~��V��lR�K'X%��k��<u�K�GW>��Ū��!s9%LL��g4b��E��������z��ߌ�OX�ܺ��%5?�I�H��d�g��9_��9��?g�{���ۼm��2�����[W��^�u�U���gg��A���A��ð�Pz+RbX_�`�ra��jJ�#H��1���t+<��/�}��vx��!CT��W_��7����%u���ѾXZ���M�����M���~N��<�ӧ��uP��% {&�be}"5��<�u�#��s����>��uF�Y$W��%Z���)2$�/A~�EHd�d���`K���9�a�>R�a�@�����bb�o}.6�i��y:V�b�O��>�3
��c��)C2���P ������@.h'u��!W�_ō����^�P���l���Ϩ >��m�
����E0�3�JGCɇ(�3!�R��C1��tL �S�tFg-q��n8�;Q��2,�ga�=	��È ����D����=�9"�2�Dm B��Ȇi���t�LΉ�E�ݹ������[��mUc[����.
,tA�2�����,sL��X��� ��]'>F�~VUq��-����$��������qy�EQ�^K�&s H#C�N]�:�2�Q϶�j���[��<i8���?�w7���rtt �v����Ĭ�j>�GyC� �i��+�5�Ȏz�}�����E+�2� �9l�H������;�w�1?!N�m#.,�l�q�]�6�����L5؃��<��F�5�[կa#�=9���X��2޷�%0�+�(��>��_nɖj��� �
��sK5�D�t򾋤ؼ*U�4�1K��L�e���uT�!��4�����9y�<,`�Zgrm�W)w��t��"0����E��o�4�^%�ËEf�ECeE�NT���Q+L�
�$q:όb���v�]��'m�V��&v�ײ<Z&�FGU����[��㵣2��fҲ:7h��'^4�0���JI���Ǎ��I�N��?���ےw�P]��4O;��Ad�єB;*�
��ǓV�C�N!4�GG�_Y�y����Y��!�9u>��߱��|��ߟ�5����".�_b㱼π�����o���$����� o\S����-�����Qp8�X
8oP�	 ψU�ṀK�/��W���F��O�a�bsu%cS���� ���(���?�Dnݸ)�aOn^��G�2�vz|�ώ�e����5��,�
Fu�E ��r�Ƶ�tlSO��/����T���g�����P��>bA.�0U0Ŭ�r��&�Y�]iѬn?\"0�[+�d���V/-s��Zln�bh��j�����z4������I�ϥ�]�/��Ϟ���*%�ЩQ��8�Eƺ#t#�
E�t �p��ɏ�Q��P �Z��� ��_	��Ǥ���lo��,�~���ZTO�!.[�y�Χ�.�-RK��j2�&�OAyC.�̳GΉA;�2�62Ȉ\�ܐ�U�),4k�A��X���X֡ ��WG���k���#*}$�v!�P*�ן��u&�.�ŀ�fc �m'��2���B�e����~�sXQ��36v��i�G���8(��{/�Y���˜�x�(�_����S<������ߋ_��iΜ5�C}M�W���mr
4�s�b'�-5��\Ct���	��u4�6��O?��0g_�ѫ��+7�1}/Pρ:�F��\Ci͘=�hF;j��^�����;׌D���?_��r��m����3�E�����0޹�R���}�s$��S�({G��e����l�
F��S�Bdύ#?Z��悦\�@�^!��6aR��q_�ؗ'��*�gwk����:�
mԃkQMM�{��QQ9E,�<�;R��S�V�o/K�i����-��#�¨i�3�R36�P�E�Uyi���}������*���>�� o���t�s�9��EnS�A�f=��p��7���GYc����/��QC�'�,��z�u��"E��m/�u�|����jW����nsW�����s�#.Md���Q?����E�ʬ����@�v؂R���\����yR�ɼ@��(��\�J�A��G��z���KIk9��f]繃��ң���C������9�Xe`��t�����K���3�Q*7��&�'���l&���#�=Ak��?�R�z�IޣN��K�͎�=an\�tU�z�-*�|}�}�ŗ����u�7�ia7\��৏��_�
Q�r�\͜�9b���CMs�Q7�׮i׽gϞ���Y�����a�d�����hJ�	״s��
� dч �k#6d A��3�z]84U���]��}f�6��`\�{`�>�/��Yǁ����
Oh{c]v��8�ᝢ軲�љ��E��P��� ���Řn����	�"8p�VG~B&��ӧ��z(;�y.u��9U��~˙L'sk�RЁ����)|ϽCϸ�;fMk8K-��Fapo(õux�|���\�	�O¹�����p���W�W_��j��S������RpmG���}�d�(���\gM ��Qp��AR��Z ���c=�k/���Dv7�M&���m���D��`�?S �{�N�E ?v8|�~���?�uLt�����c��=T����g|ﻛ�봺:�1������.���W޿4k�V���tQOҾk�9JCaT�n�Q�t��lp�M��\��c���@�����^�_������}��@�pgk��1\#{���1��j���X��l:�հ����S�t�:'ݭ��NQ������h�����r�t(���9n��x��	tH<�ۀ�C��l�d�G�"�߳s�=w�l�0���p߁W���ܐ˗v�d���Od�iҦ�/���4��!qkN��J�%�����ܬ����:����
�~�g����{�jL���)��@&�r6Q/����p�T�I��3���%�!2�o1.U�������3R<+�Z�R�ЧZ��!J�i38�`���v�ћ��'Q*���t(U���d}������ͽj�_�H�����Ҩ��&dG������c��we���}��w}~G���\4�F��߯��9F��y����8"c��"W ���-��(6̰X�s&[nc�?܋o4 ����<Y�s��x�~�qӗ�|Y�Do�&)k��Ӈ\4���V����4hYŇ�ȋ7sB|�E1\��G��O�X���9
�����������'���<�_��Wr��M��O~�Փ��my���޼�kPm�����~ ߗ�^b+����c�T�5o�D��|�ս �r�����rz2f[�MJKb�;=9�u*�+k� =�n������4~[;� Y�oߖK�w��6���gr���� ��{�?�#g�?����)rV=C����0�v�>+�����8�������Фɫ����02�
N�E�����" O�b=ꅱ<�Z-y
-��9h���Şܼ��y��������A e	�"���Us��@�T�!������T��gO|M��h�G�|Q�ҐB�����	µU�\�����?�n�5��pu�z�\@1&����^3�o���� /8u�K��P�J�-�9OͮJq��2�������+׃sy�bV8\�Q�`o�Ŭ��E o+��S笐U���ބ��uN�oDo�z{��Q>V��H���/��Ԟ�k_�nS�E�=���x��Ψ1@��b�;�m�z�y�9�����S���.u�]ҵ��������3=n��,m�KL��sP 5����zb����w���K{S��B� Ui���E�~��3�Ӂ��*S߳,�rT�*0���3��ev@/�c�-������K�v�2�����r����lVvt;s�bH w��(��j�P�R�P�:�f�٘O��R�U������� d7�WF�/r�����Pq�KZa�8����2���;��q ��p��rl��+��p�ӎ�_
 ���P��)ZPio�2̱V޾}K���k��c6��ڐ�_�T�/�NHo��#:��ހ�K�>�9H����9��(�j)3(���g�����(���1|���ށ�%ۅ3|]o4�Ia�P�>xX㙥�L$�mXڲL����#M�Ff��Н�Ѽ������@�ϯ��K~+�k�Ս��~A��N�¿�}��l/����e��.�����E1��˼s�_-�# ���d�[�\G�hRQF��4R��1H�3��:+�p�I�z��1������Ҩ�oE�Ly).� ��-�'E��h����,Q4�ǋH����g}vP��`~
��j���#�,X I�~��xĬڽ��cyđ���_ɥ+�� �F�^�^�&B_�v���!w�����i ��=�[�ܒw�z�4�w��J���+��;�7�6��V� �3E1"��i����]F۱P!�����J�J�u5�:�!��'���@���7�����zgtE��ZQd	�tоn����t������w�����r�ҥp|��S�Y����>�#������W0Ӡ�.�4ͼ��\Vs6GB��o�3u��FiP(�㣅8�sz6�3A�<5�N���
a�<�?c-��]�{�Y��\Pu�j�T����zC�Vԕ�r���3uJ��{uc'(/T�|)��EoxmA�~�t>�i�0~ �@��+��S�Wb���"�t
���L{�r�K�)�P��u�eM(֐� ��yδ�l�&Z�����5ӑe�O�%�)��3ۦ����gk���iJ�����t�W�y�&)^����]��ض7}Bڔ��G��u����D��z�^��#�����s�l�ڭeűi���w���>k��g�m=�D����3�U�˪�@[���)��3x�i@�~6N5��2��4r8��Ɇܼ~�������ۿ�6�Y���\9���D�؄�`�KM�����d<V������_�/��u�������9SͳT�3����C�]kAǳ��g�5�5D�]����2����	uC���yk����<�g/���t��Uy���1��7P� <0��¤�=:����$�R2L2�)ω���D�'ߋ~/�� �o�y�aZ�
MNpSX�;7���Q�j/V�	O��S[<����Ĳ��0�H�+S�n��k������j���X�L� �"���̷���ݾ�@�(�^���r~���X��I�5�����gw���\z/f�V�57��S�R|D0��s���>ڒ�'l;��腤(��P� �҉vl�y�H�"�[����'�m��1����/��K��Z�1߯z �w��B�i�`��=�����ѳg���)�h�����3���cfǞ>�g�����S�L���]D�Ѿ��K���S�����ތ�lAލ`�QĊ�������M���W6W	G)�:"S}D�l�,�{f��=H�C��EE�C<�Qn�� n�A�iӍ�:�znX�(S62J>>=	�� �>���bS�-{���Q�в{�h�?I�2��#Ȍִ������sHS��*�1����<�+u����O���=`]@��+�\�@��t��D�Ktذ��rqZx�E8:"���	�Fz9�'�AGe\75�a�l���\��M��\1��9��
��ar�CTj�C汬l�%FC�RD��^�q?@����J��t <�$��ɀÈ1���,�A�e�t^�(���r;����SB���%kK�z��yL����������%^K��ۥv��Yv��w�7�^��F��s��i�^�YĴˮ]�ט�<�X���☣q��z~^~-�'e�hxč�ZU��zs��lPX�K�˶�X��=�G� �^����8���Z�#�{��E�|�$�������ܱ�>{��R�~K�����Ͳ1zιL��6��#2��6&�������#:�"��Am���X�Z��:X�����z�(�����)�;j��a��{�� gI�dd,3dd*�6dEj�E$�,�F� � �wƭ�3�?o���g������'��y��[�d��]?������'aw".��/��*_S�ߋ�u8^6��זe �D ܠ-����.�'�Å�\�}�'^⻿c��˾��`,�������}<�`�,Z|�r�	]��Wv��E��?�L>��'���8 �9���,x�3�j���J84M=A����C��՟�̿�~p����y*E��/�54�� A<���� }�N��R��˳��"1�t��U���=F}
�?ߗ�gO�f%�g����C�����6;R��e�4�������S�o/��pv|&{{{��y;�*�Y��7np�;�f�E!z��T���exD�����¸畞W��B-���/D��)�2Z?2g�c�r�Ոp���_�n���1j����w��6z��1��XV��X(�Ź��U�}�Tϭ����hEN�~�^�q+k#U��k;̇��)�+ʧ-�h�++C]�����
�iOiE]�಺,��t���
��(v�6~��@���_)�;܈�yu�㨤bM��UF��{_=�2����+J�����PҲ�f}яxm�6Ły�}9�t��Yc��&��p�`/4�1����i~��Xf2^���f�M��8�����^�	P$!J�%[�<��q̗����o�	��E�d˒,[w�  b�[oU5���O֩���{J~��۵de�r�9{����3��-}��2����Zs ��n���?ePx����[�7�u����i�a�Xs�aB(����	�;�aI���sq PBa�=�����>w�5sCm�5L6���j.t�ڵC�OX���q45EV�&cu�e���S��Q.�ڭ������,����g��t��]o��:"fs!ξ8v5��Z�����:h�� @G�0�5�`���k@c�ú��.�Y��?�������o�g����!�	���5r�z�5��w��/Ȟ%ά�>�!�m1�� q6��0cMB�${؇�x�sM������U��r�zc-�_��"�^����E�9AbZ��T�}|�|��b#���.�4�Cw}_��?�@+���c�v��cl���m`?�[s<��ܳ��a��ܵ9�JJ��L�%����r$e6��� t$�M&�o	BoM|�hٸ�o��n\?v��{���������C�%�w��y|/N�u |��wH���	��S�r�5 ^��){�"��F'\V��6/���]'*>��JU�uؤp`��U"�H:�!
H!�"!u�x�\�	P라8u�'#q8�!���|%u���ƙ/7E:g���?����H$��~�nx�	3*hО{�N�В<~�D~� �܊�CiJ�������!=P��6!� ��`Uw<�s����FElU]�8א�~������l���φ�Gl��]��<CPG�6���XF=�F������@.�c~cs8� �t�	��@��v�2���,�����Ԩ/�wG$��.�i)���3��~��s�_
�g�a�.��^ x8������qO���gr��"Q�}^��4���3~��=;Lm�E��@i��@+Z���U��*M`4��Wq.H��� �d\�S�7F�R;�D�����t}Pl����) �h\w^�]����n�9#+l�i����T�\o�S�Y���x��%s�	Q�����#�><%���L����l_Y�(��B��v���~�9�t��9F:M� ��:��kkeb}�<i��&J��ǃH0y�8���5+0>~���ו�1"N ��P5ؕh����k�wK��󈗚�
r�)W��:p,�xJ��6����\��*1o��:��"8�����xD��i|����8~0k��fR/�A��g`Db������w��ᮄ;F���p�~㦴���w�1�����#�Y�_�"y����tN�,�}2o��&��BA��jP%��H�-���ٟ������4���]���Ĭ�.k;��L9j�t�s��`���;6T�*ô��@>SrR��{M}W�Χq�g�lҺw�7k�I�O��l�&]5ǁ�;Mh@� �D�=t��,��b�h4���t�[W�\<*�E ޽��;:�s�ӑ��>v�|������4�- d�y@��g�-�Q��V,������*���H߹{�ݨ#��nb�HK�&&E���X2d�v��~G�͐���o�;���N@�H��u�����<��KǅH�Jw|�Ѝ����q�~��lN�/�I�L�Z�a �,������{�衻8=�
"�yC�"�oD�����*ϱ�����y�����)��_x�@"��Zu�S׋��$0X���zw*�ѦO<����b��9q����qg��M���%��j�-zW�F��RC'@Rϰ޿��{��E▯�.܁�2D� ���;��� ~H#j�3��B�f`���G��O>҈D�e�+���1]�!�&�������ƩO���f��F~��l�*0���Qʚ�޶�q�~)�i��Rd�t�Im�˨}���3Om�y=C
�J
�0V�Kp���ļO�m�\JW��9&�J�k��c��6�.��
�R`K@��_
�s{H�<؀}��ն.k��;o||�T�����u�x�>{T��a<Rp�u��{��JBD>C��(���uj�Ҕ����Pi[��V$�e0�B�JdM����� �d}.1e�zh���S�*D�
	3����i��m���T�t��3���v�����jnnJr���q�i��b�4l8�?��c�[��)]��2��~gG �k�_��v���7�A�����}׎����k����CɊ��ݷ��"���LE�~��u�R�|D�	���-�Q��4��_�?��H�*ۭ1$��0�e)�T���kp6���T�	���&B��u��f���ZLi�N�eB'(h ��M�����-@�ρ�u ��d����M��m����ٮ��=7UKxػ����Q#�"�a1�>�ԫB�����Lv�n�4=r��q�����;>�w�������w�eh'�]1�X�D�i���l(�Ge �9�S1:(�Y�S�F�K@g�8<�Er�Ἔ1W۟�xc���!�hƻ�~�{ ���*��%�U�Dws4¢9xccc��~�@�V8�tI�H�ux����o����'�9a��������/��09�G-Ygs�޷_�4�|}�ᇞ��F��c������gR�����<�@�W�1���I�mD�4��aJ�A��C�R.8W��
v�V�?�J�Na�����U��K5��<�}�-�+*D�_&��&�R)�B"o)�D�@�D�i,v�DT��r4VB%�0�}���hp�df�\�Ǳ��s�����̛�{~�\�M��K7��dW����0I�t�3+H���LBE�8L�iv��K}����Z;eq&:pj�T��"�IYv�:���"muN͢�@�cY#�I�j��X�7Y��`��{��t�j�}�h��S�r�th2cm߭�+��,ͤ��F)�M�n�^-y�̰�Mh��0|������m"8��~�A��9��
��m��>j	��V6�V���./�k�9f�.vm��B߀�՘���&-�p��Vs�L�p�f�}�NN��z����;�NӪ4	3�ޮ����;#�Q�^8��A�k�-�{��iY�X��[3�)������f�p���^�w���8�-�5]��0��E��u�(�^��S��x"�������3�8��C��Zwzr.t6�))Q��B�b?|�DB3�8=����3IR(�1�+^�&��k*Z�V4�i��v��q��ZycY�wV��ٜZr�csT���U�b���ց� O��t���S�U��L7R��`}����Ǻ��h2�l�/��k��<�(�֎ݦ�ց�\?wNJ�H4�K�g���.�k�T�w_$��h�jķ~!f��S��p�:�s��~�ױt?��s��<A<��m�\`�l�q^�.�`�3��{.�翭�G�1^��88!�H���S���$���������i"�� �V0�s�'�M�uH��f+�vǝ�}�v����������$�_�F�bb�Q�f��BH��c�	4=t�Gߺ-��O�K��Ʉƈ���MQ��_��n��v<�����<���ڄ�zG�V�!� �G��ݝ�;}�BLb�Ep���?�zBE2�3sR���@X9�������A�}�J��f)�oH�$�s"QB�P�e Y��d}Р*{��e]����c�� ��'�f1�
�PĜ!�d$l���߀
��� H���)�
�������ԵfOx��P��*�O�>���\;$���͛�i�`p(�b�K��I��AN�W�o�J��m�^��:ҏz�	5���*�;g��>���1�e �y��o��Z�z�Xl2���M��3 ��TZH瑭[�u�?�k&�g�$��Z���X�q���'����b�n���Tm�\�vJ�J!�9�Ĉ���*4��N�I~�,�遳%�r�bԎ4�Z�y4f})k�[�����^��Gi{׾㖒b��1��=��!JY��5���Hʲ±S�D��I̎P����#���7�|S��M�q=��	��jW���M)�)�2l�ЛBs���S�f3��4D�I�JM�j'�	�[r~�0?+��mUN��d�UٿQ��6 �$9�hܢV�l��a�-)��6��W6������������;[G���o7 ֓y�M���D ���X�t1]�om�?[W�0�s�|J����a�1z�B8�LA;G$���j\�_���X������Z���Wi�dj�9R�������d������dv.	jq���ho�-[��N�QM�4��eֲ27A"��Y"�*[�(�l3r�H �9Y�x��m(�lc2�@���N0��M|Qu&���`όe+j?n���5m%�XBT� �&S��ى���G��k���޸�n�~C�&׌^�� �C ��+>�~������}�������W�S�F�}i��,xL�F��(߸!u!B���nJ�@Jb�H����/N�7�z[l���gM d�za�±y���jmH�t\�佰�,�U�,8��8̃��d��0�~�{p�R�߾O�n$*�V7���<K��߫U�e
7ꕮĞn���NU�se��6�BGM�V�� ����\�x�8C�$����g�E9��6�tH��@�NSfC�F�b�u�EX�Xp|f��, ����(D�(5I�:��C��ݔQ��f�24�o����~�Z{��&�9ZO���\�g�{���Њ�҂L����`�� K�\�������O��HZh$��}H�-�f_�X�m�������g���m+��b�-���?�hw��$�h�ع#2L0�B�6��q�B�uX~�{$ ��Gfʵ���y������~���	�<Eg�U�M�(���aI�k�s�_*{R�6�b����2vE�cL��bٹc$&K�~�4[�L86SG�42��EM��~F�K\K�2>a�D�w�o��}t���=-�Y&b���C�5 ������meļ"h �ǖ����*��B :�>���L�,�	�XL�`��v=����i�J\���N^���Q(��*r�Mg3@�c'�]�W��+9��=���c�"�p�c)�]G
������Z���'�{�'�r}��vqxߐ�䞵N���\�h�f���q�w��w��	0TmԄ )#�k�Y�GH�ǅ:�!1̷��z�O�[�ɗ�<�k%��4�������<��ݘW�I�I嶝�Ts�u!	}~�����R��%c�ѧ�zGA:�d C¶6!�}������_%�`�ņ��HB{�b�V��ж�>=u�?�j8��Va>M\]N��b��3w���"�Xm@x��T�-́����;����X_�YH���H�p�K��*����Z��9�9�\���K�������
�,H�	F��  ������"��62���	�:rv"7�jO�#q����67bQ�Nc��L1ّO;R��'Fj㏙�Z\��A�B��Y�li�:����L�H�;��<�92��%׊a�4�$�[@>�����@
+IN�d�\î�uk��Apӣq�N��~��w���	�rR���z��u�;m�po�@{�s���u��Z����m��3m_�DT�>��c�(\��h��Bs�D���zϑc}�M����=s<[�9������M�S����ϟ9W�6��E3��l�
)L�9fMX[��u9��G��M%7���Y?^K�t*4����B�ip �s������*j�P���j��q t�.���Uk�5�9ah��1����R�� ��x�D�����i�FLe�C?(�-#���bK�}�J��}��Zi��0\j�֛�,���,�"hE����!t@��v˦I�MXn>j��m���6LL��n�������7�����P_��DNZ���Gց��m��M�3l����{�[^[6�|��	�_�ю�q�a'lWMJ��!=;~!��缿�o��O��/�g�A=�+E��N�v�T~5��Zs]���_��3��[ܞ�rr��+�(� _	�<Ay���H>z+�uE4��&��
��8��x�l�F.)��#1J;u�z�^�����+���H5Q"ޥ�o����5�'x���c��&�]J13�����'?�G�H$8�j6�R'��<������^{�F؝��~>�d��7$�@(L�UA��C��K_37�h|���]���L����P��h%�K �&RͨT'˶	ڱ6�_/��{� m19��Ih�ٰM*���]���BiX�j]he��܌�m��sQ��0^��L�	1cj%��������3N�Rޡ�.�@F���3�������`v�q��|�H�9����C��{!q���N�)M��R�<���M%����"�i+�2�Ԝ��Z�aMkRp�cpH+-p���{Y	mn�a�L��\�+�uMۘ2�ӫ������7۟��m�sk�3l�/�I���r��$�.j����kN׈8����E�덾uv���P--�p�]�gb����{z��jcd�,K�� �F�p9.Թ�2�Sp�V&���K������6�"|�q�sŎ��m�%�4�2�aZ��4������OM�hB5sR5H;����.�{���{q�!%��q���=�##Ĥa��3�ۯ�a���G��8*7*H\�D�j%:���I�u^m���mj�j����ڿy]4YB���jr�8G��4^��Dg�JDb�s�J��w�{m6�XO�7��X�6mG^����g�����i�c����`�*�游{�Φ��E�g=�H�< ;,���3Q�S�F�.�n�x�7;=q��ﺏ�x�>���'p��!��{R�>�m���1O��e���릲�u��h{ܦǃT\�9���8g�H�K5�pA�g�r�4�8Ԏ��~��	��p�n�0M
��tلh#q{kЗ�.{��07� �d�}�𲖘�b����0IY6�V�,ΰ˞L�l�����xbӆ$��h������3 ��l��Ӑ,Mw{��6f�8EY2w�c~�fQ0U��U��*�4u��k##lTM�F-�l.�dG<w�6��;g�i�����z� �lȈ�!�����ԁ�%���%�Qu��\�l$)mA�j���1��p>��;6i���/|.C�o�z�	C	5:���X;x�fh�w����y�����g*I��N�q-����ɬײ���\L�jۛ�3������ټ6���ؽ��w*M��Az.G?�N{�^���o��5�z$����1����y��jh��^0�͐6S+����~/�����[7=p?���𲈬5?B�s�j"�C��Ӌs����;;$[�	�d(,N�LI�$jM2{�ߚ��>ڔ�V�o�b$�`�C��7�z� 4�޾������?�A�Y,��3��!rqJoW�!�`�PG`5B!�]�pC���<�)l����E�u�ь��vv��{"&X;{Sw||$tm:��dy.�'
����M�j6��e]�	׶ϝ�*x�J�RNR�87��n���vPʫ����:1�Y�i�L�]C��������qK@�����H�!��XɊ���� �~R�Ԣ��}�(ص�6�o��� ��	�����"Ū�����ֻo��=q}�H�|H���7�����]F��2e[f��˧��3o+��U�׊<��m<cM3� ���7&���� (E���SH�Ŕ�Ј"��O*qzE�ID%�DI��� �.ƿ��J�QCP/k�AW��U̘76!�FHl4Rg l`h�l�~�a�R��_�]!h������B���B�n=���1w.�K	VGKO��B��1�+6Q����-G�ŔN�V꽻��A�X����QH���@���@tclk��8�Z�0V���q��kwv��aGY�MgT��)h��3d��T����"��$C:_���y~ K�y(E��_��|g�]0�B��\�i�$E�^�ؔ.h}��i$�no��pG6: ������A�SED5Z�q�/�{H�����I���vU����}[��{V
 ��v�o|֫�Kʰ��TSPe�(<J�-ﵒ�>�O{-�c=�Y��W�̊�)CC���iiޔ�Ymzϴ�اc+�մ�	T���H2�J���&&�D�W�G�GjZQ��D�|�a��ˇ�%���o��޺��h�^��g1��!��Däy3��z>8�w�n�s��R�0���{86���QਓV(��2xcf+��q������ �	��}vv.�>泥d���-���w���b���ͅ��!����T��,�-������lu�����l��S]��U���(nG-���9��S7��z-��Cz���V�ўۙ�@2�1�(�TUI����8�מ�V˦Y���:�D�izqTW��4~ӽq��c��^���%�4��ͽ=�>{U �	lg�O�
x��M��>�x��F ���m��b��h���O�=B\ۘ�"ɆX�&\V!F|�Z�Q�$��E�޿qt�޹{G$���n�)n��M�F�ƨ3
��㜴~�槕�߿�bۗ;��P�s�R�yt� @ￆ,�2�5��:� Y7����Ѓ�a� 얭n��RwEu.��1/�[E�V�tR�E���i��1��h$��&��w��1AF��v�p*��6B��:;W��a8II�Uh��GaW!&��h��o��^��e>c����LB����	�8ei�+�8�I¢ō�[O"��QS2:�
���?Cb�F�.���0���"���y�"�CFWn>86�m�{sCLc�V%g2�Bl��y���[Q2 �$+	&X�Ur��$��j5���:Hڗ�Ax/���g�XЧ��}$��y���C�oE�!HgR)o��K	P�SP٧���<��tߴ��=�JO-#�ci6��~���lo�z�=����zۯ�~�3�s���ϕ�Ʀ�[��\_��,L¢�����+�g��W�x]S��\}�|��J��m�9�IX$ҔR�Y��1\���G�
�~o�y˯�3��`�3�
ݩf���e�#���h�9���\��kb�]_C���m礍��׿����o>���/ ��ޏŜ�&L1�B`�`.jmG5*�<��.
�b��o�x��Ό�YSQ�y�k��O1�;�d�ye�_�%�)�ĩG�$�k�=1y�u�ؽ��-����Y4G@�l��r��yy	�|o)��E1�rj7�`�_���R�=�bZ�ctAX�awm�x/�Ά�".��zq���%W-�6���%,}�muv�6�b	hZON��{,Q�t���:���6a,bJ�+�"@�ԎfL��qL"p?�v8!�b�.a��h��X��7�ݽo��~��O������������@��߰��ʼ���]ӵe�u1���tS��Q5�;�=V.d�l�`�!�S�&	(�(�6�*V����HCR+�,N�/��U�`�RG�Rm�Y��P����1Ku΍�$���.��W�<�D��ּ�����$T��\�*�ܠ̀:����u���H�Q�C��Ѕؔj1g9�c����l6����/e\�����~��,ř��ᥛz�/��37�8&� "�@���h3���?<p���z"�X��L
 ��Ξ0`�"����{x	��q���е(��ǥ�(F�%Xt}>=.�PM�l�acR$ǂt}o�����������g���?wϟ*p8����g�̊����x�.��k:vΣȬ�:�ɤ�6���߶�{���$�{Q���>�'�"�L�g
���F��c�*��N���3�wg��Y�g���>�	�61Q*	�zצu۶���p�_�]�?h��#ɚj�31I�Or��"�k$I�8H���e\C�b �<D��ݾ��г��O�/~�_�����0�`J��"򌄔�L.v���Ԧ*����t9����R���|�ڌO�4��/�O6j�#G�����ۿ�k~*t�v�@)�cpfU$�E�9mc0u)��<^Q�~ǐ�U�"X�a�W�7d�����_Bu�9m��t�^N%��������J�k�3�������\�a��w�/~z>.Fz����>N1p�.���VR"a��� ě�n?ꇵb}I
.�P��(�ĻHMh\1$JW))�c��� ��c����°-��u��(}Mx�9��t�G7�q�ڥ�Nz�	�+ٜ	� �C��'���������z��`Gc��+��^����{o��~��}!���)�1�?�x0ҏ@���c����ù��`����`My�*EU�}؏g�`�D*qA��a�	l��c4ٓ�J�W1���Rz�y�+�Z�v~�� 0�i4*Pp޶��g$�_�����B�l�T������V��*kB�"�\�G�p�L�ay����
9K&ik��6�S��L�6�����H�wwg4�g���h�~�"μ��)$�R�@-��b��$��x'$%r����طY$���E'V�8�7޸#�%�=Q���vׯ��|�\����u�V����E $�����D�{W�5��@e�l)�b螕�롉 `�zq�ӈ�O�r������w���oݼ�o
����d������?��}�`_2ܶ���n��@�}��T��~Ҹ土�~�m�u��5���޴��k>�֟
Z�9[,c�P�ƾd,t�ߋ�od��ۿ-s��e�˽��3��{���hd.�A�6
s���M,�J�
1�%"v�&��HW���%�k[��hfN���~��r_|q�}����?�1 :����}�f9ߝN��������d"� ����Ɏq�M��LǧC�3�^_���D�� m�-�G;b��F�{��_�B�W�E/�Be4�2~sՁ0�'�q�U�NJ�̄�dgg�T�8s�S<	>z����}��J��EF�֭[B� H������o����C.���M��o�g��|g嶔�&4�jZOF�;q.H+Q/��a[	ȕ�Q
�uj������:�tA� �{O'���ݸ����>ޟJ�X$��F0v�~�l�U2{�(���Ñ���!�_jY'@׾��I7��{(��ڔ��1�^��Q0�4��!�C!Q{��e4�9Tj��$��膌W`G����C�؁q���z%�
HAFաzy# �b@��xN�ڑ�qt�>}�A�ΑD�����&Νک�N�$���0����s?�Qo��6��:Z�����6(�J�@�H�X CK6ԑ1�	ểT�m�A]A��
 kQ���dUg;H`j��D��jτ�`Z���0�`(���тم���lǗ��9���H`��Yu*���1Z�`~B����1
N��M�{A�)�&cɑ���s��Y�_��� *	I��i����\�r�o��ݩ�������s�<h��g��+ ��cTv��p�lL�1�7�+T�
�7�L���Cٴ�ᩏA+�^P��{�T�M8`����$���t��߶�\3�;w�k��i�F/�\
����8D�X�$��d����5����4¼�A;�9&��[�Km�@�`��ƿT�GՄ���J
��Ͻ�$��x�X��<*�?L�"��ɮdLD
�����qU2u�E�.1�kT+���󙛎Gb�"1���#Ү�s+���5�am���KP�� ��J��ܢ}`Zh��u����6��Y}(T��C��:����s�P��^��(>S�d�O���s�'�v���̐Qʨ b���l�F�Q�۾O��V�=��k�T>ex�(�M��h$��sW$��4����o�&SHH��hZ���4 M��%s �C^�I�{��ҏ�[o�����}��G�O>��w�v�.|�<����1���^�D�.��oL���� G���:1���e�"�I#&u��C��]0�n�SFB2�|ж�������pz~�sO�}��ZG�R|��դw�*r�B��VZ^N�Ƴ��9���YEq���G�Ej8޲s��u��a�c�:�~�a��	�� (�2���#�ϒċ0�\����/��%$�p�*"�0�dM�h� �*�u+��qz6y��ا�>�ۿ�kY�RAlC	�O�ĿS�<�1�;w�-9�^i��m���T�#��ڴmLy/�	�5��hO��pb�vt6�LtP1\2�e�VH%��۷oK��$������v���[�H����]�LG *s�I�
c�<hT:�9�2Hi��'k���2L��ú�9�+�w�������#�Z�w-��2p��jJΙp��t��VA�Ө�H"� ��H����5�aJL�B��j,
u�E}�d�ԵҞ&l0��1G�*8��[�F� @3 ��N�8�|G��0���Wt��H�E�D������Y�H�� �jZ�<�<I��	:AW�6�`� �ֆ4�S\GG�N�;����z�~��2G�Ǟi�!�3��iL�݌%��@�明�����4cU0�@��&H6��.@=0
a�]Ag%�`�<�����ܩ�O=�T�.q�@
/��?p������p�ȾPUv6�)H���5�Jr�ᦌ��F��g;k֨�#��$�:�q��C;�X����O�
�g6��5 ��i��������H�a���c�iT	�,���QZl���pOa8������Z.t�8��j��V�=X���J�X	��k��	���8q�x�0A��~!K9r^�v���]�����(3�7��MwT&�B��C#����u}�!���E������S�5��u�@ֹ>.����9��w�����p���J��<J�0OB�i��fr��Ț��ߜ�pJ�}<�I�\��o��q[�K�-F��E3��<��_m���h�s6�����3^篽v�j�2�e����A��_`��iz�:�k���5%���J�ׁsy�rxͺ��{���V�1|ǌT�׾��(��
v��"�9Ph�ɩh��a7 ��%S�0LFrŒ�oU���a�B}��#Kk��|&�J��RA:V������H���$1
��v��DvXr)b��r���ߙ���5�{�5g[w޷���:b���^Wޡ5�j�.!#�d���p �+��`�kK�5M�ߤ�����/ȸ��t:M{1:H�m0��K���jP��Y�j �Q����D ��G'TJ-)��Q�=��B�:5�>�^���^��X@�kᴉ��̣� U�b�=�)]/� �*Ǵ	��B4 �A
i��muAB[�9��a�*���m4q	\/�~��a�㙄�������;y��]��^�Ш���fT�q�{���?��藀sVҌ��D�T��|�3��9�a>�u�Z'CV-}���گd[Zi�-�i�{X��އ�漳�� ����q\G��1Vvb��ֳ�q�{��vc8�Rg��8�M�,�fH��a<DĒ�,h7Ơ^�	��6���T�s_��h�yY�|�6�u�p�{i�6��o'�6�(^Daظ��㾤����zB�^�.]���׆D�)��<NK4%m�p�7��AӰfw����g�C.z���uu�_�va�vlxX��Ø������x�F�چ�u^��`"=���G�tZ:0ҽ6 ��k��Օ�ԫ�g�z�ܻ/��:��卬G�&9l� ��d�V�ऒ����k,x��6��%�|�=���H�|����n�X[��藭���O��]C�j3�b� ]�ql��;+������J'D�6�}����]X&��"�z�MA"z�b��=����	4�5,�����_�*�1�鵹b7={]����_�y,\�	ӆ��M�;�Jr��<@�6�R���9�gҏmؼ���L�Wr�H��p���������Qִ��vkI��J�j 2a����U�b.r~r���ԃq��u�$S�0 tlrX+����v���u �x6�<�  ��T�K�j2!Z�`3+�>�`��D���NǺ��c�7���ܚ��ab5�C�����'�R�Y�<z$���4g���[o���ݻ�����}���b����)�$2R���j��Ƅ���2�rf������o2b��m�<��;s�Q�xN�c�̧�5>)�`� �S�`���MƇ���(�%7R����f*���r�}���+� �;an��Ϸ�E�� �=�Κ���ϋ�\�	�c8��:�Im�;H#�z����FZ���s:�:��1PT�ƇC�-$�k���e��7�S_>+�L��~?D��1��1=n���aeT�;��ШeM�c���m���Z�'�d�|�UG_?����/��X��2���R�g}��y�\�T�tk"tj�ǆ��&��P��'W����_��s[	�F	� ������0X��e��UJ��[<��Ik|B����oޛ�m`��/�.(9'/����}�2��*�d��>(;�S�Q�č���ҡT�oǊL>��� `��zS�y��R38Dv*4�2�L��Ġ��B`���&Ɇ�����K�|L}�i�go�!@�iϷf܅2��ۦZ�-s�-��^oY0
����)�o�䇛�-V�Q�����J�,A.B�����[��z�|zL@�T�γ�Ft��^�>3�!~��ԭ�~�Z^ĶXAl��s�w|������z��S"��t�?@�"�6J�6`^�H8�>�ƥ;=��5��!�z�n�z���fE)cWar��)H=I�A�^M��N���o&l:��bir�H5��35�;�w7n�tG����_�N�_�����J� 2&��(1��xZ{��¿yނR���2��@��)�;��М��stڨ�(9�����ԅ9�B!���x�^~�Xr��%�,���`{S�5���/����/�I� ���
�,�oJ��7eǤ�\z-���߾嚇O�W��[Ŕ��5��@���
#ꇯ�j���;�ۗ�,��\LB�/���t\�>Fj3�&SA帇��M}Rb��߿��6��|I�ojmz��:a��fU���2yz^�mH �I؇����?���֧=!�ٰו�������A9G�] :�h՝�y'`��
74�\篡�!�ok�Wι������Vu]�N�x�o�ۗ�3,��()��$��M��M��w�{��M��}e������Ia����e ��L����i]i���S�1��uIc�X.�}mmV	�h���f<�h�����(�\7Ҋ6���R�,��&^`�$��|7��*��!g�L���S����nP�5�q����Y��tR�2��Xw��M�1�A�ڑ�Y�����m�q/������ʹsS���)�W�t�~,�u�>���.��m��!���O_kS�g��{�ܗ�׺��6��(�~���Z<��(l^�"l�0���
��i�(�Ֆ���U���l#�l;��Zp\�$t�u��0�k���- �7 j9����6���o���ȭ:� 
�e�R��u�=����S@�B�����&��|��Oi�Epn����>�R}��r�s�cϰw �����o�V�/��}�:�`���q�Vȃ��q����w������XƂ�,)���u�>s��
~�i]����2&�kb[(P0D��~tM�R}�B׻��Q��Oig�fw��h���!I���{�S?N������_�w�׏�o�vS�t#b˃�_j��H�;px䬐%�Hj8
Q\
��]4�!�����S���q�������dެ[+i���	L��	�Z3g�С�I58g�5��6�k�On0��o��{���C���ʎT�E���I���W���Fe�'H��[۰2�m��P����,{ϵ QC�2a)����r�)�̼� ��6�k�:���X�*�������]R��+3N��lb�R��]�m�<��ܒZ~<��$�5[P.�h"�j�O�8칝鞀���*�rԵQ��<�c7?
���lԶ��H�)��3V#���M��%�}I�[bC A�
7m�����D�s=�jC�������n�IM������2ӳ�൒w�H˦�m��Q	N�m���}Q�2��A]��!%���qx�\ƜТ4��?��\ì�V��~���P�����uӎ��i�C�*0�!�Z���>�@(C}gg��H�<��+�0�H��l[0Mٍ��Qm7�5�tA������f~͖nR)H�������m�,1�Wn�(�F�4Hà��\'�ѓ�$`�kýc��&'X��f�i!��m���������ݻ'��1b�ٳ�=�ρ� �G?��C *x�"�0��_��_H8C1���f���s`
������~2�Os���������@�k^`�:��{0���7e��ߩ�.e�C��3$Ë%ō�flG�L*l� ����>+Ȋ 6<�^��L:a�5�k�Ƶc��z�ڑ;	Z�$D�ܝ�^����mT���Ѕh�i��QתuVF�'d��Դs��f���\��%M�B_*���L��B�w$�0}�{BY�9��2�+R�{����脮���t�u��wi}P�o�s�(���X�ķI�T�e}��z[}�"�ծYD��9_7��{U ߶��T�D����3z�b'D@Rj��q]��.�h�I�{`+s>�>ۖm�~��u�/kBc9�t�61���k�&`O"�^G�^'F��&Ln}���w��r�(4��z}��\(9l�;�h?�R4*�~����4QШ舼dhmu�E � �-Rx��K3vRw�����s�4�A�9F4B��h��#��`lkC����g��7���BX�aMt�M	�H����<C��P��	
��]��!C+���l��6�AمM��L}ʘp��ZC0�� �)F�rȫG���&,�'$��V�;(��X/V�D N)�sݺ�}��pB�kP�I��R�����?�a�D�G��!A7�Mt��cA�k����xU�59`�;!�8.��2 ��uʥj."��~�I������ <���~���L(����}��CÀ��F�(����~�o�3�?�P�;B�B"�9��������yC��yD�.�k��c�{8��>����Am�n�ǉ}g�3��3)O�1��>�����oh��D?M�E"i��Uj�b���d�#���%�6aûovH�u���$������-������{��Cw��7݃�ݯ~�+�����O�"D��k�287ݩ4L/��/��vm����H�Z�� m��1E ��k�o�-�.1�-)�������ow ���x�AX;8���k��˽O�e�ԺL��&5��v~6�Zh���J�k��	Ylʲ���t�w|QɎ]L�����܂�/���I�۸x:���d9DU�)Y¢`��8��.tP�-� ����+%YWϦ䲅m^Wo
��k�Ҥ�϶JgH�{�R�:E8D���(��c DC�`U� ����7�-'=y�����X�8���:����-[$�GfA�YD@#`���M��n"E� ��D��]��\��Y +Q�"��a�+7i$FZ�/���$%Z"�&6�V}�
}VP����!��c�$ٔ ɵ!��a�Z�:�	6�
���5��:[��F�H�������2ך�A�He��Y��ֶ�2�Uc�m��8s���o������tZ���b�L(#���s�x��ٶ�D&�;���)�A����8��7�-q]��/h�PDӑ�d׃R����נ��ԁ-���D�`��d��-a5�(�Ms 2��u�vx�I��f���h�3@3	���?u�=@�]�	EI�ġF߈cZi�lJq	�P�Pq=r����Tpd��'&8<�sV��6ZS�TIF͂c�' n 6H�A9���r�ʬ�i�>��I���V��Y�o��3�0��5�B�R��m�`d�l�I��%-GQ��ƙ�UtN��GN�Xs{7%��_�b�{t�-#���_�$��K��>�cDr�vOa�����b'ء�j-8�	!�T�W8	�p����w���~O� ��8�v����1�U�"�R�UܿD0E�������$����}j���s��yQ8C��`W�a_;�u> ?�Z�19&��_���>,c��������2�ے��K�K�жҍ����K~ $_�DY�'c�I:�Qpw������H#s�����ℶ��)���� ����]��c��=o�1۞M�����C�3	 #`|��}�$
�����ST]|y+�AA��IFē��LL�D:�3�8���P���B<���%i��7u�5}��&_�L���$��{��vvG���H�W��3wv>s3O���4B�l[Ǩ,e�A��H`a���|�&�b+ ��6��)$�~�$m����
��EKF�n�d�))q��0\��]�r7�B��7%n���m��e7��JSz��Q���6����+/UǺsvm���Y`�-�&�o��\�����	6���K�)|7n��i��_
R�o��y���>���1�k �����q�2/t�m'ӂ> ���Pb.щ���@�k �Ї��eS
@���#���}h�O-
���}l����1Ϲw�H�:�`]?��c��)�g�m��q�4X��"h�+&���I�1�X�zoNq.�n �e�4h��
䴝u�ª#�_�_{�3���4�����0od��^�%Z� �,:�sw���˭�\_�+�1���t{������ڜ�v�\��sǒߛ�f���&H�FKw���/�j�s��$5�h��	b�溤�vC���(K <۽ͬ���ɜ�M �2%޷���mcr5�W}f�$���)��P��[`�ؙ�����kpfCV�U��(�NL�D�s@�&�ҝ��@#9�j9� ��ўz�v����4�F��>�5%&j�QC��%:� V��H���������0�8�jOx��~����pw�|����Ã���8��O�?��#��g�KJQI����ж��m�96�-�){NLa���Ƶ���ny^nI��8:�$����l��m 	�r���ډ��E���ؽ$-���^��򅒳�K"h�y���H��IK�?�)� ������ƴ�䨼�_����	oo�6�Y�m�T�"Ψ!�+�Mu;T��P�'�R�s�������]�;o����8���ԯ+��׳0]���!?�	��7�����<����6�1�Ůz6Ќ:	}I:L�> 8��_��_���g&��00���O~"����*��0�"
�(���+�C�x>������ߞ�y��J�L�$�ƍJ�Q�p�3� ��(�����M�����N��#�7d=mkcb��
�N�6dJI��
��~�۝�HTO�>v�'g�?wd�Z�`#�`\фL�����~�1���������s{����m�2�kO���������D��734)棩�!�~s�D-m�ͫI�Qʢ�l �;(�z�h�躐Z(��{�X���JS`o�r����9����u��cD�z�ݓ;���v��J�Ӹ�$��(T�h+�q�&K���:{Rd���ZT"˄���t��457L�����E�H�HF.)�Rl�	T�,�5}�v�N�l+������8~�����D����|׽���QZ��w�kǇQ�(����Ń�bn���S�bu"�7@��O�$�E4}��J�;'���cޙU���r00���pT�|��a�0���7e�����K��c�f�> ���eIGi�>�J�dn�*��mm+�L(�c���E����4���7m59�go��md\��o ����g�ۋ�i~��퇴��I[_$�u�O�dr�GV:���ז>�]c�LA&��3 ������N��;����H[�����5�����?)6Q���q�'�|"��`��O�D���s�ߨń�����ܿ�˿�5����b�G��  [d��C-��dRXF-+`�0&pv��/~! ���i��۷�J}'�)�DI|�k�;�/uW��O&��0 �mȾ�c��B#�E'�V4ŒXЏ�=�UV��i75T��U����!K�uh�u�Z� d�L�^�n���$��*��^E�<�0c�����=]빺�_�x�F��x3.�Ka�ma$c��/7���H)����.T^c�Y���B�
xO��v�U�`�'u�����@�e�6 ��sR0��Uu[�-z�C������ra�F�n�ܜ��,ũm�o�K	��~p[��j)�mI.4�s"7o$Ǔ���L�Jb�����(KMX�}�ߛ}b��� 6�]��|�ܳ�_������'����ﺻw�p�x�߀���_;�w�م��A�Q�l�rO�>w�| �}#�m.Ħ��G���p6Sۧ��&�l��Cb7�"����@nt�M��	V�Y��G�e�i*���#p,��AYC�"�h;{Q�\J���~�1�@�q�q��]o|}��~O�P-C��XC�)d�HL��R�U�O��kM[e%�)�R��Q�0VE ����@�ߣ� A8�A�c�����p�@dXIy#Ќ`R:6F^ن4��g�Yi1
�R&���ԧ�s�oH���_��������ݻwu������dU�{?���}<����i������oЙ��_ ?��i`{pMdPp})�N�l�a"A��Pk�HѼ��sP/���cS���z��gF(l��姦���S�6�5:��]�|ߟ��7�㑮�H|���q�1/s7�����3��9b�c�݋��b�5ɾ�|���˕�C��]^Y��WK-�HM	��㐮�C���su]�x�����$ʦ�{}��n�˯D��2x��V�w�>��G�;���|v�U���|u _`�*~�E�J!�q��M�`�!�7����9b��c[o��~�ɛk��g�J��ms��^�9�6�u �t2���HoJ�K��r�r�č�n��uָ����쬻};zJ����2<����N@�#��]��zfC���������*YU}��$��W�<�ʳgO<�, �㯞�/=q}��al=+���V��&&���ݓF��}#8#���s
�'�j���n���k��p���}�0�q�!kn1\��ƈ?��CE;ۺo6����2�V�c��}8x��,��'�������_�8'�%�O`���6���Mmd���3���m߸v��L�A���;%����5B02�8��5��sh>C:���Լ��TR����8OS�Ȓ:�1\#A�u&Ž8�H)p�_��_�6��x9�>F��`HJ���G	���-@?���Wm�+�4��B��������Q��ӣ�ڡ�ՎO:^�ɲ�G����,@w�*�B.�8���s���mHWef7�2��y3�!j�� ���8�,Wg����a$�X�F?��Zu�eѶ��8aB�]�}z\C�RZ��������n�0����u�����0��g��KTmSUe�.Q�x�h���z�I�r�o�h齩�.�T�f�^dS�p�r�E�;���k�e���c�}�wL�Jϩt��ı
qVy��Z)����G���֫���Z�_�n2Bܩd���,'c�j�5�'*G�����s��=	��XE-
���T�����3��C��[7o��&���}��%i��x0�v p�y
ςM��oh'77�֌D{(uq�c�l;?t����W����}��#hҺ���4ěs`��'}N\Vz�~G%U��l�V˾Th�0:v.�k�!����E���O>��L�ٹC��v�Ka�49M�hՉ�B#��P��~W ӗsJ�D�
�Dc��.l��A�����w�t��*Z��mf� �[F�����n��}���~��_
؆��KC�7��J�)1O�iqݽ{��NH��<�[3�b)��ڈo)�F}��{�'&<``~C���n�����o�>o���_-Z��ڑ$;1��.%����FPT�7��~n�J�Mw�� ����q6����S�����m�`�ua�z�ɘ�H1��I����x.0��6m*W�$IK6�!���6/I�����8׶�=����GQ��:�m3Ȅ��.F�,ʺ�:Lh4��*n���j�6�tI�_���lد^[��\������Ly����mJ�r����:��m��Rn��t>moL�~������J[�������̐���N��Vfn�)������]S�eM�|��d(���2��tN�5́$r�8���>|/� �[���&H�?���wX��+�G|��M�{x�拕l����j�!d���D���I~���Ԉ<�H���-��~HG��h~��q�R�X��QpJ#���s�@�Ώ�<� (�s�L~g
��vچ��L��6)���OYO_�}������$T��C�|W�c!�/�3�0@9�$ː	*�N���`į��c��f�*\����( 0�0��ׯ]�55s�[�Cә�POЙڼ�߱��Ě}D�u=�fA<����O�$�81��������s�N�0P�K3ؔC����X�0�) <m�5؆��������y:�G�Gr��A%p�/M5R�mK�����{}�;߉�a�����BaǺB�F*��A��K['2Hs��5�R���Ztɼ`�9���|&!Z'�J���`���dHߔ��Z!�%��n*1���i�y]�qQ3u�nGe_�� 
m��j+�(f#UE �M?�hZ.+ ��ҕm߉�B򖬣����z:�n�J)��~�í҄~�Lt���"�
�E��b�żn����lx!t�l���������M >�����E�$�H��$�1�kR�t����T��	"�>-�����	����{�M`;}�\�����u�ʴc�M� �Q hG)�5M��"!*M/dG%7�Z�_^��!}?=?s��#�V$~8��y�/��w���	0tYY�S��d�g'"����yM�!�Lb�kf9��QP]����t�f�Bv��M����@��!]v+6������c�';c�q�kq�l���w9�@����}��osqNCf�]�^��_�n����8���=�9�t�Y8����	O�D!i��D���F�4�8��`�`��>���f�e3v�έ�&�����m���s��}��˶��b���p1$[x��q������זFkP&QYZl�m4�]��s?ꌧ�hRժv��\��"�����ޡv'����Ls>�g�8�v_��uY�\�!HY��8�ɭ��hQ9.0V�5�g"���[ݻ�t�3�0ch��`����w�a��2��]��+4�?w�P��k��BD�Bv�-�v:��4��� ��)	F��"�=M.3@�G@n�$@Kh�t_ ����QG���x���[o�%������^Ö����!@�:��������2P���O3�N�- �a�J&s"h��"Q�M�di>�
u�p!��Ц��%-Uՙ��tM����Ò�$��d�w�{nQ�Y��{ә� �!Mv$i�����t�U�|�l�JC8�1�p.]o)	���_4��7��a+�'�y��E^'�t�/��E{�s�!��X轄��z�Zľ�!?��im�#��5}HaGG<�~�TR��
kڜ�ƚ��V�A�t�[��Ŋ����)\��Qć.2�C�k5�M�^���	~�=��ޟ��w�¼��ì�gT2&���W?�e�5���ܪрaA�*m.��N�f��jaҬ�Ϛǐ �v�JiIXm��1͕`�4Y/+;X�L,9鏝,��M@?�7�m?[gJ\@H�ݞ%��iD���dG�jDl�FwQH ��� ƕ s1�1��=-Md����8�� 'R�:b!F���5��_8�1�J%	9[������W 
�e��+��a�汚/�{b��������}�=|(��p�k��t�����߽�~���܃�?s_~q_T�;����w�8{�)�k��&�HT����ҶO`�5o{+���R�M�_��Mp{����a�]�����J���-5���g�Ǯ�55�7�\V�����fmXs���,�޳� ��~[Kd�zmozצ��w�Jִ[��!_�1S��ӐD#<�S�r�ϞE@j� H�EB�A�y0�clq���äMi�w ���,��I����$��O�6�>Yb��	,QRzg������\�i��JqikOZC-(i2�b�6�~�q=1�F�&�i�G�7}�I�o�)3���u�p�[S6���c��l�g�?#��=%n��VQ�T��T��O��S0�K�fb�V���k��m��ZD�B���8���v�v�D#Zf
����n�������98(����\��DSb"��!=lz�����a��`�+�j|/���u�p���|w��r�<��>a�μ+��4�f�i���hb�fΘѲ,��F2<.ۊ�n_GI%�� {,�)^0/��]�~x�E��?/��|61W]X9��x�"��0�)I���}vS�b���w��H� �HzQ�dH$M �#%Ԓ�UT�F%^�yK�:bOGXr��^E��Vb�f(��}��<�q|$q硲D��G��g����q��W�'�2��s��H���k�n<�{�������_�c��񠏮Kԁ�~s=�����Mwt�;:�����;=y�
թ��gb3��7u�sD��]�#��U�λ�L�E�LBB�t�l�f�.i«���l���1�6���$t�;�qXOot���KF��*�e��z �y�g����J��E�NM&� �s�$��QZ�{i�b�}��N��]4!h�LKW�6�� %@ڿx�L��s�5��22*dVxm��I[t�v���������
<p�WY����[@�2"����O4�>N���>���.�sn����~�xͺ��>��Ta�H�͉f�=yq&��p<ݗ�O-�S̗	ړq��:�t�ֱD�Ǖ��<{�{���{�����J�'gn1�VM��\��e�.���@U~��G;���_����u�$}�\ɢ�b�x}YESr+�4ɽ�z����>�m�"����m���3F6.�S�g3ᶝɯ�X��c�da���{�����ɹ����Mv�ޤS�G
�P�]g2�o;P�$՛6�����~37x���!I�M\_��*�Y��\S�k70jH�Ô݌l|n�@��/:瘺q��T5W;�hMYm�j�)��H�X�1ȶ׶�1F�9HCJc��2��w��-��k7�[w�]D�X,E��'��Ï>q3�/��6�)E2��RBr���~W6���3��;<p�}����w왃����)�$��8I%le�?�>��#�8?q7�x@(ɡ`�/>G��S�nKY��n��~�=+h�4�&�d����[�g`��L�tE����%��Ϧ��d���s�3Z�~_WI�p�����L�s}z�ˬ����]���	�5R��z��\��jUX��9���(' ڧ�/	�����Ӊ��۷n�1j������jx����N۹!]��V��V�l����X�h��������o�g5����}�l+�g}��t�e{h�c�g��m��R�㜷93$�I�c�W|�N��>lE�j��v�>`�;���c��=��}FD��hM�� T������/��C�3_�"H�ar�|�x�o4��[�6�Z�D��������+���o��.�O%̫4��5w��-���������.<~Ӧ��8�����yL��f��)=�;�����Ӓb��-ٿ��}}z�ْ����u�®y�����}10G��� Ht����W�BӶ��m�a�����ܶ.bJeA��D�%��Ӂ�G�w����DھǺ�o+��6嚷՗�]���,�,'�%�6
%MT�Z�NF���vcJۼ��:��Y�K�4Nb��bԩ���ΰ��^>���^�|���w�9 �����޷�7<��������cq8������!�w�&����Ϟ>u?��O�{����s���w|�g��/>v?���H����C����r?��?q�Yp���/~������~K���ﹻ�߼��gf�b�p�׎�G�=|ꚺ�.L�R��Jc�s��cׅ �}�۾�������Mw��Վ���מ"}7����zO^�LG/�oO�3d�71��v��zꎧY?e=��:m��l<���K�"������#�}���A�b��`xi���� o,� G��d�:24�t�~.�����I�P'@*��4��������T�Мł}~	��û�9������J�SK�)��
�=oMx8NV�h�",m$��_- �{���o;����'�#�F���_����	���O�a4�n!�J�W��"6�k`�	6�~���-��}��y�Kw�����tǝ�=Qr���;��Q��
 ��vud^���@�&?�u��U�,QH�9g�Άߵ�֎���B]�w�v��� >��������'l[�f᷂��7��v�n�u�$��N��z��$����}+�z܌_�����69�U���Q8R��L�&�<�g� ��\z��˔��o&��\}W� ��ۊ�uR�mL�&��#���<�9Y�~�Ɍ�B切��Dt�Ѥ���\�v�n\jnz�}��]��l�W�?�f�b�x���{b{|�P�߰U�bĹ[�n�O��RѦ8��~�B%����s���T��ː�C�����o~�+w���}Z�w�s0/���p����/~���O>r����ݻ�C*B���g'��7������h(�\J��a�k;�i0ꭋYiUZ����?�N(wE:~b�x�R�%����Eې����{�?}��]�G�x�v
#DqW�b�'sF$�u���o�ȴ��ym�u	�&�$� ^׮]�k�<�7��8�}�FƲN�9Z��+G�r�'w���X'�a�BG��h���KjJ����������Q:����,Ɯ�s�,\�(?�W������u�ж��LYF#�W��cKY���Mc��i5 ���k_%�`1!mǻ��RC!uЯɅ�M��������w1v�q����s������G���?��{���w/<���~�.�<??Ӝ����֋~�q�뽸v�aY&}��o��3�w}a�:̴�f�>�}޿�դ�IP�k{��6�M��XM��,=z�ъ���pY7m�z�k4��H�ٜ�6�������P��f�9.�M�9���ޛ�)��I҉r�	��=���mJ�m[t�y�����U�H��sc�ԋ���H`�l{�E�F�Y�0ֵ�����[��v&a��d�Za��ym��Y����h@꿻����^<��f6-%V���	�gZ�B;8�"J"�<y�Lb
�����f�����BLu� ���}�>��A4-@��Z/N܍���w�'�V��?�Ll+��y��1���o��K�"UB�6�*Ԩ+]GuR����!(㼊tE�~�И��;m�JnM��^��8lG)WX�!mʵ�ϳ��H�@��HG����z	��k�%���������:�kT3�m-��O�fle�C#��Ȝy�ڝk �6�zR:vZ:���9b��RG�t�l�O�LZ�o�uꧏNj����t��+�	KK����0�`vPǝ!"F����qJ�t���#QP^�p��/��N������c��w���54�}����<�cf�V�w����} 㦩b�R�4��6�Xva%c]��ס�a'�+h^St�X���l.�߯���~����?����;��> �(8�.��~HT0V��.�&��2~*��n��zǴ�����1�	(�	�}�ӗq�&� ���w�I�6c"�1d4��	���RO[��6�∋B{)(p.�i����K��b1�^����R�ǔ�����;.6LZ{Lv�K�K(,aL���s%�@�ݴs�lc�ҎM%}�o���5�I�O4y�*M�X� �eJ�P���S5�:Ŏv����$]�Cl\-ǀ8�f1#�l�f����b�G�zz��ڳ�]2����'����v��L�k#M�S��g<.κ�ը��Q7��@�Ap�;i�t��`@�%_��_�5�/B�͖�R�p�h�H+���o��EC��c�sm{5Iy6RI"5�q��y���vJn-�I[���ۊ�{Q�_��#�4�;ޗ&v�M[/)�xٶ�����к6�م�SI`V{�abQ �J�w��c��u��$�0aHE]31�i����3<#�+Gs617.(`��D�Raj�f���f0~P@E@���2�u���gH�������?
 7��Eh������{-���q�+�����}�B���矻��ۿ�~fd<�@$!ԇ��������v�Ґ�b_��R`i1��5��j@P�1D�^"��f���$��9K!����H7{��N؎  �L��`�TJ���^�%��_���������.̾yzq*�
5���>�&���~IFa�o�q����
��e���ڣ�^%р�0�������_2>���s-7wY����4
�x��?-�Iq��;��i�vQ{���,�W�bfL%q|���9�}���;����n��� 0�l�f$1��&�%�(��^׽O<["b����ؿs���9����,�g�v���l[/�Ȥ��GjObh�]4��ċҢ�[P.&nA�α��	��d�������vv�y#�VMԡ�Y��+6Zث7��ԉ	�RDqo��H��إ<�l\�) �~���-�p�_�
�uh��}��{��$�A$�e�Y/氩�f��OB8��8�J��j���X7��H�K�X��Vr��(C��7u3v_=9q7^��]���s�7����g'/��b�J��F\�w6�)Q�M�fpô�׌Jz�gGƩ�4+u0��c��W�����Z���K�#T��vÝ��jR���t�k���L��u Bl�]@�fU�6p��>��4��V�T�������Xwz�0��v�����hJ�:`H��>-  h�g�@��5�f���A��*]Wgj��,[$ *d�*�/u�f��b q|�>� HH~iS�����R�-7ik�aۛ�x-ǋ�t�,�o�Gq|ӑ� �k�C��0(�Sz��}u���"uGΈ��G��@�������ےu�e��C��馗x	L�>�: ����;���I�xܾ{
���+���A*x�@��6����X��~����7aDʎ�`.Bs�y�k���]���Eف/��N�ψs�<��ܲ^��ږ���}��w(mB�.h�F�8��gg"l���É �o~��J���p��eв]R�����tM������\"j&��J���SY
��m�8�eT�B@H
9��!>��ubUB&�!Wt�}ԜX,Wў�m��&�S"�f�d�i��iP�O-F,�o��z5m�_�k���0�w��� ��	_�+D�	��jr��]����m
"r�m�z�����|nQ��w��׏G~��1 ��M�k+?�IŪ�ҒίѨ[�(��d�gǔp��TW �Blk�[#M�����*)�5;� H��`��4z-���񧟹����������޴I�#9�̬�t7�� Hΐskd��a2�f������ߦ�kk��һ��F�j.��gH� q��uWfl<�ᑞQY��z���FU�qx<����=qD�C.��Q�e�؃�@<u�q!�7#�s\tEsf3q�@Q*f_u��� Xyx9\�g�����7��b,�}7�/_�[���[ˇ(Fne,y_9g*&�+�Ⱥ5��Ǻ���W���5kHD��C��U�U�}�9�&��C˦fY�j�¬��2^�}�t��ĵF����l��\u.+�U�s^��+=3y�k_j}/+b�KVg�n�֪��[yi
��[_�M��,�
��m�	��b�뭢 E�/��w M l ��l9�9���s�� ���E�u�+84T3�h6���6ꢓ*lm�WV9J���]�?��O��$nۯ��S�P����j����3[�h�W�XR��!.�r�
����A�s��Nghv��ߨ�_w�@:�ٚĊ��%�7׋�W.8���U+��o(�Ѧt_u��m�~Z@��|:^�o�KR��*X�����Ԯ�鏶C�DJ��\О��e��Ƹ��wX�iM����e�T���z�SCJ�op���u{R�&�����]x�N�~��3���U��MYx����T��{���7�2���tҷ�5}�����*ݘ�)p�ܶ��4��Ӎ4�$b.�_]�^�:���V6�D�6\g�\f��z���\�7�y��0����G3Z�+� ������s:�8g��n��3_Hi��|��堢.����i������*����&Ѷ�hJϟq���mNo��;�.P��s:�
���Zq�!�� �F3')�Vۣ�����k�M5���
�r
H˲���u���|N͹��!��s����,;R� Hs��!�Ti39�"��֌ZU����$���ZV*���k �\�f3�Ȃ`�>���Z]�Q����]����7l��>�ބ������v�Ή��|U5e��i�8��-O��}�V-���2O�о��mV�c-���zc3�a>i�%��9���{��oU������fB�������m{�T�ٚ��*C��.�i��g�s���Ad�u{}P]��懁'�.O��3����{�y7����J�ͣ`��pwq�y��a��?PJP�Z���VOb����b�"s�̰J�؟1뉝�|��9Y	�* ^|�k�I�n���r��n�q��Zf=��˹�z�����|Ԟ��P\�y�w*�e��d^��b�F�C躷 +(��7�
y�G�K�OK8O��2�6b�q�/����}סc�I!��
1Z"��LnB�3��9�^���n��mU;W]ߦ��=w�>J�L����6��N�u�_���n�g�[��&eŭ�L�l�[���j�jbM����E�����`^�C!�*<�
�0�x^̦��n;`��|g!|'��t"��s�@}����]0��6
&������?yP?2�X���O��Ş䮆���g4V�<=�o��B0lo���B �J)Z���1��~��k,̟<{NϞ?es9��FH�T�}%[��Cc6=�琂�҄��m��?���v ����Xo-
j�-~ճ���Ǧ9�1<u�]�XZ�L��Uώ�)Ld3��Yۣ�報|c�j[���\PX�&����h�����<�;O��~lھ�~��rϲ��!�L;���&g-���h`��V�b����-���Y�BA�f�����{J���}������?��7�\f ��z�-����ֶZ7;5�n4�g�,>\i<x��E6���~��~���y������V!��p�Y�1�m�='�uk��Q��:&��)mЅB��3���Ʉ&�(�ȋX�'�����nF�9c�8CjJ����w;�\+�k�Q���ʹ��ه����-o͹%\ε�A�:�{�X���,T��s�VQH��Yf�i�lj�5W�Ҩ�D��K����/��<�h������y� �t{3P�����>NW
��:l�uV#n[��&o67m��m�i{���6��}m�l`U���m�D����ǫ*iv�ҍU�R n�`�D}�X�8lօ3�S^X�6\eՉz͛Ҭ⪫8,x0GV���gXÜ��cp���(�_�ۑ4�.�/!� �K��	���3N�ґ�O��j:�r6!7�r�n��Yh�Z������魯��,��Ǐ��]"`����hk{�^�u���i<���Ő&���C�@
�������x����^P����]��I� YE���3�=f~a�{�X���z|�C�ͽ7��7c��Y�rO�l�F�
җ�A5��&���X���m�k,�f�жc��$����$�G��3�2gt�i�[�A���U�F��I_�g�H�9�*�@�{D@ܬ�,&��g��`,kiNn�(y��SA�*��E��%�=�?�w���N[�U|7����)g��|��i�Ҙ.�Ɓ�4�4ּ0�c��������?�3�� �O��O9�U��+�����*
�5<������>��S����&�W�ɛy�m�h�*Aa���/��M�N۾o��&���2j��~}�Zqk�[<���B�Ľ��n;1�+��/�X��/�e��Ɉ-�|N�v��Y���b4g������19���ӹ����B�g��s�
Ě���y��ےXó ������ծl�2�f�K�;���40Q�`�b�@\5\�T6����a��t,�����f�fF������X5eE立m#�x�� 5�!�Z�K��Fv��\w���_� �궍�����x�spXJ���pX��_ �mOa���j������U�n� U@Ys�
ݘ�qK7S�7�&�����R��&����|N�L�{,re���� �g4�x�;�j���b�Xn0r~G��~��3���s't���ΙɅ�ԃ���3{��֣KZ�߯\pN�k�s�M@���ݝ>\�s����./z�:��X/z������g2��� ��t���^.Gtzt�ۀʁ���Un>`�!�`q��nI�-xY�<h�{����w,<��)���w�$�s4]��������A��S��*�
��z�	��³����ĴQ�J�W���5��[����X�B�� ֢�׮ʈU�N��<V&[v�+�m�}o���m >����[5&z-�C�q�^��u�4%/�W�����k�&z��ʂe�vd����*L�m8W�FZ`S+z�������L�*P�"j�Q�� =��m{��٪��*8v����ޑ�)��Yg�1�b��E����ޒ�yXɸSpY�����mpL��}���T�n,��l@�y𺕋�Z�	A���*;�e|/+}S8_�]M����ʽ6��� G�5�k�Fm��:�y��� *2����9 ��x����ҿ&�P��1ɖ��g�q,�p�⒘��%�#�N�9�j�Ўa�턌���s��������1�9���[�n�ܗ��盗Y<��w���$�� xz�U߷��n\��u����6��0H�IM�)��z��I���{\u�=��� W*��{�zf*�q�����mfj۶�E��롛��xf%��®6t�K�NQ�� <����q ��g4�< �y,+A/��)d��5%��4�,�%s0O��H��ym�.{��5�_��ۄ�^A��G����g0"~�Ay��.Ύ�w�5e�މ��BZ�2d��7��Oh8:c�K��y�...�_�Ib;��<��Zz�~�d��Cf��K���jZ���W;^��Ͼ���U���օ+e�6��d�5�zS���\/����������j`su��=�S�f��#;�P�1p� �j�Uٴ�&���33�5ڿ�нcUX+o��~Mmu��6�+Z�h��n�k�|�+l&�ҭ�w�����n=϶���M
��¢̲*��(�Z)�o�U��m �ZB���nE�`�սF+�*��@=U5ݥ=W?��_�lᔺ)�>�DN��e�>h��:P�*Jm�⪽L�Y�2\�U�l�4�g^[\x~�_���c��SgB�F�~��k ���Iȥh��ո�7�*�v,j�j�?��\iXλ;���i�������%� u&i���w�U�+�[�pP�pЗ��?h���(3Q���6GX�mYW�PHX����X�{���AyV��A���j����NP
kA��3w���bs��t��=�ʅFo���l �PMA�f-����h�L72����Q��IA���Y��t��Z�x�	����9���h��Ҿ��bo
J�jSC�[R��s4��e��>�B^�����}�gw�f��=��>Xo���y1h픅MLs({@>��x:���_���X�]M��gK]�C�>ݻ��޻���GǼf�g ~�X9���.�8�NE5�ˣ�&%\%��U��I;P��]`2���e�;[}�M��?��R�*g,Vp���п섮������k795X��x,=��3���?��<(��I�G�`�F����<~.<
nJ6�+ ���fb^l9��R_��s��13���%��̗Xت���Ɗ��ir[��A��lS�4�J��*"`�m�6���Zaic�O�	�Qs�;h�kp�QW/�.�r@�&
^*���3g+��u�\s����˾ Ñ�d:������Wr;�k˅�X�=
���&Pے�cھ��Z�c���V9$����^���`!��d)��n*VQнF�qE���f�������	 τB���Uy���1�����T����p�Ax������+����%�m�{�=�*,�a�s�}=�FE�c3���z�X5H7W�'��9�?NpiA�Ҩ4�h�kr�;�?*z~�-zL�h��y�(憛%�� ��L�?X��L�4�]\��~N\;n���T.D.�8�M�Z'��xI!��B[��qQ:���ױ�cQ�����o��c��~������\���U!P]�?{5��������5`�����=��_C�͝��!	��Z銢W+P�e,�E�a��>c 2�h}�/U��P��R�	9���8isA�*�QY� ��x�n���xL"��U\r=��.07	�j��]��6;F�Z�P}�@�6mlqN2,`"��V�2X���0Yt��:�fŅ+���2ۄv�2.� q����k�[k�ڿq2�96Y�����C|�$�f�(xq�����H�%�������7d�Y��Fp֖_�g~#�{��v�F'8޸N�|�r�v��t�,'0�������3�.���������n�ypi,�s�EW�u0Ν��3NF�_�A?������6���q�T_�`�G�'�|B������|N49������É�C��`��d��j��=�����}��)}\r^`�L���ؕ\�fL����������?���~��D�;�tz���τ�φ^��Q���,>�Ùh���P�;u� ����Eɥ�9;H@l&V
v��D�\�k)�w*�wS�8�G�`�Ed+������j>�WBe8�u��J�_ *96�h2fH�{a�P�.I�1�Y[�j�\*����uczS�����}��<�3�k�����uM���A�dr��b���
��̯+X{�\Ue�`�Yv��^�%c�A�W�EV���s~f�eN�S5ec�k���_Gh�ti.��z��w�`���9�w"���֮w|Ry`���>�K�z@&%v��]��~�������OD���gk@���Yq/x���k����c�r���=l�uW0\[cԟ^�����wT�ZЫ�V�O���f�����a�7�Y���@j?��|�E���4�����h�>����'��w��]���G��n�x)�V�j�a�S��Ĺ�1?����_��_�����g ϖ>�u��{)9�������UѲ��*3���h��J��U�����q0����1�/��g�*8ފ+g"���K
 ��G]���ȳ�
T8���x�wG��{�S���N��2b�5Rwv_�6�/�^<����ْ3�A�y�>'��s�k}J��z4_d�Pu\K��������wd���TM��LMl�*�������4�������x�{!�!������V�~���$�ᬶXR�A�����k��X㺮~��
�a7��"\b�����.�Cv&ART���Z\X>t�1�G^wU!��an-X���b1��;1i����2�a츝/��C8/l�FU�@&*���+��ڴ==좶�[5�Nǵ.̫�Ʀ��%����)���8����VW�X��9x��h�&��g��������Lo�b0�3l�Yr��(K��;�x8�+Ng��[RP�����و�{;,�>|��������?D�RRB�af����p��WJ�0\���|2��'�h��{].�s��uz��[���u��/�-w߹G���7X8��3.m>���^�Pf[��gĊ`���ҿy��t�o��6��^���Bi@�o�������u*�����'��~AϞ�M�Y�z�p��~�f�ϸI�>�y��Z霣�=r8�i��Z��r_�SA�~�ɤ䵣(��ۘ��M�Ϊ���Y��D������!�"�6l�]�ו�:�u�:�'I06���@le�q��������E{�<�M
��G؄��"��c�B� eϦ�P)�/�:�MV ���kH���+6O��w1�ү�U�_�a����*{	[�st���)[b�d宊�
L�_K�ܠHv*q}�Ռ�"|�1��=@�e/�%e<�u��{
f����-�Qt���B*זҦ�R�;�������%:.�w�ԧ�R jY}��?*/����8�����Q��1x_��?����������-��Ֆ �iCQQK��5X}�Okh����W��V(��-,�.k�o��o�*v��ۉ�U��� ,�/��~ p��Z8�0Zi�HF8q1���̻X<q`��W2;����]�2�s��{�O�g���$`��R��F7�e�]rJV`:�N1(mD\&4�w3�jqXs��b:V�-h'�a�={qĊ(�@Yw���`^3��.��5��cYn��su�?8�y�DݱW����
����� �v���L��	��r�}��39��'�Bܚ�`AȂ�>�G!^a�tA�Щ_Dlu;��QR��6OҶ��c���S��@ `�u������j��B��N�IA���u2'�w(N�y* ��R0Y��6Н�����L{�Eڳ�H��D���>V�v�Q��݊<��;���I�<� �'���A  ���p|��g����o���Xly�]�g�B�i��.*h@M3f�aʻs�&���}�7���S:9;�s�/�p
R��J A��}O�����3�+P*��C�E��D�p��B�
�A��wFj8TE_Nؔ}trB'^��Pw���9���`����W>�£d��f!�L�B�U�:���U� ��W���.��r�I��ss-�c2�Po�fn��u�R�pww���F~��)[k��`z�V����z�{{�92
�����3\��M���]���{{�"e���r�l��f��3M�[y���j�oPx��=�E�/����K;�қ/Kg��ϼ2c���Wkr,����ܨ�,�7��#�G����`��S?����Ps�* .F(jVu�2܄0�ܭs��P�����r�n���m�
�yf׏�7
��Y�
Va�Pt,�{�0�u��@1S���4�
^�Bi����ZyTd�Zn�P(�y"�%��<��<���j(A����oӵ�o�[gm�Y72Q���)�{��'����jN�2,8'��J�d1#���jCz��XM�@����2 ��OŠ�İ#{�	+س��}��蝷��ώ�����TRC���>�l`�A��	�0��m�V�]�=��nY��;gꨤ��7�%��ߪt ��_��_0���Ӈy��g2���ken`,���H�� ˌ��?�ZXy���2�e&�2T�P$ �*fR��>�P��Q���&�83�,����V�z�Q�wz��J�I(d\g�[�/r���PC�����Ĺk��-�.42?�_�i^�2n�m��U��U�Ƕ��"�xzͪv�c�ׁ���V@�-sb�����=�2?��Z����ۮK�KY�UǪCY�u��wˆ(����&/w���dO��`V��q������L�o�������N���O�s:=:���͕U��*g|Cq���f(M�bwu���	?��:O=x{�
|$� �!�;]��G�F�h�Mn?01o sv��tz���ؿ�G�v�1M<����tt|��aQy����K�}�[l�|qr��ǾM^����8� ૬�.u8Xg9�Rz��;>?3�8�?�[���z�&J��	U�A�����+)~��%G�â�3�ǽ����L;~���ɦt�c@��A�� �$��p����|���ǵC�����((ry��b���q���k|ù����Wb�>d,�%&�y|�w�d<������O��Y�?��}T�y*U� ���Ʃ ���:�ݢ ��o�ńS�.�f2�t���B@��*w��8�Պ�l�u��:È�t�ā~n�5e�e�4�4�g��j<nT��{(�U+U64{�Xv
Syz�>�����]�}�M�Zq����/��k�5�T�mToc�l
O�j- �&ݫW�^��잢>�:n�����D��e���}xNϏ#r��AN�{������%�ߺ����9g�w]�H=|1���}�[ߤ�~�=����.8�έ[��9��9m��@"a-Cfh��R��>�g[�uǦr6=�ZL��25�f��7���߿�{zv������s��mR�*�`�t��<&2�&��<�q�-�����s��Z���s	�^�B?���z���(S���ܛxf׫���������w�������=�ϕ�l;�
��N�k�(<$������x���q�W�|�,�t���G
��`���
N+T����\��^Ϸ?��]F���}U�ڞ�N���6:ڮM��U�W�F,I�k (0|�\=��jA���4lʈ0���%>�!`6c����>��_���K�ͯ?�
C����߸�}��%L:F��"(�,v;`r���+{���G����9�~��h�)@>*���n4���O������EO���`4�`��W���\�s3��U�}�� 
���)=qD}�}��1?��5�B���}}z�σyQ�Eh@ �)�#G���u��yȱ n)+�G�n5��%ڨ��>�)��La�[�ZW�,��Y�2 �ݼ�"h��/��'����d� h�LƤ~�:�q���"c���V|��;�D�PJ)1�Mx>_Ġn	��f����^ �H�pyy���P2 ��o�\�MU��=�I���r��B�Ȧ�Ԛ�S`�"n���}?_��G7��\F��1��G�w=~�����c��tw ���;ʾ�AEct��w��;��g��LOI�T���, �@s�?�
��ZWϱ`�ᘉ_0�E��g8�m�i�p������>����8�`�*6��c@I��TR��!X�?~@���� A��'�E��~��k� $U��m��89h�_d|�y�C�r%���G�V�r������!������y	PLN�Ϋ0��a����߹ Dޟ�z�� P���M?����7��}?�3z�����G��0~7�����=���ag�k{ Q�0��^���"	f��y�·�v�G;���Ι���G_YI��i̙;��֕�d$^ y1�J�sNҀ�z~&��Ӌ�`�����1��U�*v!�9%iP�����8A�\8����lm���n{�����\��.�Q��V��l�B�r=�6co�����ݻ�Koݿ-�<��qU�D����,������<��١!�y���Gc �/��ȑ�s�)��˥��6�ژ�8jY����u��/M7 ��L|�{�H-�3�#{�n��v�Dz�t�Y����X�F�h����]��RW�LΏ���:X��-0: 8�~�k[�&�ty`����������߿�E5�����L�3(�����<�#*�$�,|˱�	=?=�O>��l:��JDׯ &��$G%���cz��a�X�2Om��ge�!l8�%��u���O>��<��g���Cz��3g���%&vdYy���倐�����TܖEͮ�*����.mfo�7���,+j���~Vϻ�=6�Cms>2�Y!�L����z�� �z޵���ʃ��a&�Gs�㥊N����!�̺��{������E(<LU*;j2�^Ӹ6D�~��KU��3X6p�ٽ&��X��s�_�g={v��&/L��n:�0K���'e��k������5��ξ�4�a_c�����)��^�����	`"�< ,���l��6�� 7uUA{U��}��
�3P��w�ۂnƭ��s��{h1�޽K��� .W?�������-�	�� +_XRP�	�����>��/�qJ�����-�я~D���o�o��o����︿p�h��Z�+�.%
b��F��A���O���ן����I\M?2�:_q=W�&��A�o]]�����1$�}��۵����oUA�r�M)U�,���T�=��B�um�\h��8�k���r.c
�%9�R�8�����=z�����G7����ǿ�_�����-.0���үm(�Hl��݊
������ڴY��68���*���.�
Z嚁��N�=�s`s	8F-��7o�Yp�E��|��أ�A=��Ɔh�L�^���qf�P��2�t��E�������ӣ-��)�ĉ�5�.^��{�x]�sV�q=l����؃Usljd��� ˪�
���FN����`jn��׿:������i�mr�	PێT{����E�ߩb ��)l�m�W2���._[0���nRsw�5Ñ�U�jcI�����
�o��
dT0���*$
�8�H(l��
7fj1��h*�嶙x 0��_�?��/�_������Kd+��_�N�j����H~Wf,9M��G|E=������L����ևّ�F^���	a��4�Q̴Z�xH�]ga�T<�|�W�e0��=~�.�/���r<��&�rf�|���m�C�#䯯���;�
�b2|:_�Z�
,G��L��@wj�X�\��;��U�:梙ǹf|!g����M�����K�҆T����nk�޹�����=^x�rH�|B�"b���)+H�ɜ�9b9�̘�����6�O�CA���2k�J�;R`~���^���?�~�l$���+�`�����G���n�JTe� 7ˢ{��8�~׎Kd�7��]b�*o�|�+&�ݽ�� V�&ke׫J�� @���DAvT%����oV�5�?֓��4�,8��)���[@hp*[��S�%���]`A5ӏ>�(��aC��| � x��o|�A�*���R�	�V(��i��Ksk��I���:�����J�4��
�pP�:��N!����ù�NvmY�6r��ʥy��Az%$�"aqB�8���>���\���P�xL����rV�Iq��
�������֛�<PߡgO��~@/�>�{ń�������M^���@�9��D٩$v(3��4(�y��,};ؗ\�Y��5��Zf
�i�}��U8/+�S���B���IX90�aa���X 8�|�Ӛn7\�8 ��e������q�ۍ)��B��v�k	d�W�������T��!�
�L�������5 �N�ʃ̥< �+��2��� e��AP����W-=ܗ�Ue(�����t/e����U������}�=US�=v!�-ݴ������w�|�x���݌�곴�z�ׯ�O+�d4�ڲi�l���~�!�G���΁���^���j��@� Q#}&N�.�Ï>���������c����+�#��6����E��$KI�5�%*ȞP�F}�j����P.��>��B�ӡ_'sKX7شNώ�� z�ƛ5�!�1Ѝ� ���p��� ��8׉��������V�5'�����G��� *�٠ګ��e�����뿿*I���cĦц�^Ug�� ��@�l�������c#�?�g��{)�R�}�@	sc� -w��}��#�Ժn���m�Y\i�VW�⇍��v �Ϲy�:�P���l4���gJ^�Q�������o`neY7 ���ɩ܊؎求��q��Aɤ������9*�; �7�����gb��6 )؊�M�Ay��}Ҹ ��~&zV���D��Z>5��^g�~��H���Ӕ��L����U�e����fP,)
P�^+�W9�m��ӡ�M}�!GaI�V���_2 �K�͂0x�∯�;�-Y}f���3�~()�Fua����i��(��9v��`-^��j��;;F�7�&��Sո�X��B*�R��Q��\��Y�AQɀE���M���k����O~G�=�;]?�F��.=��@N�6X{�B��e>R#j߫UO��sJ�Ԃu�T��H�����\O:�,���]Tu,戦x�g ��J̯��Ӹ_)�4��2����p���c޽{'ĚH�,��$ר)��%����J��汽lIe���:qN
,���-y��,�m�ǎ�mݞX���s9�hCV�lz�U�bs�o��R}����տWުm;�&�n4��J��i��-�^�"�
�j[�w�Y�X�n�}���n �����ۮ��� ��z+�؂UmЯ��v��ϱ�2֏4�#�h⹩\g� �j�ρ�1��2dT��3V����~��_�����IO�����jEm���")�ݙ����J�A���:�x.�� `9��\�6�I��)�B �U247T -�=��}YwrP:�B,�͚7�9�KΦF>�]� 7/ܡ�gy��Ae�>o�s�:6.���0`M7x0���l���o����֘�]7'���))3���EQo�6��t�����V����@��1 �̄�A��@9�8 �� 0��)�<������ސ��ò3+��_#b�v �ݸN$��qI	2����[�����:�	l�3)d2�)����(�y�.*��4��<��P<��ςզ���Qܦ��c�?�D<S�u�f,\q㨤v6��[�o���vh��pM���w�o�MN����1�=�<<<��y��BQ2v��D �~�M?ȗ~�dE���E,����ZH�����?��2� Ē=�b^a��(c��W`�\7���y���{h��k�q���3� �Vh�������Н�^g�Ɨ��u�بJ	VF5L�����{3ک������E���k.{����~���%Iװ���{[1U��^���{��?d����f�(A��H,l�M�|Lʘ2���R������-���m�s����y�'�6����k�y�{��d,!��y�����2r��w���߁{����C��F�,W���z�=R|�5�QS!m��jeG�B��r�#�BU�V��r�5X΁�ϱMh6�qf6�o�"�	.����E���?�!�y���׿����:׎`�{)�.��~��@ �~�<ƽO�|E��t>��"qKpL������QV#� �*먫����I�_�Wߖ��'Sz�+p��C�Ȃ�V���is�\fu7e��X��eɳ҉���X����M����u���M�JIh;���d&���I�U|����Ŭ�L��#��M�
p�-3�����sy��]�w׃�)��_���(���?��_��^�<�No��8�E�t�^vÉ��$e%X'�0�|�省��/���D�сc=�Tp��)���ٜ���0M<���Is�a���CS�Yx����r���MK�\d��Ki��o}�v���h��A��]/|���B|�!8����(�ng��x5 ���e����G_��侭����-$S
VIbUp08�M���W��Q��a��චl�2��J����Fva�̼�KR�U1+
��cz�%`c����N���1c|ȱI��.3�v��"@���L�X)?� @%�x΄�>P�;8U�E]���'� 1-HX�Jd�A����m���.�dr��\n�w`an��CzOd��\m���:�8+c�O��!V��S;��[b������m#�p��b8������χ�@�� `���?����<���@�B��X��k1=�e�\���������f�����)�[=0�?<�C~�Hh6!>��.+��:.���M�g	"��vll0��1KD��_팼~/n^)�sfx9� E%C5Z��{`��kG�I� z�3��ы�4���ޝ��k��
����G4.�z��jn�D���;կ�c�i���ݲE��?�:��5�@�E�/���N�:��ź�^\M*��q���H�;M0�����`^\
���a-<z �iH���o}��{�=����7����^I����_�o]G����.���!)5s\�Q,(�u�C쪵;�����nQM�l��|ƽ�b{��l��~��ھO�V��Za��c8ڴ��{ʾl:�����
����5��߹���}���鯘��Ҷ��aS���6�lW��A*��Uv�!�`�������=/ ��<��_����/M���s /`�I���U(Ԕ���ŀSf���B%����� �wv�o���I�_��@�>u�?����7��ǣK��=��s�����@�0���N����J��K�z�3Q_�W��yp��ޢ��ڻ�G{��<���zj�]�կ?�?�8���gPVВ���M�7 lc����������8ڼb�+V�Q�3 �՛i^��)&���6l��.�E���`ir�E`��S׋�Gw���e�|fʅ8�����z(VB;쩦u0�c �����*(��K��W�� ��5a8e���⯚�[iF	��\,ˏ�[�8a���Tۏj/��`�z]vc;� ��Ϟ��%��f�,?L��տD5?���_�����?�Gܷ�adv�nPW�5�|���jM7��T��X7뢢��㚂KKJعi�$��;���" �!�����������<�z��X��M�x�"�j�k0� 6���y��߄L�@6�G9���e+����s���`���3�{Z�@�Īϻ*�zX%�I�4��vOK�	{?]�)�g]��~�����8���Ok��skWʻJ�Tt��>��w��^���AS��9'B��������1[�������0Vd���Y���2㶻ӹ��e�T��
�=���S\��VQN86�w�/����i�(�w��YS�b?��86a<��<�wָ��bׯkE��@���Sz������n�`WB(M��X�o�Ƅ�������C=����r��+ǬDdu���D"�β�J��sY� ^֠�U���_���g��]~W�:�����B^�����!5{n�`��^u�jS[_]u�u}�����B|Y�.W^���y�2�d��6F�2Sڦ��6��3��������2T����	���?����}��8T�s����np�ȅ^��e�����:�����f_<���6��ߥ�o�A���w�����'���{tqz�� ^=��?�-�T��NdJ�e�Y��-5i��3a>�_ߦk�{t��z��}�9{�����7i�w/�����G�9��{�9�;0S�� ����V�/�z�|-Y2�6��݇�b�C�OYr�j ��t�b+S���\��@1َ<C	���!��0���cs�y0ӷ���7�,8Z�	���C�VQ,"ӟB'|�~�;v� ��ܽ~o+(\9�b�k(�(Tx�`1�B!@P�*��^߁i���� �*��b�V���-�Z�NdB�@���ѱ_#�s~�!� ,fSV$^Av��޺��(%�{:���].q?X�����(*Q�XQ
��ܱ�O]+��#�h��T����x�?��~ue�:����膣��*7ս@�Vk���* ���s���j�Q �ʫ������y��7 ���Pp���fj#�RI��>���35M��̿j�UkEU�{�K�ϼ��+�;�9-�"�'�R��$G9(����Z:f�@A;�YtsYw�o�&���*-j̂Қg��J� �Qp�Q����=��Z��M�IӪu������yǁ����S��ZW 2��u��8g�[ P�Ce�]䴕^^#������C)�����`;�{�7��m*�ϟ���^�✱��}0P��Tp��#����ty&��68�`�K����Q�U-1}��5��j�ױ�m���k҅mM�m~��༊}~գm���������\�{��U�K�3�m�Ch���c�ץ�
��iE� ܃%a6����;*�!h����=�������n3y�����V-8�S��� <�g���|V(q�Y�K��"3?s��-�!/&��R�k�����
�5��J�sB" b�Pnݺi���[�Ι����y:�8tc,����������ea2@��������5/�^{�������sr�yuq����� q��!�)[�"`�9���_����ŭ
s�ꏨd���.��i�$��qE�1�\ME�!��a;�sdvrJ��K��B�@���	o� ���OG�<�|�:C������(ˠ�i>�t�5�$@�e��`�
���r�D����:>9���J��l��0/����_zV��|��7� �kY�ʺ-ؿ����hBg�=3*��y�c 3�WB�������ː��1��I�6�s�T� �����<�a\�,V`h�4NG�m�/�{��Շ�?�T��<�
���Eۡq5��
��@�2Y�`aP�x"+'~/s���uc,y(���w�$���G�xuw�<��>䟮;��(��{���ݷS�nAO�p��A���5��F���E�����(D�3�aj�d��3�#2נ3���u��	qYP�Ύ������9ƪr�	���k!�8(�(�WQN�+ɐ������/�� ���x�g4	=u3�qʲv9�)�ѱV��f���\!زR�V��r�z*���G�g���a�c�\�1���S���{�����r� �u�a��G�?�1��;�T�ۻ���� ��|�M����qTх�E�6��$�	�$Q���SU���Fv-��/��i��v:P�6�UǺ���~��H���x����Mڷ����ژ�W9�����_����%���F�s��Q�g��O��l|4�*�"i7� w���_L���g�駟ұ�����n�r��q(Ā,���������Ѿ��a��ʙ����̒�{ I����z{�G�酸xP4�nqe՗G��MUb t�����У������Kۘ�#��p?����?�o����cf�.�Oi>��A�Ϟ=ḀA_J:�_�؁��y0$y�sv?� %eX�U����:O�Wy8L��ղ��ujEp�{��]~<���3��8���\&��	��3�p1��� ���]�P�5JY3bZ�C7,X
���u]��9��(B2����G�Xsf"�W2�b��J��<n&����q͂n]��-JV
2���sG	��c�S�$��kƐ��}�뭃~��9� �Hf�P��ZDL

��l��\��/;���e��d_���4����X�f(�l�A*�t|�u�������=�>p�ߐm ����ׇ�|�V�B���'�O�����5X[�ގ ��9��{ ��{�-&�X��F���ܯ������=��Umqh&�h.l䴷��
h,�c�Βt��=2���u����p�U>���m���܀��-6p����g)�����p�{�w!ݠ����"�%�Y�� ��]�ɋ��{���01p�s�����(!,x\;�ۍ}��[��k��
�OR��N�5�y�c�H��8Χ�ځ={�`  ��~gs�����bI��M�?������Vr\�Z��6�է��8f���Z�{�mz��)�?}@7Qx̓$�@���8b|���`Q�&=vI�y%>M<Tg�+à}y 7��0v0�bs�� �2�vKB+�U����Um]w\Ũ�������:��C�N7ƶ�69�w�J�r��>��N�s�}�Z<�M�J�f�O)����Yc���~�чt�,
ΰ��I&���"�hG�]U��ߋL�z����������2��)�S �̜����z�A���)�G=�Ñٜ̋�ܹM{78�N7dV���\ ��Ӷ�\y��4V��-�:� �6_��Qa�Ϸ�ŋg����]�;�tp��.�cfz��^�`�P�B�W�������+�ێt>���b��L�A���%L.~gNdMnTQ���s��2Ь���璱 ����ΰ�P�e-D&>�p�7W3��I�(� 1�>��c�@8d�.$Eۄ�Y�
0��}Ƶ�4��LW����O~_G1��5����L]�`׃�J��S�y 	��(>�[�+���ً�#�u�s��m2�����̉�/��&(�a����}�Z^�{���2P���9 |�aak�Ձ�E�'�
j�x��u�Y���oGP����V�U�n"���ԙ�"7�,(b�����w��t�8mPE���Z-��ďu��rV9�joM��t,R����=�k4�*�A�*�g<���G�F�}���1^�|#�*��PKu�� �"ޤ����ꭷ���������j߼���?;�s���W�87��H�:t����(�<��Z�餏
��X�5Ta�	?���zI �]�Ă0��ݙ�lg�k�,���̃�Yc�,��Y�PA[	����A�xL1�����1����+e���>�s/�wO�>�f�kY��Z���ϊ�T�n��TUY���i�?��������Ӂi,�����U�} ܔ9�kӍ%etS0�jr�����-��:�q�g��˺��ژ��v�G��yW��\r�G�gٕ���i�]���(ϣ�l�7���2r�Nf������䄦HW�ا�`q�� � ,.��-�R�M�N�|R���&����Ym�C|�B�	�yU6S���������������P9�� ẑek[���/���HLoC �xĮ��Y�U�q9�h4m2K���#�+|�O�.���<���?g���Ƌ�G�U'G/����3-6q
`2��������\S%�B���I�p�j�^�8�����o�i�Vt�цbj�����8-sI��v12������c����`�K���-�X��;�_2PZpZ8QT��n���{�%9�����iDXke�"�v��# J��t��vs��ӃK�f�����%\��
Pܴ�<ډ��u
Մ`YYC�T@*�?��g�`ݰY!?6wV,yǅR\n����T�i�Z#p1�	�?����⹎bLS��`lP����z��%���?�7�ܤ��ޤÃ}��{9��/�sQ��%6gɬ�8N�J�6����ٵ�zl75A�薑��b�u_¹�%���� 0�m�T��.��:�Բ�l��Q���:��U�;�����ˢ����-�oܳ�� �T��I�heX}GM]�.�	K挞Wϗ<��5a�Z�m�r�}ՕǮ!;z^��՟�H���%���������yؑ�>��$��*��"ʥ����=yvD�y ��
�>�q�w2�l��z��{�����W�h����:opqr�#uͺ�5�T���u��X�Y�	~��{�T܍v�lv����5t�����nq!B�w\���+�����(�չ:{�E�f|ÿ�Ca�%�ɀ�vM�gl�h<��L�y<>z���sM����y(nY�kQ��!�R�6����&R�ٽ?[囔k�X;��Ӫ��	��Ѝ[&/�:���_����6-~�i�i5�0��uYw��I��6�RJ�귶�oʪˆ�I��&���dA�,��f�!F\�M=�3b�;��@*�؍N�԰9q��)A��@�%�`f@�tq�9��Α������=�XH�E�H�uش�����}aI�R	luR��/E` ܯyM�����=�x��L-`�3��V�� 2a??��?g����=�c���)ͦt���h
w���_it9f�BA,?a/�x.�Լ@����3�U����}^�������	]�ʧ��R��M�������Xv�(%K�����lV�	��9T+�)�Z@#(�}��n&11N�6F�
���Xk��vqb���L/�<7��6��Q_S)E�e�9��i[�s/:rբ� ��O{���Ty�~~vD��W��3Vs'� �R��p.5��@�����N���;a���!É�Ӏƪ�Ao ԋRlCy'�K@V�|��~6И-G�.?[���}��r���q�I�� uJ'�{��Ǝ��p]):���w�死4B5[(챎�;���X���(9a����"�?���uBIs��(��5�bNp��Xy��os��(����g/��\�w���w綿Y���,dF���	����6���>�_�eܹ��<����*K6�^��l(\u1��澖k��sd'R0�m��"c������k<����x��R�9�Hv�ೝ����<�f�t�]���{ #(V���nj�������(�o�'�&�CޯvOh�K��k��)���g��^]TƠ�c�����4�w"���A���㩎��H,W�)ʅgi�o
UH�
Ra.��ώN�w�=���k���t�����C:�=����o���=z�I�
�)@'�A�c���yWy'��/j�"��̙��X�k��G��T���b@��+YfYH�)�jX�v<H�����K��<�pe������jw�Ɯi���t�1F�_�~�1 \L�9�X?�����<�{z�q�f43Q��No�k��c3:99e%���3���eI�"J�`�p����>�5M�H�Сs	b��X�B��Q������,��G
��b[rS`�PYY)�OA�0�ڰ�X��oz~����f��}��U��>��R���-kH�D@T��#])y�]���<���Z1��,����2a�E��c�͚�9߃���,�<#����51��獼�y�4u��g����D�E��`�����V�i$37��:>A�h,d��6�>�������4�������5��<�89o"�E%I�&
|#!@>�࿼0� k��9[��JЅnR;$9����XI�JK1���'y؄I�)���M��mg�W��(p�:�#��K�irG����f��m�bn<E���䕱\�D��+�,N�����ss׎������lm�t�!	.��~v��[�NjR����u��$Gj!�2S~ �kP�W� �ǐX���]}̇���x<<�T���-�M�o�Ѝ��h�l;��(�P��>�%��e��|�7f��r�֌+�k��d��<�+l�`YkC�Wj�~w1�x%�����{�����j�g�!. ����.�e�2������/%g Z`�r����9�o���>[��5?�����<�D��ǂb��jA�~������s�||�km�q(���j�?�˺ޤ�l_�mJ�k�����̴ͺ����v���l�Y���P���p1��g9c���=��F~~���� ����Ӎ�;4<96����'g@�z��d�����=�HJ�"�Q��I�������+�W_�G��W�3�ĺ���(���߅�h�~�sd�
ܪ�A!b"�(��X���2:�
>!�����B*c�x�t΂�,�U��co��o`�;x~x&|�q.[�.��.��wϘ@�r�tڪ�.��0��{��<���F�����ت��X���	t� �63N�gm�;�V8��zY�^g�6���{�9��v"p�*mY��W�K��ֱP�e�x�祖e:�c|x�PY����PHE��2�<�/��TFE��.a�eJ-��H@=/6�u������u��ڧ��'S"}~�rP�~e�^��Ԇ���҄���������g�?3�A���1�Hᇳ?p^`C�La1�|E(F��9G���'c<�i݆��"pug�r�F�E���R��
��)kز)�݋sWM�q<��ʮ��aٷ��ɘg�iΝ��U5taS͋��<tu~�F�h���kv���.*^���#��t ȧcQւk�����%��T���(�v���Uq��L`�zq����q<�;5~�� �ϊ�3EW\���v��p��a�̸�v�\|��:��w6���B���eP���N�W�(�Xy��3�|��\��9@�w�y��M�ɳ�o�8�t�fA�׽CI�Ӿo�ef���|��o��\++S���O�i�r�5�f=?�L��ɺ����lX`�
[Y�Y�YP��]l�l?��������c��mmoS4N$Ulx�ec��̝d���`E����)�ĭl�UJl�[��+Cty1bK��-���gr
E���~��c:=��ݝ=`��x>��,��dU�d������b�^��k�wۼh;�pݺsSV��2���l*{ t>ru_S@�� �:0���R�k�����λH(�j�y v���:�3b�����J��4[bE(���=��CT�-X4�YJ�~��\�bű����N�ЦǺkRF)����i�m������u��U�!����U��MA����l忛�n�(�����e��fs��tq�����5�}����N(]� �4���%��yA����¹�`%�tp��y�W6G��^�s]�8,��H �������,�;��`Z��:� P�����[����|��G_�;B:E�$�e���Q\�
��ݢ���Y��lA��3/����ہ"7�L���
f2�$��WP@l���M*:kڴ�����q�C�k�Q3=mo����!�A��LM����%<[��N*�&����w�y��H�$�o�`�����:){R?��G�;�[�H��HJ�oS�9�s3�Ђ��t�=���z��u�t�=�
`�g��L%`��ǟ�{�8G3s�:@��oɋ-�v5)��ʃB�����Z徒1�5n`\VE�0~�m_��fq��@1�,~�u��6�m�%j����1� ����H���*�TF�p\g���gi�t.���\���/���9��ɕ�f"m��Ah[�=�s۔�t}�
���	�\k��z(8KE��I�ʱ�Yz]�D��L<��;!f����9�Ɨ4���''g����Rok�ױ���u�('J����Aj��e��	"���*����^� �-����Y�0���u}�>��u��Y+��i;C�\��qh�0>�߬y%
��k��*̧ϩ���̴���2�\������$�A�V����i�c���ʅ&g3�1�Q�4U�KWV*�^U	H�N*�R�*���p3��8<��<���^u��ݝ��V�[*(6��K���(��L��d,y����2�Jsy3�����l�U�E^ݨ��])Yk�!�$Lm����	�n45 ɠ��h�J
���zzvN��^`\�/��C�້k�&�0�$Wr����6g�(�r����n���ADs0�����+�uF��D����r���?%I�Àꉓ��uaƛz��/g�E�����]��g�}��o����t~>�h;�vA�/\ E%W~*ܳP�g��������R�e�v���,��zmη���^��,2�1��5!�V�@?�9:�}��#Ѿp��	���膠D�>ˡ0s@���h ����$��yM���&�c�ݜ#ʮ~���y�e���wb���w��ݢ����#������c�}��Y��ۼ��Q
>�N>ӹjB͐�iy�P�m�s��
z\����a�̹�w�+��|�R���녵6��Q�ڦ���C�|�c���=�r���1IV��C��3'm�9�U���A�����}Z��*�6�c��lS�*Z���X�A�V)��1�S�$�Ԍ���(k��N�������+�D�]3�2������ �˳cz��Sz��[�{\E��9;N��q�I�4�$<5AH�0���誵�����9;��杽���\p���V�����.NK:����˗G��0nY$��Q� �|6g�=�-��8ָ�^�\��� ��<p����|�]�y������3:�J:�j.?e]��f��ؘ�k�H 8ǛdetN����U������x�� ��/r�i��6�g5v+��в���Z�� �J��:^��_垫���X�B��=69,ȳ�el����wU\l誦��* DJ"!�- <~�q/�B�+�#`����h�5��xBs���WwB�0��N�)�X�3�_{�>����hwǃ�@LFCz��=�4T��s/X��N�<+i\�!����%�~�y��*y6B����蹘!�!f^yA��*��{�M��Td7��������\�f7��?����q�B M�!� ��8�2gw��
�a�^e�pG�ծ��f�EA1����g��c�i|��T�yP:��u���Wf/s �#�c�`��jၬ�nz�:��6<3�r���π�^2D9S����x�I ��s��9*���M�Tj��.r$R%V�D���}��d����&Cά1洓X< ��"K�}�����́��~�<2H��,��u�<��,.;��_�ٷ��F}h������<�b_H��WV��1?Q۠Ű�1�(�o���*E��l�}�g�^�nmJV
rW��Q�JD�s�ZP��[�&�֜�w=%T�iN8���ާf�.`(���{������T�j e�8����YI������C�V�8��#�c&N���Y
�S�!%"�Ir�!]'�E��>G��3���Ƌ Z���-֤n'�]V�=�5�~敂LE�K��Ht�gE�Z��m�}�u,���p��+����C��5��(F�Z��'����H�5b�}ͅ�º� b���������ݻƗ��QW ��]4˘Ť���;~8�X�8�dU.��q���(��������r��Eh@ɂ�e��=��<�m��.«��a'��,�^�̓}F����7��W�/
�7����Uml[\����ev��3샖-]dV�6r+G��ׅ���
��9��&�>T0�ܰ������PfW�x��R��MY��ǀHƔ��CHΦ<�)?_d�w���ݾy���:=|�;�.�^l� ��<��~�1=y��KG'/��&�W��������J�Ԥ#��O�ݡ�@*��d�e ���[w^��_�]�w�>ݽw���:d�z~yI�?}��C�C�۠_�z�������-m�
Z�$�(¸���UL���F5_��1
2!���5+d������a�����s1��������R}�g�_�
P�Mix����{�mN*�N�SLu�(���\�̇��P��s�[ ��M�4���?g�A����ϛ
@sͫ+
��4�׺x��	W��ncH8��ؔ{��m�m��'�}N'��T�?�̐������т��Dڥ)7)�W*�X��y��.�tQ^��"*I�\��y��+�E��M��8�q(�Ħ��E|`{���Ɯֱ6M7)�ڦ�z?+�V��qo�)����$��W�O�>��v���iz�:G��,(�R���+mk���)��/)Lz������c��5v�=.m�=�}a��߂em����	�[$�5����m7e�u�&��熹�i�I���2�u{�L��<�x���sd�\F�dX)%��B�E��U*3{z�L^[�9�~�ί����&V@�i!���'��9��ڪ�b<�ZcB���1z�L����sٚaR�^^�<�?�T��n�Ɗ������믾�BR� o(�84k�|'�㢎�O�� �iV�y�z�c���/M��+],m���6��~�ڳ� ���Ѕ�
�/{�«&�*���~�z�c)�9mq�جӦ�=?eW�c��[�n>껛�,��$( 9�!�$��j�y�ߕ�}/���Z)��L��]4ڙ��@�~�q^��},9�"%����
���E�^
\�}�^����+����W�ׯ���.}���d����1}���������HXվ��6��$a$|�P��D���o�N�����W�Egk�O׼q�A(\hFH�ǩ��\,mg��I��YΩ&!�+�TR��֬�(�?�2n�n
�J����../��u�+�,[ZS��0�U�n��0�ra�U��=q�@�md(�o�i;�֧��p�z��tp��c���1o(� �5A�]\��Z�IR�A�X*`o�����L��1j�MG���PU�j�UHDwtz�7��_{�υ��˙��Ŭr� �U�k�E��=��!�5<W'�|x[V�+���V� .>���j�E\���(�Vp��S��ڭ���lm
����*�u����f)JYi\o�ܤl�}��Ղt63F[0i�w�ޡϷ>�6�/�G��V�m߶��H����YO�Þ�Z)4ݠ���%���
�����吼���eV���l���z]De�(Ɣ�OH6�ʥ˗����.Wō���l%}$���YX_e�����U�Sڷ��}ދ��2E�IH	bE]�Fñ��e�Ɯ�x����+�/b�[角im�e�5u?�o��0R`���Ww[��;������BjG� #�� �A��p�4�,0���ӬJ�L�+�O��D�lQ̿<�L�3T�
�
b�g�qlHUQdc�ib��m��M�(X0�B@4��!Y�L;�y��`o�c��
EUI�mm�U�g��m����Tp�Zt�\����Z�V�T-Z#��k#ƕ�`߱J&:�30*ſ��`Y�릒���\\I`ʬx�/"�^���f��`�L�q��EFIy����@��@���-8�񜃈�r��;tp��E8�y!�=����`���}z��w���{�ɃO���Gtzv�
J�#�b��'U�ҩ���n!i����޽7����������~������͕�N��� P���8�� �e�A@�̿�DΛ3D�0o�'��~
���2-ͪ<�  ��IDAT���D�1�,*�e��&� ��X�>�!���#���
v\�Y�K� ��$�$WO�4��W?Vw�XݽN>��˼�W����k�!!�I>X����: hTʰ�d=g�����s�z6������؜y�RT�5�,ϣL�k�5��b-���B���:�1���X����턴lVB��1�R1VM�
F�n�SKN�)p=s�S2�CQ)��ݝB����>�\�k]ŮP�%]^��ɪ��Q<m{�st�:������O�*�⽃;I(n��ڹҦ �; i������xT@b�YW}���L/���>��T5縶M��Ne��WUu��/c�S} @���0��߸S��Q�}��
�پ���5׿�v2�����J�J��wr~���4�
���ts1��޼��Y֠�'a��F{P�[%[;��U��s�ل `��Z'�~� z�?��g�����H� �>�eY�qs��F�"K]��X!% �p�*�`�U�n\~�Ng�<�1�2S�~��Nc��Ŵǩ$�~��2X�秣KY�����̽{��h#�@����'�����\PVI0���23�+@<~뜲5!pH��i�sI�,iF0���*\;�*�d�{��O#	ϡn�S�V��R� ��+33ȫ@�cݽj�Y��~o'N���*f~�"���\rl9�A�sճ���]c��U�������ӪEm͡v1�6�)@�ބ:X6�ւ�������Ȣ/X�G����Ts��+J`ߐ��O�*���a�#9���"�g��G��ǿ���^�i6����&������I4��:HxA���߹�8y&dd-j�CZi�By'�.�Fstr�7�����?���Gl�ʯ����p<�g/^r{P �
c}��Ң<��jr� ���Z�y«���'c�s�o�qvG� �B+�ο6�[ob���F���U��"0��vQ�������Y�'��ݽ�e������a���o���υ��6��jIѸe�4��������K7�Fp��cA3��̴�m�n6eT��8�oT���; ���O��u2a��:d���.�.��-��`��
��u��q�2��<�M:�D5x����������r��f%)k���)r��w�!�2�`y�Y�V���=G?#Z���6�J� ?e�-`Jm�N}�w��
|lV��U&�)���؂w�/m�ܯ\��}3U�����|J�x��>G�]����w�Ji��A�GY�t����g��V)h���A*VllR�y��;�v>��8���i�M���;����-ݻǤ�J:� @$���7��W���
�u�&�#��3$c��{\���Ò̅��}q ������9-��7(�>.�9Q4��Ot��*
o��&+ �ݣ�S�E�;���#�� �W�������J���]h�v:��,��&5~�ф&c:X頦�m����N�U Q&x�z�=o�|�q_�vA��7�Xu�X�u���,�U�[�]e���.�& ��j�/�e�ՖՒ4���ُ�������,ɑ.�Y���FkX,�b�%�hƗ�����K3��H�����Qu�l�]*3��HϨ�>�r�LuUeeF���\}�P�."���������x��b���j��1s�g�mm�*�+6rb-I�,}mj��圾��=;:�����R�ӵ�wwi?-���3:yq�z��7��rqj�y���7($�/�%dnX:�(*ICR��2�OOh+�����_�����Q�o5����p�z�nɓ�)E?�yϸ�*�W��D�nw�"V`�i�@���pBH���*���dc[So����杁?�_�3��չJ�ay}W�@�s�Ja���<	X�D��rh�*�K�J��{��xjV+И{\%����JQ1{5W�������� ̃/��~�,�QCy��R���b'=����e�(K8p�_P�f��
�{Q��1K7��]p�=��d^�q@Fm`�T���:&�m]S�2[�*��֛��@pm�m���|h��y˷�����O�S�L�z�]
�vo���+�I���1�_oh���0�A��*���\�E9e�)�e^���χ��_����k~n���YLY��C"]p�1���	���Y�ᬼ��A�*��|�1Ix���W\��f6���c�(d�{v(��U�����^g,�@޼/��&W�Qh{���r���=�9d���g��q��
�{Ii���d<^�n���3�ݒ���?��󁐻������;��%���������[<�^<{���;�*�'V�o{���c+`E���럘��b�L�t ?����X*J�y����j�_u\T�;Ga�[�~�6���Wi����jc�y_�����^u/�����Қ�*�_�揄L�6�ߞ�7�>3KW�A�5	p� .յ.ȑ�5�|6ި1q� V��aUb1�5��k7k��	-֋��(
Q7����m��+���>������)&�ܴNB;��8f�זU��@%O>�Ę��щ(!I)f�1�ERh&�D� ���B=�7 �eR�=|D��������-��_҃GOӽ�?��6��b�p������NϤ�+��[�H�a��D�`V�oh[5	ks��ר����[~7��n�i�O��Tr��]}A�.Yw�1��\�Gߜ]\rȐYP��q޸��g�@.Ū.�lP0��h�b�S����>V��
�?}�~FAb�94H6n���
��;k�F��[��R��'Ў�A�2�Ƨ�g���#�l���y9ƛ��$�9|`��r�n��*W������X�aw���W�.�g^��(���l���0����6^���܈377����2׮g�f�s�O���L~�⟁�a�|o5Kpym���Q�@i�fx��vMS|�Ǥ����d\XN	�k�4�b]]�~�u���� 	�Ű��稀��̦�B'N�ÒuږY�4��F��Q���KB?������Tތ��1���7��*L1�D���L.�
^�1$�ZTiFӴ�Nϋ�n{��2? y���J _���c(HP��I-VqhB��6���#��1�C���\�iw��"��ȉx���֕؜w�{��~����o�KN_��u�l���v
�c=i�U˂�ǃ�k7�b�_��R;�Ekn`���?;����7�럥}�^��v��o�g�=e?]�/}A7B�V�̒���[Ğ��r�Q��/�n��3�����n����.��Z������Z0Z��f,4r̾�^��K�� $������P+I�M���[:0{ƽ�cNZ��h�cs��Ê�b&����Ԯ��b~�����IpL�R���Q�b���=,I��|C����}�����������UU�8L��Ij<('ј$�Pr>N(�AvS��t�zBq]q_2ЌRJ�7�5U9���l
	>��V-�L��ϖ"�4ǰۘdnj�{6 V����~�HƤ�e�ܙfЭ�Gb��Ի�mV�á�Տ����Z�xi��fۼq�Vq6��x�����٘�w��myMD��Y��T���[3tH���Nփ�+O&5�	��y���,m�Y�u�����l�`��!��b���c��XЧ��ll[[:��.@�z)	�	������Dr�n;Ug�c�� �^}�p.�<�IjմC���z��jUv�_ra�g	-`��
��<h��Yb�y��!�0�k}s��h� ����[���>�e��B�ʂ����c���-c��B�Cxx\��g�)�g�j��÷�LH��y��3��|���e�ٳ0��9&������[��=�)D���Y+���*�p�^xa���p�P�ٗ�j?Wi�(j�T��nl̪��Z-�6�1H���x <���h[W���[�C��U�̟3��^���u�cVxȥ�Ŝ��N��7��S��V��r:�c��Պ�4�����ay�}�}����o��ԇ��_s��R-�����)�H���B
���/�2
P[��j��R�jp
�Nr{�w~4x����T-r��N$E���O�w�!�W�UZ����L�}�촫�����c&�u���y�y��oOi�+�/8���V��o����N���)h�Aو��&�B� �[s�����MIw���ہ�m�7�"J��r||D�Xԛ"���m$��U�C�Q��ph� ��y:?����"��2�� "a�濆�߹\���I^ڜ�&��/�M�L���Q�@�xƠ�������7�Bb���5���m��W��������.r��v�n���L���F�?�l�K�gﳀ�j����n��vh�BDz���$���d�Ș��緙��x:��I���ZУ3,�y��6��$`[36�}(�uG�l	����5e� u"�
]�PH�i��>?��'EV<�����Ηb����0"�u)�e��
Tn��`xg��3fz�S�[�dk�Jv��i�F���ժ�˲묎�~|�@|���w��J��r��w���I���� �U�r8�Z)}�Q�F�Y6c �Ǣ� �>+E�����\�"���>����� �}f�����ǫ��|]���1`�<�kH��k�2A?�cן�����~W���J^J��tŭZ�_�d5����Ʋ7n��8��V�PN�M�J��]Z7�)�s��o9>Cse��c( ��V<�<���|EB+���,ABvV5c�af�F��A�Wt0������7�x�!7�1/�	�?ľ?x�DBt.����^C^
୪:ƏCk�����a6�J���}�۽����W���9,�	����ӗ���ߐ,|u9��r!�~H(-�&\<}�lv��W��U�W�W}U����);W������b��p����C���� ���,��ja��^(Ժpk���٫�V��և��'k���ƚ���.M�#ڿ�M��M���OOD�  o,V_y[Hg-�[|d+������ ��q�%����; XK�l�h%{�6n�`!C�b��:C�T=��(�Ig�4cc������}���4�a�B"��EQ��ÆU�n%�ڦ��-7�WQ����ö��S�Z�{eiR�qg��[�M����[f�}j�R˿u�V��d�s&�BG�9 �w{{������OҼ�O7�&p��k39�����`X��A+��7�;~l�K?HN_'�a���H��f��'���R��>`����Xl�a0��0��zG�^�"i��Q�������=�M��4'b��u)�3��c����-䯰���[�����JX@�R��;��t�cf��P�q�I������"�e�u@�e���r,��}؏���]>Tf(��\�Bg)� �[�zo��q�kx�i	�K��UJ>����eܺ�J�g�?N�Kp94n����k��j�\���}�Q7c^�5�+vm�W�J^#���1�ʆ�A�YԬ`��޴�Qm����qZ�D�}��{�~����N9���1E@�Dê���Ċz�͖󶷷�	���`cb���c�����C��
��Ç�����Q��~��y��-������c������Q�#(�e����p�è6nBzz�W�X�U|���W[�W�h�6�!@-q��~����������@ƴ[��2�	@��	1���dM�G�Zv��V��x;hi��=�RZ|���o�疰g.7{�v�t�<"����2_�ʏ���}��P�u�cl�k�����F�dn��h	�\���l)�4b���8�;��(2�9�,[|",1���Лo�����s�۷nҍ�������/y3�_�-�g�0���,�M���ʫq�]��� ��ZQ��lZ����H����ig3��FK�Dy�ɲm�̰d���yj��o�R�A&̂ӊE!
Ue�����k�=�o�3���e_��7ֵV�4��Y��W�t����fХam	H��˨�b�Y"�u����\�c��C�p��`�B,(�i�U��sp��sT��Jt6�8.��MB�L��7oަ�t�ɟI�;;��n߾Mw����;å��&�\��ZҰ�P���eem�l]����W��6C����8gOv1���b�.����ͪ���1W(�a����]���xw��ʌ'?�,�?:�7��$�Z/cj��/��+FNl����u��δ��<��������Q6���o$P��:�ǿqš�����A��+�����|���r�s?�5�yh�1��)��vM3dX�؛L.)�����5�~���h�݌�/Yņ�g!jCVx>փwS<���߷�������Y��2���i�9PkmbJȦ3@�>uekr�D镸�n�Q�2�R6ʐSP���mi�:�Z�^/z��Wh"ѩ\���!�n���h��:��b���'�K���G;����yc�����H�Ys���'����` �m0N��[��s� q��P�8�#&#�L^0W��ɽ,�����Bmq@v�B���4H�eV��cB��KL��&<9ow��~>���C��E+6| -����Y�����ҲP@�Q&��$���b����Sto6a ��EW4�֢1M  ����C�\$FU�>ҁ�f�Cr`�D:��?���M	�w����G���E��+H8Q�It���zV�U��*�r#�<�׏y�{���9o�,2�#�jd�1����Zָm$��|�A�oXKN����MN$p���}@ڻy�K.#�V�)k�k�tG.���^{�5�I������ɓ't|���]��ݢi:ś`� �:��ɮ,G�дƳ���3 H�gh3�]������Dl��t6Q��ER�,h,3I;Vh7�l`���..�s ��Q��!YU,�`T�'�s�N��ŲA��V��X�%f9�m$��Ym�ʤ<�+6�����N�̾a}�
��x�_nSߦ���Q�
������@�Yn�b�qi%V�*�����4��n	ˊ�Ú���,֋5-/� ^F^�A�XPȈ��*d+��$e(�$% )sȋ����Sj��+cq��=�t۶�X]y劭P�R?��;v��?PE0�f �H�sqz�	tX�!tn~)�%���Qk~�m�ԅ90pL�_,p�����"
����n�~����!�j�^���I�Y�������D7�0|/�����ft�b�g�C�+ q^��Լ�7*�Ef��Uu�f��'����ʊ��V3�sR�S��!CK'�6��OR�}��H��v����Z�s";v��b��w3s�{�go$���~�)��em���|7^r��¶��ٽzu>B?��+H��3km�\	��s�M��De���1lP*]9����N��)r����+�	
��[k�T�%�q@��"� �X��P��z�-k�_Z������+��MmOX��.��`+�SW�^��σ}d6���z`ސZR���b+�R��������٢`^C>�-����.w�VM��.�;󭓰 ����oo�2uc+�����J`z1_�������>��u�O��!����G`��u}� �֐��:?��rh��%�<�g�a52���	����"��"ɟ�4���+�v�����2A�	f�Y�ۉ�ٶ�9�I�|;��[�x�O����(AW�O��2�PWY3�:����a@�/T��,��1�K����'o�P���� ]P��ڹ���y�['��M� ^��y�ܲ�6B� ��´T�Z�Rѱ�*?ǹO4u ���D���n��k�1����!sww�v��6�!+�	N��r,nL�fT��P�P���WM��[$����I��MX�о����sv��@�*S�2���1����@�#�{�vR"\�'��u��Qa��_]����g;Wl�?�Bk-b�$����`)"U��L����o�`����i��@���O���5�x� ��} �(�C ���-��ƀC���
���K�_wƒ����z.xM&��֛�q�cvK�kuc��T j�bC�������j���N��,�w�<1/��@���9��Ǩ�$����=(��cǝ+t]M8iX�e̪��MD\�l'�:S�(T�[PC�4m���H��YI���@�j�2��<*�KZ�2S�U^ǻn=�Bge�8[>O@[��6
ۊ=�H���kx��%pA��;�78/�>�(��*���1$a��FxL!L���Rd��y�	O�ɊրE��R�b�� EPJ֚&
7v]+x���*�u�u����W���H/eZi����~or��&[Yݽ�B,��Ã�~��[�3`�1�l��ş����q�lYV�o���e�f�F�X�u��_����r�c�ztqU�kc� p�4�d���K���WJ����^�Y�B��lI�P��]�3��"�Mα^M�1IJ+����X&��zޣa���ࡅJ���^�\��q������m�A1=�=!�q.ޔ��e��gtrvN�s:�Drhzz����'�~yv����"��1�mA����g�,_�4^K�,f�����\��;�5=OBM��A$���;[�`�s�M�������.����]�i+�����`}�.F��Z��ˣ�Wp���M���@��K6�ʧZ\e22�d-|$�Op�qa�:�AƵƕ�v.c���m6��P~'����� =�t*ˆ�^�d�J L]+D��e-��Q;�x\�|�w����a����oZ��)�" ��BN��/�/����u2�>�+�-k�_E[�v{pc�����q�.=?����������ƱrS��/h�&���]t{w�v�����_�˗/�g?�)�q�_,��`X���*Td,"��Ԇ��ٔ,[ʠI7�F�UR����kwtL������Qs	��Q%q�u-��K����%1l.+H$&�6��P=�-��r���m��
��zTȡo�2V6*-84��{�nU_�WYQus�$��Uts��;�ju�
l$�|��❙�0(@��p��%_��hE�Fh 2�zƳ��\<H�E�l��Z�Wil&y���4�IR�.�l�콫ho:�Y�b,���/�c�ů.��R}q#�*����'������+�vԅ�g�B\
`�"-۳�����bc��Y��bt��	x �'I�[����/ߗ!|��e��Ҥ�-V q	��u���;�o6��
�=o쬏є�qx�~x-�oS)�"g�
��1�0��U��e�|������U�u���%����?+����)����:��TB��|��:o��/K��GVtQ`�CB�k�WR]��s��M��v/+�׏ٷ6N��s�4Ӝ�º;I
�|�99̚5���~���Xv������F����|ڌ�׏�_56f$��{� ����w?|���9�����1~��Pe�fx>;���΃�Z��Ӊ�z>_tޟԔE����e/�*m0ƫu�Y%Zm(��9��ڗ���I�0�>���5�66\���f�ڵ�}�O!���f�(ۦ}��_W�@�K���?�4��W����6+C'�l��[`�x�%  $�L i%d?Ic�䜾5� ���J,[�Bdd��Vܲ9�ƹ���ɾ%�S���,
�S�V�d����g�+��6���)�|��c,�e���0[�d��Nm�0���V��ʮK\8�<{J�/_��G���v�I���q�73� ����M�٣O>�D��Ŏ��fw�	~��s��=W��K��2f9�� �i��4�}���w� �S�#$ڜ%�`�+�/i�Hʓg��Yx6ۦ��g��RX-Q6]sg_������ �Ų��V����Y�|X~aee�yQns(��h����AB!���M��Z���X�eT~��W���.��D�m����F(� �-�
���>��W�i�U�'H.��4jL�g����:Ɍ��L#n�\?�saw�f{;j��_+,4�ژO*v÷J[H� ��b�;�� ��-���d6o�j��h���ƭ/cc1yf�6��D�Y28����ɷ"�2KF����� �*0�zEXy��!4�\�%~~�+E?WQc>5���xTy�>,�Pv��pQ�|Ei�Zg",�uԥ�B،>R5mhx~�	�y �@�\+����u�j@�@���`uH~�J�>�����3ߦ!��������U��?ǃm�;;,��[<��:�ZW%���(�&��J�g1��6��=d
B�D�l-��h��Qb��^�?��>��=lA�r�;� ���V�$��W/{���jl��Y�~",���RR=(��1�A�ؾ|qH��K���/L߈�aL='�t�/�s�c$��C�Xar^ݨ�yu����3�1��Q4"�  {j˟�wh+�s5 �o�X�|5o1�ui��g��jڜ����z9�dۏ>x��z��4�c��2��Z��P�j[W�����_ך��̻~@��H{%�/�.'�O�ה�	 l@3M�j��o�"t�]��Lm� �aI&Y�k��I����`q��T+G2.cL|:6�r�n�A������h��U@�|���g�p�>*Kcw��6�
�����:b�,x\9�j$w�^\w\	�b�����￣�O�уgG	�F��X�d��C<!�qgX�O�N�믿�>x�F�FN����gKx����'��&��@x���
�8KB�FR@U�����#m�<f�1��T ���h�z�d� B�Z�:a��sh�����\
����\�	q��=p�蟞����q�HG��t�:�O~�`T�rn���W�	��꒩�J�g^ �|�i��:g��VE5���	pO�T���sB����RI�E���%-P��
N���5x��fW����R���2�"'I�(Ō#a$bYQ1hE�ڥXr�٥�d����mI���BJp>�!+����$�J��J�(
��F=B�*�X{Q��|��ͭV%9�ƌ���\#9�&+ V\-vsEP������Y�k����xұ���
8�7�TQ�;�����x�����D��1Ҥ�����i�rq0��C{S9Vt(��{0]z��yŮに�C��7e�E�|�|��U
���W ��+��}�O�謢�0$�f���%�������;��^P1��2 �(۟�28�B�<c����~1o�a��3V�,�c2F�e��rΥ
y/eo�꒽���ӳ񈗳̗��g�YW)UC}EẂ!|�ca�!~��=z�����{{A��u+�I�3���9��m���9e��4�^){Q+���4��;�[��w�X�*0�.>Ɖ͂�%j�_���5���<���f�#$0��<��5���=��|�7�~���wYƬ������Iڊ*�'s��d<�7�?���6
:-�_�~"\7��Ǧ �i��1��Qk��r�Xf��i��0�^a+�ovmސ���W�QԨ�V�xcN�����5~W'�fhM.���g(�e�}�M��ׁ���vt���qpW��@r���C�VG��vy]38 �BA�_�BGkU�(��4	5(fO^ы�G�cO0�#ʋ
pamnɊ��|I���c�����b�a�Uo3(]��Hӕ����o&���?�ݼq� ^ Ԋ-���b7_e ��w�Q�u������'�
֘C��Q�I/�����{���-��^�a�Gr����r�
�q2I��^����$�ۗ_G/�o��ZC�k�z���F���l��Y_P�olNBs]-X���hɧ�A�l7��Hg���c�#癐&ܶb�
���UfQҹ�A� �J�cԬ`n�J+ JF���`�ieC$�2�b�^�%[��* �"!�� �iX�U�H�h��&e�0%��L[�|���z��jW�)mTJU�/�����e���r$����p�Jb�<�
٨�)u��0Q�Z9�G-�d��BP�ʅP)RJXo��<���D2�Fe���W����T��ԕ���WZ?n�o�~����*�畈��<�6XL�y9���!�?4��#�R��m��tO�Çٞ�ߗ9�6��O�����ljr$��2��
̺�1po%�k9��n\�7^~�i�C�=	WP��x�j9R��d�*s�O��xO�*�dS��~�b`l�[dWTު^?��Y��^�5��='�70�4Ք"�@&�Oϱ�I���B�)�x��t=��Q1��hk;��f����o�S�m��c�j� �I��Y�ϑ����xq�|`��M�^��<X��9p0�������k�3�[�'Buv4�~H��͕Ԯ&)I�x�H��ct�O�)]��-�r �����um����z �wm����6��0�ZL����o�!/v6�9K0oNk��6|E,�-��1c�XΣ�b����hA�,vw�$sr��cw��g�CW�����u���̟���^�e���x,c6�*q��F�!7����X5�x��(�ɞ�XO+`P06�%`?�q����>��p�$�D^TcQ��ڿi|�=}JQ�� �����9+l��cū��x��^�ϛ��[o�E�}�[���&���%]Γ�p��BiŜ�$i#�a9yq��M�{w{�
�=�!���D��������:=?�p��K��K�i�����oӝ;w���1[AVQ�3�HL��RL��
9���BU&�[E��ұ�['سn\�����+QD�gjP%_:�{.�D���s0�:`X)7�$�ۦi��n�i*�k|-<S�J!88GudOO%�9��� O��္j���zٹ�m���R����d�����q����5��d� �M+���^�gGM�f��s�W%U����R_~�"G#�%(cW2rB���RU�!!��T9ӲB��� �a�P�R�Ek!c�Q�X�:tRqM�5jG^Pe���c1nZ��*�]�ӻ�~V/�\(��е=X5�{�Q���᥷�[�����T�6�� ����P�]q�������f���Z;qx�C��Ezk��T��j�����y���ZYN�f�2�I�0�4��F[S����"Fp}���c�*F��aT�Ḣ�$�W4'���4ׄs�"������g�W�Y71C���WT�����/�믿N?������Ǽ��Q�"�m���H���c��O����q�s(�Xw2'<���0����l��@�� �-�#�Ӱ�#gl\�^ؙ�����S*H.*�)c6MXc	O/�ޔ0�]H*�[5	Z0i����j��d����kb�+���>d�A,��7����B��mm1�qh�v�����+��%����U��uY�,0�cWi3]ۢw��Y�P���
�p;m+�>��Y�D�I-LK�� Ik����,8�Z�}k�5C]�Ɇ���ތ6����Sn
�%�7Kώƀ��?�����UZi��=/�0ְa�XqhB�t�&��Kдi"�i���e����C ��X�G�on�%U���df��bN�'/�)+�����x������{��_.�f���X�Ⱦ_�<lVB����d���}�~��H�������@�_2��/��Wzy����	�����υ�����ޫ����ҧ?��nߢ	oNK�:�	��$��bt%�
Q����BbH��m��"�3�"Ef�Y���&�bf�CȖU��.�@7���֕���X�*a��M>_VCM7mQlmW܉�� .8�ބW$�AQdƶt!P`�s(�p[�dF!�9[���0�'}��]���!����*�@�F�*�k��QiE�k����eXݱ7I��d:!(�.,���\"��� �l8l���5�C�
.pru%,EY~���C�5_���m��mf�a�6Q=/��*��`~�r��{yL�w Vvs�gP�t������.���!��U{R9^׽�1�s��z ���*e��۱�������}CJ�1�|��y�,�8��K|p����{���2sx��m����?Nv�R��>!G�����2��ب��P��y���)�i�v9���f<u ���c�'8����ִ� \,ʕ?���|������qHCS1�x��)h��|��K.",���/��͛�pV0��RQk���L�� ��ۭ˩��#Ut8?�y6�ggO;u�mc�T�T����(��y�ٓZI8%"6�z��o�Cr�:��ؓ��ɲ,
s!�N4�p�{�2Q
�!��Ǡ��� 4��#S��̗!O.�F����@dUS����v�	�����X聈NNO��T�:�p�Aihƶ���y^�8VZ
�����(Ek^,�Z-�Z�G���a��j,�#�(H-��uވ����Ƭ�!v��i!7m[���E����#q���y�O]R�-�rS�ަf>����ұ#�]��<���������[�aض�yLR�/�s&�r���
x�$6h���.V�O�\���8�J�-��q��F�p��T������9����n#�a���{�% ����<��P�嗭/�F�ˀ�rw{Ɗ�V��|�+��'�in�gk�Uw��dqy�"a2�`6a1��\�Y����_�g?��^�8��������ߎ��l:?>���iRzD�7�k��f�Cz��g��c^����_���2)R��gg�Ⱥ�]G[LU�Pa>pA�~\)KD��>�;&s��6�S+V�u�0O��5��-w5	u&�y��T�w�C��(9G?���smJm���UB�ƕV�
�9W�����9ppc���<z9�����<=��W�?�=Q�V"�RZ�V��E3\�fe
}^�$m1�[d�ޅ J?ʚ:����G��CN�u���`��q�+��5k6S~V1{(lZG��$�5%���P�J��ϘG=��#{Ǫ4W��? 2	 Q6z��c~�c%r���s��dVgfPo!�9�e�1�� �Tp����Q(��c�3ވ�e�����b[j�2��V��'J�F���z#��e��7�-�/<���<ݞ���4��Rk��OJ���+�˿K�������u��R����^9~n�6��2�{�i��|�pO۫j��u{l�ʪ�0v��fj`\��މW�ø��B�<�sK�7p�/
�Y^�j��0M�k���t�:m�2��q��6���iQe"��v�_���*l*��|Rn��՟
��v�'����3�Ř=�����w�߾���Ƨ���@�f &�-���ܮ���H���X�4�
�3g<u�KZ��8��~�5�Af���7ޗ�M��A�x��ؐWOF�2w'���J �9�����`r�
�0����)/�Z�m�![?�R���Ͽ�"m,#�J��b>�����gk='�e�7��J�)B5)��:��Sc���"g+B�ܝ�dZ)!O� 1���X���,�箝� ���}l/J�7u�F���,!�>.��=S�������k�Y5U6�+��
H6}������e\'���I'5s��`�y[X�g;���h�����x��Ɣi8�8M������{�e���[�j��@�����Y���O�/�R1�h�>D��ͯ�Z>^��x(�� =��m-�|IN�o�����	%Pϧ�.3b�Ф~��ݺ�Gwn���q3)�n2h?L ����t�k����г�/����] �eLb�F�F�Б8��]V 5d�$I�nE���U��;@��1K�I!A��h��V�����[�B�������������sɃ�Ȭ�Wg	�?{��N�}���v�wޢ��cz��iR�.����o�Ia1����(�2���i�{�k��=��C��9�sk���yd���#k6�d��b
0@b��v�~!ݤ]2�/B�4G�S+��@�wrzB�=����FK�XRh��E����3Q��saG��q(ϐ'���w�V���@X9��m���Q�+Q�`��ۄ�v� uX�PI�vs�@����pJn�r��=��x?֞O��=��>����r�� ��%�*��}���s{�9e�dy��\�W�t{�og���k��҃a�(��߳�`˶���S^�Tu�]�✵q�G��,��̃����}�M^E�X^�T���%G,sqR��Y������*�rZ�$�_畤����9���{����Y�9=4H;����`�C���Ąik�{Y�{�*.���꼃ͯU�/Y��Qۃ��X�@��R�G}�l�h���"[�_���v�%9���n�����|��'�*�mA-My
���x��?�(����@��"���E^���������T1nd���+	5 s�KW�_���`���4:��FӬ�,y
~pxY�c\�_�Yi(g"��۲�](׍K��(J/T^Ϣq��V}�-/W��w�dM�6��v�/-D�����B�@��?,�[��$0Sl�2=�&�¢m��5^��Z!����q��sso"�Ijkw���}B��S���X%��-㜈�<v��$ �yz�xp�������1x��آ��}�{`-��o�U\1� @�����sI�����GN�N����`�J
�{o�A|�>_ɦ'G�t��}���t����n�Kx��.z������6}��{|���V( ��L�}�z��>N`fF?�{D����� E5S^3A����\c~�#��-i��I����V��.���9y1HU�Q�!+sӳ�xi��
���i�z���SP����6��Ѝ� ��Cݼ�d�̿nhҚP��vIw��������=���y���&�>;�[��?+a�P*Zqco����i綽j��פ{J[�fm���(b�Tv��	D�J�{���߷����z��iS}��%�����ӗ��n�%]|�-]&yy1_r�S���Z!�����φ�*�����[�k9�=*,Hg%s-�Qh���)"�Yf7`���E���Wj���8�HYV֛�C��:�����]�x9]���ރz�R`�����?���oki���*�.�l�!�r������*����/�R������<�F�i��Zc�dn+�2��h�a�%���mlfJ��W�JrqpH�Ȕ-����%�w
��v����	�K'fdiO��`��I�UmN��c�O|��gC���c�4#|N+����)�s��?:X�9-��Шe�s�ԚZ���t ���֒�{�)�&+Pgq�r�BѶ:0ٝ��,�����˹���<&1uH��/n��j ?�	�V5�U�I�b:�U^�^��=�y\g��VTJ��2A����B=��X��s�� 9j��Z"�B�b6�.�yحݬu�G־���5�u�0t.��j�i!3͠X��Q�hp}#>�+$��Z��� !��6�ڕ�0�4��� A4M.^�~?uJTiUbM׹��kx����0���wD��ѻ�ͺnnJ���; �X��(���\+���P�`�`����O�gT%�9��uYK�r�i|\j�R�.>���$d�%,	{ �/����{z����������L; :[��r��ﬄ�W_}Š~, �<X���_ӭ�4�<�ݴv>����O?e���mz��|5?�����@$��Ã�Ԯ洷=M�K����}���_H_9�8Ks������W�p��Oh��K;���oS�~PvM�� �4�RB��\�F�s�ֈ��V�S@�j�cg��X�4�����ݓML̪�R&�����Y����a�c�Q���'�.͟G�g����q��>�������/���zr�>{AV�	�G9>7j�+��Wn�~^1S�U�]/לbȯd
�nHLw��Yk�:wo�a����k;zZ�gQ�@�ከ�T�
�Øs4w��2����P�
g{E�l�Ɵ���)�ش�
��9ؠ�O��>b�#���<W垏76�;��]������l�V�Pe��Xƭ���kj;��|�ۖ���Y�B~��[V�Za�i�9�� %(,A��k��˘jxKx6�����BC{�P��k�g�����N	(cɯz>{�i˘�����yH���+�t}H���Py�YI�އ�=�"�p��8�5a��Zۊ�TUG^����n�{2�W�X)��%�&ٓ���圖��M�9V�sc��t����0vKk��m��t�1���2��r��:�ME(�"4����.�7�L��0j\:i��Rk>X8�oаA�q�]��Nn����5�K���Y�w9<f��}������2���7'��Z�'���d2�?⸚�fT����[{Ys2Z9�m��9rH9A��(dhk<(�����	P mV`���%o�k�����I$麠��G��a�OL�'�M�~�N#�pf��8m��]�[�H�e]��j� �l)�ǻr�:��;�m=bO�9|�]��� M�XG������M�R�ds脬	��Ja��\xS +�q�x��YHs,`���i�%�����&�>�0���xk7���Q�]pr��̩�L��e�h�#�D�`+!LV`�99|Iϟ<�'wo3h���8����w��C,�H�āq���	h��\��dok��z�6m϶X!�8=�9upc��fcz���?��g{3���[w8������S{�|����ý{o|rzD>d�l>���aM��	����ֈ���SȼԞ��ǻ��h ��E��Lȉ�6v��/��V�֕+�]�l���Xk�<�~�j��(�j��9��$s,D�)t��2G�yYr���md"O�B%
�Jr�z�������:�����ß��d���٣������B[�+�XU�
���0Gt�~�/�8�+f�Mvx�
�!�LT��<T+p��A�;�ާ	 ��%�|���h�b�* �ؘZ-��r{D� �#�	Ė!X�G��-���_R���^,8��6Pi�v4G��y��\��k%>l������uQ��8���D�����Ɨ(�UX��9�X5e�w<� ��E��߁��!�9�˸�`{�=���^����U�ǆ̵Ѯo@}(����V;ǿ����]���n)/W��?�����c��{]���PK	�-lA?�S�T���9��3��͡�'WW�ʺ�Чu�l+{7��1�����Au�]~��~2��ch�֫�v�~7(��vE�g%]�k����/n����c1�̎�۞�+@>?g��7�f�j\�D�`�J�T����x�9�
Ҧ���5�Y���O!}�ש�������j �q���&�Y���:V���j0����H��ܲ�ѣ�Սqﳭ��;�X{�ΕFm?��tx|�6�/�F폼X���^�h/�� ��q �n�:���;��Db��5��5O�L��Q��5F%�.Ku�uRQ7��b�����Nt��/4D��fL5�һ�:!fU�A��Y��	�2�ƾ�*����������V��
p l~��̃
6[H��h��ACm��j�X09�g��G��*�yO�����H$�J��Rg�v������b��	��Ա��B�F�����r�3����Wa�G"��8��̻��=�˟����oEo޾��)B1�/����(ͭ�$`���l2(���=��ѭ$�g��Fw^��
(��d���[z�@�'�����o�����I	���Ω�4S�ئ�=?:�D��Ź.�9##x�HY��	;�*�I�����`�x҃d���
�*s �w-�Cn�d���&�g�n��H�T�G�o���
+����'��,(yN�6�Z�qE)<HJ���������ߢ��|�E�~��_����c�t\�uI��c����Ģ��m�xo�a���zRLcD��&��ʛ�}$׽�
ft��ڼN��S�kO��K�����1��97�'/���lN�RQV������$�A�5j�bE,��J
��4�كL�3v���J]��v�[U�_�\�+1R��ZK�Kn����P�6�׽��?%H���������������C�o[)��->I��Gi��
��>�Qe;���W��u���<(/��?C)�M���3���)V�oٖ+�x�箋��\X[]Z����q�΄./�أoF0T�b�Q�	��+l���\�E[����5�򪣧�(y�CpI����]�q����X?�G�������_kr()u�J~��j�ȼc�y�[Q����cGb���|(����c��	��f ��/���Ũ�|G�G�;�qm1���EH�p�K�>M���.�"��0/�=&��wn���+�������'�|�b�����i�<�O?��~��獝[Ig�d�+.�7?s���� xtF��/_���O��c&d�C+O�F�Mzl:����B1���jΠ���� ��'�|L����Db���P��<ǘK2e ��-\�(}_�x��3��Ǳ܄�9�}߳��İ����>��g?��Řc�u��C��H���?xBO_�C]�E-AF,4[yF�@��c�r$�ZEV��]�G�^w�Ŭ�!LB���$�',ǰ�/[ ʿ�կ�=w�>8ا'�˗�eNF���}ܣY3�E��m?���˟}���\|jg&V{.�~�p�����ެ�Ԯ$�w'����c�[b~��b\� y�ͻt3]���q�Vz�ی�����������+X_�\�n-B�R�:XB�2*Զys1�f�\T��E&*�b3�#N?����eE��"ZA^��!fb�Cf}��e�-������@��ֈH� OjUaZA����"m�O��?��?xNwnr�#����C��k�؋C���"��[b9�CY�8��������6-�
C�Q���@E>ֽ���~ύ�q�g� W�9f��Л^��٥V�l�,	����д�J?�w���(jh�y����B��K�D�񨖺\Qϕ(�9�9o�Y�*v�_C�:�����L��>֑(l��`�1/)�{)�}L���͏�J��U��<tn���׷�Y��{Y���C�\z(<@��d�� ���U�Dm��Ua��#��S��vcvo^���&�6��g��o��6=~�`e�l������J��("+�f4 �R�cS<����}�х@��5�4�|7>u]߹���YR��6�{6������HMo��)PQ�<���!���\鏛� ƨ�2ʚ����M�@�׭�5t��O!�A��9�	��� �i&i���	L���Ӥ�3��reG�X/ TD�{��<H�@�V�T����K������(tl�N� ���''t�6�g/^�ޭ[���߸I��!]F�P/ٵ�g-
���������G���k��Wg	;^\�-���?,�xz��/N8=���溌\�������"��r��%ڿ����iR(�� ��w�~��C�;[�>#s��+��,�X��	Z|gVo+�l�6οϸ��r����>d�9O��]�cs���]e<VT�ƹ���Ν�	�
���ޏ$t���;zztN��g�����x�q�a"�RIN�r����@��[�fG�6��,.^@|4Q݊i\@˸����O>f����{� �����r�	(����Ļ����?��#���~M��L_}�9mOj��g�2�F�����*���d,�i<h�*:��O/^N8w ~�=�����\3N�z��;l�����5Fq��d�ý����i6�."��Fܧ}kH1�8�J��#9�T)`߄-[�%�p��\�,�&���"l�OR4GՁt����B��ն��lU���_u�p}f���V����1_�K]�0��"���,a^!�
 omO���O.���1=y���k��k="Sˢz�,Μ��
�����e�ްֲgȟ�s5��N�	�B;0��̔���@Q�$�c�Q%F�����p"RzPVF+�� �
�@��4���`�O�1&���E1m�~�%����|3Ќl��5MQ��$\<0��yk�.)�U�XkD��(!f��8U� �����.�6���^O�X���w��{P�b�K Z���V��A�6��]7�/WA�l���P�}�?��W��{��γ�(�.�ڑ_��e`F�����H��1�8P(n_�wΓ�����c��@,�-׎�'J�kF�	[�}�m�;��o���g't�,o0�Q�iLP0��H?
U-Kp��,����,�����>���R�a�z�Q���������e5��&�rt��'�C�!����������B���~��(Yۆ��g��c{��kS��}7t%�lmĚ�v�U+�#�A �n\�o���1M y<�(����qX���e�0��[�&�1�8u�R5�f�N���e�C�j�H_������E�����҃�=������۷�f�X���w�y���1}��9&�|k�$k+�e[�(�<cv�&)[�hԴɷ�Ejw��9mOG��c���zJ���[�s�M���ڵ&��	y�����:<��/ġ2 ��O/����j'a$	�uY���|N�?x���g����?���1r8IKr��4X�X�-����Y��QvC@���Z&18e�����dQ$�20O��)UIz��!X��~�M��6t�~	�ih��˲�d����7(��$euFN�]��dj��UR /�=ѓ�pC!� �vk� �H� �s I�=?gp�vji{�-;'3r�2I�nT�|,|�mj+�~	��t�'/�қo���Ø�<�O�|�Z�y�ۀ�����N��|�_oܠ_������C	l������/�����wޤO>z3-�4/'!��h��	 �(�t	�h��Л�����^H����U����7k59�w�y�^>y�~?��;J���;�/�  �ʷ m5G(s�H�@�2i���m����?�Q��F?��+{�*���M�l��4��Ѿ�j�WW��qR��v[�GeL�ȴ�E[�ZY�*��)H#C�Z��>��Ɯ��>j��X�Ҽ^s<�ĲC>���j�nHs����nq*V�F�k"+h�mz�|�C����8]�L����QόU��#����+����[�Y:Z�[���"���9�'�>�$���K�!�f$i2�.b޷���X���BE�W-��+6�D�It�7?�hu�d��n��jsӱ�a���>Ux)�Ӛ@zycݵ���c����� rI���L9�1U����y*͚�A���`�[�s��X[z�����x��C�N�U�'��1�
���������z��%̚G���[��������C`�+�l��O���d�F����덍��Iox(��f������2f�W�s�s4dk(�î�p�H�є���xQ�i�n�g?����Gi��Ӌ�O�qړp�Ύ/i�8�-(ݳɔ��'�5Һ\p�)��X�emޠ΃��=�tʜ�R!�M[��34�96G��*��`=Y���>4I��ś��a��]��HU�{��o�L��,s�6&����v�>��t��U��=��9�QB�����gI�Ro"jusG7�d3�A�u3��&����c���,.�^ �	�ۻ�)���=�kX� �j���B���&0Be���D���:k ���D�� ��۸�Aa��Z���➘$psk��1�ߺM���靟5n1z|�4) i�Z �(YϠ!㤧ɔ7��bA;���� ���X����i�h,�PB��C8@{�\܁���6��F�-TRFwU���$�M��)\�`�A��tޓg/��~G�ݹM�$D&V�!�`�A8����BY�B���@�̓��6�ER���$D&c���t�A�!$����*�;X=|�@�mM��(�p`�qRr�3M@w2q�~{zq�9k'I0t'������|���`f��7�1�A+����3b�#��0�0'��m�+�r�V��y��XPo%�`���{?�����zy|̱�u������Cz���Ï?��[w��|X���}�z���8�!7���*��wi6���7g+l�1m���c:><��x����n�#�����{ ^{�\��&�5;���O��OOΓ�|�ݥ��_���H�	k�Vz�[���w�ss
��
�?*�6����3 T�X�RϮ��O(���� �9�$�E�1���p�m�e�i��&��bc+��čW\}LU���Q����[�|U(rR���:�l��%˕-����}�}9PU-,�&���)�y�Hb�,`ٜ��Y|9��C�S�T�.v�z��2�q��Y���b�q��z`P7;N����.9\Y�6@Jw�8 _�"2|���w�d�	�ϩ��Ӝ�lȑ�hC�w�R�w��l�e�X;��WX�X��VG:KNy��{����v�24�{��~{��F�TUo��9�����_�yx�wC���.�}ٮl_՞a+���K=�6�� ��L��v�T�s��=��Ֆl�����ϔ�l	���D˧�D��$:'�0�=}���F[�	�f�Z�������.dӝm�_��T̋%+��lλ��̒�nDU���oQ2ڦ?ό��{X�_��܈�6:�K'�$DFB��]���"mPK��~� J'{Ǖ��F5P��Q̟���y~l{�8�#�v`\�:����:?ػ��}�˙��g^r�Kx��*N�d�������o�_���*�ݼE���7�Zs2�dV	[)0��	�s���D\DDCx�Dq]�=�� R}4�j���Xs.YϓI�W��RB��rAU����ً��hVl�E�*�
 ��ĺ�jȰ����)��a=�}w�ӆ;?��%>TQX,�*wI��������1��G�[;׎O,���+X�W�~��5,A ���!��Ao�v�~�W���������%������r!!FQ`�]|;[FH�]2�n9�E&3�=��F��X`���Xl϶��>ҢYk�ȅ�}.G\x	! #|�d�Q��p��o߽K�� >}������%e(��HM)*p�r}�v���JJ�BhT&���J��TQ��Hw�-o:K�ɳ�#��Ͽ����T}��g����Mj�Qz�������_9A��wҳ��υg�Nvҵ����#z��8���VjB4ƴ\!<k��%l�_����4)>'�����u;��O�x��3�@88��ˑ��"�~K�J�û�'�+:_��i4_4�@��[L!�5�N�7K |$I�ˆ�,�J�z��M�ZC�$b����@ro�R~�d��*�B��,̛�ֈE�%�S���prK*B`xo��5�������U�+�ho�憍����Z+����h���;�7�J�Q����YK[M�6�>h`an!��9�kP�˺������Nd֟��Bz�1���;f��s����xo�����=��!o��	MVP��gnD��!���Z���Q��{ݦ�i<q�7�᭻@��t�)Lkf�� ��0TI���BT��D�s���]HI����0����Hoɼ
�Z< 5���La}��c�-�����{�B 
P��/���u��C�C����U�떿5��僙���	L��r�0��F���3��k`��m�=��T��p��$��}5uDA=i����xr����ϿJJ�H��i�Y�'ǧl�C���J<|Jr�����b�� �t�~F�(���1��`��/�~M�5$R擝Ѝ5��,q��iՋ��)�Ÿҍ���3���W�}��0 �Bэ�R��F��n���*�b7�B߮*+c�b����Mc���S�c��)��i�.�>lv�Õ�8������[��&i�ߺq3��V��QN��d�%��4��P�?�5Ն�~�s}�Ν��Z�0����D-��\�J]聭�L��r�<�r`R �oM�i���y�ՂC@/��M���P�k�0kF%���z�N/�ѣ'tzzN�wv����;�n��
��l	�Rp���''O����	D!�d*�d0T���!^ZTD\��}a��h���s�dM,��k���9��߾�[�_��n�H��>E$��bүE!'��41�) V��J(HX�H�E(��(R�XQ�.)���e���#L2����Ԑ7ť�ligk�	��,0�R�e=���.[�F�����I@}�}��}zvrNm��j�����	%e�9$aY
�+��6�{��좋y fRb]���N�r�]��	H?��!�.[�^��߿���:88����5=?:��/��O�	����Ӌ���ϿNJ@C_~�%�\b��(�Ӑ��d��錞��?J�"	�qR̾���x���Hm��I�s��I�D�E����/�5k��u%��$}���YR�Q=�蘓�g�;�s|B��iR�1%,��4���I߽�9�x��aX��Z���&�J� rf`�S���3�Z6+<'�j�<���ƫ5)Td$�t��7\���@b��i��Hm�b����f-5��7�5=��K��$�j�{�}'� X�)�X�M;'"M��D7���Ь�"{����b�L]q+y߰|� ��h�K~���'�ؖ,I�![���J���eb@�{P�$o�X�*V]��<�y5���w��ԿJ�G�{ֆC�T���L��A�;�8��I�	���ZY����b��2�=��؅Fx`b�[��x��#��Zx�]ܺY�=�/�2\�~o�-_�-�3\	J�nm�
ȐU�:��������4����uH���w�������g5���4ԍ9���״{O�*�xN��!�B<Ve��Qp�I��Y���Zp�0�Й+^o�1ĥPx�sM��-',�`�ʂD�,a���9�GX)�K�A���m��/5S�9H�� �{���1�.0)AV�y�
Â�FvV�����y�pR��Qm&1G�{e��rf�<�>�9�k���e�Ƙ�v��u#�%�^x�F�a@��q�7o�:h�3H�q����ż�a4�)0�@�[l
(����W`4Գ����~5�ŋ�|�O���/�	�k�yڽNQt���~�bz�Z�V��69�X&K#���L��-z�Re! �m|uq�-��x��Ń�I����y7Q�6�E���1�j)/�z�n|.v�$6Xs�|&����"�G����K�cF[,@'���+�?��zF�L<y��������c�k�łtS�O��2�q_f�5�&-<�Q@q��K �;��uM�����������[��w���.�A�#��?��
�DȰ�¬K�a@c)]�~B".�.�I 䣖JnH�mu�\���$	���@��N�p�`�f��+T�-� D��`yO�����-V6B���/�_�y@�����/i^o���6+q���H��U�����~�E��9��O7�V.�ȉ�>Eڴ�/�{X�<MJE�P=����G���B���7_�b��f��s�ݡ˴9���<)$��J^GP�Nh+IZ/���W������ϟ2�=;;�i�,.� �|��`�(����m	�������	ݻw����f���zqyA�ǇL1�M���4M�0͏��/$�	���>� ����<M�=���Z`"��jW~4���:e���홻y�Ц6�(��-�A�T���*��V*e熵�:a���}U��]'�=����A�pG읓�I��jC)����m�s���\��H)�yϩ��Y���π�?Fn���mO����Խy��$no�]���x�g��B@4�Jv0��s{	��K{��.�'�!¦���~i�!2Vx�6��Ŋـa���tq m@ۄPz�n��[{�5z�6`����Z+��?��������+�s�oY�W�!/A����k%��sLY)���|�'�ޡ���{^z�����A �m����j�:-��C��.纉�H8����
����0��m���{*����c�&�5�}�c�Ӟ{yyJ���$�7��m�t�h߂	*.ig{;�zXԺ�{�Zn����Y�$ �;�����J�h,Qz�tkFbU�dP�,[lx�d���6������Ń��=FW�-��ug��(K�W���	m������/vs�Y��j��[��R��C�#��1�0	�����닪?{��7�t �6��*.���/[�#Q`�f�4A�8���Hl�����D�V�
'��u�h��ƩT���Q􄬩H�Ud�'t��_Σ�P�=b��%k��@bGT@�����Qj��Y�I>��'g�O��ٿ����ݧ��1-Ρ/9rg�������_|M���8���4�N4 �
���YI�J\B`��C��_`M%t�P��i�yv��L������[�4I �Y^��^�Q+�j�S����A�c�P�59��2I��e�<$	#a-���=T �f�>C� Z�)�!H���w.?(*O_ӿ}�=��_ѽ�4G�{Z�H$^�ؑ�	�U�2�ՂZ�����U��tƄQ��>]Q�Z�Z!��i~-�Ni�ܘ+�V��X���N&:NB���']���������ܹ8:ᖃ}���\Hj�%^���w?|C����t���W&�?F���9.�i����M��w�6��?���_��?~L���-=��+�G�%=��K�bF{]g��s�B�4��-�AL���.�l��+ުߩEF8�5�,MT���ת!�)���񤁶np�l�����V����Q��//X(X k
����n�R!W~�c��"�y�?���������םڿG���E�E(��`�"���g.� �F{7@f�w�3���9��&���/�Z�B��+|��C���1$Ԉ�4��e�,}(ඕ��Iz���аlmM=�Ф.����}�x�i ��=E�x�K���e�o�Ʀ�֯ex�W�]�~�kx ?d���g�tXLy�:ۅ����Mvn�Ԕ
�y2����I���B<١�<�F�Mi_F�Lm׮�M-��A�� �8��j*���WLC����-�Dw�K
�A9	fH{�N�d�~^:lԼ1/�d��!����okV؉������0� 'Qgq�y�u4MUF*@7ۤb��3��9'U���%��x4�͡�x�>O��B�ll�oYOݸn�J8]S����X1�nV����[X�
b��|��e,ARAWB�o��_+�E�iKXn�A��#�$ոa��|�:��v��k�Y |��G�M�
�`Bd�"M���Q�}��ַ4!��q�F���
�'��q#�U���V75O�FBj�[r�+��k=��P!io�s%�pV+kLԺ�\��k�c�����$�Y��$��/�(q�I����ik���5�P�|�����_%��5}��Y�q��쩦�8춆���v!iV71^bp�1�߂8b�L�F�t�==>������^��������o��5�/�D�ea�uP	ޏ��Y���Ո�e�wN�ys�W"|n�������/�͙��%�Yq!�F������ui����Ǉ��w�R�}C?<yJ�+P"�; ,[h�w��=x�Y��3K4i5-�-���+�b���j9X+���c�����S�n$/�i��<��LwEy���ϏbFH�0غq�V�s��h{�<���n��6�������-?�\�}�QU����/��Œ�،�E ŀ�d���U�E�l��&�Y�@$#��E g%$V�b�iE)�"9�z��YU'��{T���͈��t���nթ��}�����{�F�͊i"��ڒ҉?y�ʦ5#�����t��t�./��o���������h|J�6��~����]va8a�xh�%��Yh�����v_���{�K_q�Å;����E�uMS��@� �=�V阉����AP�(�,�|�j:�^�����;
^?������2�J�G'#��gAǉm�y�5��@���n �3��н2P9ָw�W֧+,+ND�� �,��)��\A?WQ|���#��خ�)kw��#1�Bd�ɇ�8�~�h
�rE˵�mdp>KtfQ�U\�D	a|�A�~��<�h�i�Z y|�}��Vi ���eTs��?˛!�:@l �^��f��vĎo�_~��M�ǚt�w�����3�j��]?_��O#��9����h�O�4f�����e��Oކ�9ZB=�Y��F�jv��]��+ʶQmi͌_��x��Y0w�n@�6�����ԑ���62>����&���z1M0�� �e`�Unq|����(��l>�8�B-�Xx<�M����Y��dK�Z�� ��3,t@q[�k0��n������ot�n5�Ѯ�n;��6T ��^>�'���\;�}G�%.2��üYr#9S}&H5���L�e�����V�7��i:b�	3�2|�c��.`/�-V�����t�?q���@�9�}������: ��m,=\TV�BO��Qe����ڂV�UL��%M��E~��`P��-?�BϓMʹ�bf vC�x���&'B
��\2{)�@��1��I��M�����sC;�ۏ	�?z�̽�ӷ��wn�#$�!��$�z���������~5�B���-�v ։3�S�*����8xݳFubA\����S3�[�NP���<#P��O~�f�����W^y�̙�S�BLСQ+l�3������8�$�Mܰɭ��\	U#\BL�~�8b���j���f ��<1 �X��%-&��|���ܟ���{���n	y��S���$кk�q#e!t6
[��W�׶�TN.���W�AI�(�6�I����/��f�M&2��.//�q!����S�ZM�5g�	��+׬-M�5�룳3��w���w^~�ݽ��K6\w�x��$���p�p�����3��7�po���#�W�k�(�Q����������`�f�D`�[ v�Y~<ǅ�&�鿢g���|����#wzvNS2���	�3�n��aU��
u�b7��c�F0l���E�Cd�E�â O�� >����k�W�#�m�L���W�����,c#Ȟ���6��6^7q�^��3˒�9{���+���Sꁾ��n��[ЮS�@˪�qN7�@�u���*������]��ޯ+��>���@C�kM��eh��f�N�@͸���h�~��L�U�L̚���o�)�Ϧɧ2�(ܺY���R �6�/մ^oh`�¸=<�SJ=/i�}�H�?���դ��\�Ԍ9�6ņ��8����g>׼��Ah���� n0�n�5�����:�9�N^�8r ��YY��7�,w��8果�~\��[�Q|�ur�ZN*�|7����wK�k�*7�f��"���EGJ �4��D��MR�F㌕J���x��z�&�q�5|���^Y,����=�3����	��ɭ[�L#I�]h&q��7�I8����f����C���1�A@&�;U,$@�+�q�9VTPV�+TqM�GX߃����� ��+c�{o$!)�_�\z���ϕ#�e�ZRvdW�Ԩ5����w��Z,����LG(x��ϷF��sKԬ�v����OX�u���l��I��h� q��֭�Xo�g�rm� NMJ#�*iY�\��l������|ȁ�ȈTZ%��hnXs*�m�$* `ӉiHTR���q�����n�L~ʠ����=��o��;׊�� pu �|�h# V% >�0��+o1����܋���ţ6�@�Znٔd�L��h�>���'4�������Sw�$1lQ�֔8�̣ދ`U[�Z�����N�c�Yf��B�e��(���uͼ����HpK�A��Қ@�����<9�t?~�m� �U)K�^���O�v���RQ�����&K�fIݘ�
�'g�)��/*ׁ�k\� �9^0����<�D)�Fm����cB3]8ay��w܃8	�$˪$k�
�� �_�`�t�M�I�X8:=��n��KY��
Иn��=��-޹�n��� �T輈�6�7�`�>|�" �@=��@0�-�Iql1(` ��}睌�f-	�f`�QKX�qi�"=�.�}J����$��4�B}*�|Y�Ep��P#.��p�%�y-
}���"V(�iҤ�vs�H�8��P��L�8tMS��mܽ�G�{t����lt����{9ͻ!Sճ@j.g����ȉ�<�_n/jjF?�h�-e�'�	:e�V���> ��ot��et=]M��s�W�� �x�̙-�͋[s�����@v���ʛ\��A�1/���~��(Psm}�Ek������x�}�)�a���o|�,M~����k����� ��?��������e.I&,���?�|�����3��[�v낗|s�sem��
�o2g�asmO�]�k�y��5x~��[�y/,v{�JC�t���N�
�н�(21	o�����ٙ���[�z��홉+�Di]6b(��)$zp�0�EU��!Xw٧�5J�X06|�� =�R�sm����ޥ���[���n��N��D����%�L�]�@єi��"��=.��8�u?v���q�;��v��!C2H{t��ño�*�[�F�,��<'���p����6���}�_��}²�Se�?��?\(��A{�`�Ի�M�0�D��Te׵��-��6=�U����G4������B��>WǴ��Tk���=i|�	�:���sYYH�p�[�d|��q'�B�n h���,@h�H/~_�)Μd��������?�o�����T���Ep�h�Wt�j~@�\�s�o|��=��p�?z�^ ���������� H���tlC7e�A!�Qe0u4j6Mve\��-K#)-!Jww+!! ݽtw*-K#ݹ.�Hww.�K-��}���|��|��sΜѪf`��u~X��G.�yH#�ð'��Թtϯ3no�$\�bIsH�rp�о������!��$��Πa4�3����L>�x�b��`?�Mɭ��mַR��D��`��]S�C��,�J� �/,}�|����ozZ��mW��.��C��wfG������Y���6�Ri7�BY{3 �X��?��_�42a���6��:�N���r�������9R�73���1�̒�Q��v"2z�L-��j'�g2 y)�=o�M��tʽx�Eq��l��=���(�7�ؒ\�y
ŹsEh}������&
���{����~_J��Ƀ��-]�^�;��!�ic���}��AR�x��;U<�'@�ǀ�8�#���na�,�P��=r��h�j�T��86u:��E��l�&���=�H�V�h[�n��N�ɀ1����>�}�HF�#yS�4�+���ٗ2e[O1��lR[F���:C�W��f�G�P�Ů���������V�)I���Ehk6FIO�HՒ�����c���iq�$��s�Q���d9`r_��Nco��;�%۪y������K�|Q�O@G���H>S'̢^T�X��{bf;��G߶0�D�~���;h��S����&�V$�k�;{�Ȯ|�'z�(��/�-a0��)�~�m8AE#��R-���!ds����V���������>G�O���L�$WF=Qr��n�M%ȋ��oif�����_�zhv�J�Dِ���u�F���j�3H&��T����^^xK�DL4�7�G�L�	G�*�iI����Q�.���H��o�7�����s:O{��=4cy��o9�Z��8 k��<.i���3R�C�!|p�]���дބ����d��d
�y��_��SmA�a+R�SFH��;^6�$����TH��_������y�����#��ӻ�!������!����p����}��r�v�=�>~ˡ[�5З��Up�1ؤ�y0�˩l�DN�]�U�1�d�G�F��h�t���h��^���Z���p�W'Hl���T��'B�7}U$Ç�h|�iE�,>$zS^�T�{���>�Q��pLe1���75�����fI�%K?��j�AWn�mdp�z׎��c������2>�X�.��9��Ta��k���ڸM�{C<:��3�k���ϣ���Rө��RϹ:UӼ2f=�G��ܔ�f+�ռI.� �=JqaS�\)��l�Fa̦֩��;��Pk"!zbu7��s�����BEʴU��eM���#�AU�J��s�Ϫc���~ !�ғm��b��s@�Ў�ll�U2�orRMQ�E37/��6u�C��M~c�m��l��������sN��w�s��:�LL�+'���O)ԫ�9�co�i���̙��<\�����+��E88����if��0/�F�����	���{�׸ ݄���� }
�?H��{i�b#p��� �����JlQ˴wt#'y(�Flyؼ6@�|������S�_Р���mM�������J�`��ǵ� ������,��a��ZJ�I�T�)G�*Q�P�Gn~	@r�,D��2OZ�4!7���u��M�qoP2�oZ}B^�$�H�2']���4��Z����@cLl������H��hL��JuP7�@���9���}tK�,�Q���PA|�\��Ov��/��hy���cV���OS�E�oI�r¦����Fq*��=,����&k}͚��g�;����='�g�1k��F8�#^kr�u�P�B<r�����@iF��n�X�ќP	����s(9���_���ҏ���&�
taU�u5�4����[3�λ3��S���5�.�Uws�IpR�e����ĩQ*M<'9��?#�K��d���A�b�%�<q,1������0�bS6(��+Y�1M�[���m�q�]�T)���9?P7�� �1��{ �F��Mk�ƪ��ҩu`��`F��5�-��Ci������0�����kf��	"O4ZNto�I�_�
T#-;�w���
,ES� �DN!hk��U�$�1[4N�9��B���Scv45��]� 6p{�L�S�4�I̎梓�3�m�:�k!zj�L!��u��_�o�@4�M����MB�+0�|"7	��>�.2һ*&
��d�&��T�JC���/�T\�F@�sՀ�m�N������$�+�/"��)r6�x[!������n�eF��5(gk)��5\?ؙ���Y$u=�+ݨ�3)Wm�,_�4���
���@;x�7^�&���wAϿ�p�� ��N	𯍽t��r*��gI�x
̸���l�H�V��8(nk���}��έa|��T�z�!�[1�����< ��臅�ʞ��uSp:����K���K;��@�k�&��q��`���KV��v!�FtR�����q��S���k���Q�T"����"Ě��Qb(�g�t7l��U����up��:`?S����m5#�5���˳�D--���5�VRxМ�!�������s���Gz��F˄d���:���� u`'Wg�T���͐�پ��S�WQϰA���o���P��j�Jd�Yh��9��s.wѸ�[(��W��%oYbl{�u�&ޮГUO쭔��9��(��$��S|��J$�`����v�6��D�B��S�{>&��ٓ�`A����j���X���!�ߍ7��з�7=/U5�E-%�Ygn?��m����鷉�����z�{H\j��]�K([
u��K��E(��F�����
�-���Z��9|~�6^|q�-����y�:���Lfei"p�Pr_��Ǟ��,^<5�<�D$�6���'���X��dh �&9��,$�mey+���T�j�K�`�N����X$�ĩT���ra��3��R����F.�=y���yQ(�������a�}c�ƅo쩐[i݌6���H�u4�����q�X�4��n�]���P3���m�1��CI��m�ቲ�f�:��O�2��	b���Q&��T���-�&b ��a8�����F�x�	��΂���{�#
�xP�}(�ZFJ;!����X��,Xd�)uE팅iY�3�)7q��7�6���&�>����L�.��\A�]iө|�<��q�d7�	J��^1���mG�gH��C�k��x@Q�/;R��Ӓ>VT��)���fM��"�_�#�޾Ia	o�����纴*JTW9�'a�@�7�E�ǌ~��c�a�Z�ג�|�n%k���ֽ�b��'��DkK�&����JͺD�[�jH���S}\�#�ɂ�՛�����{M���wǨX��7p�)�ߘ�)�<8�ͲIKK��s�["\F'�L��J�7��\�,r̻��lK=ů����tt"���|d��wy56ONC�9:O���Y���Fa��|]��]� ��jw]b˚a�ʰ`���b�e�=�������l����6�t�-�$�;8}m}pb1w�� �k������X���b��BJT�Q����>Ȍ�Ȫ�Hz�!U�	����1�nTs%!��Z��c�������F�&$�̱DO&e��*��փ6�U�H���@�md�������D*l��d_X���ߋ���q�e!ãێצfꃛ�_�^��K4'��xO�kN�1�t����j
mK7�q�hT���y�=]�/��L�E���'��%�<��J��L�U��bc�'�IH�@���vvΉ	{,��o1ʮU����'vh���������j#��g�[M��h��KH?ׇ��Mƚi�?���"�12T�f �N2ҙ�$��A~�����F���wۣ��8�!��bf�����µ%j�o�Rg �f���1�3'��n,l�9D����3˶�/%�fO���߂�l��D}�����Z��*͢e_����垪g,�b+�V*�#��U+WQ�l$�"��~�{��a�j�̧��LM[���Dڤ5Ɍ�a.T��ys��ʔ	-�V�cd��ef��Obi�L�.����T&�+�9� ����4$�D4<Sֱ���ws@��߽s�=(�DQx�V�8T]'������KUr�#���w]�yGo��0�)[�O�vi?�}k-+��I��-��wi�6䖃 ��|;�R�� 2�5}Yq����K�P��/�Bbx�ma��i����^Z~f�����+��8.ZΏ*^W��Ŭ�������&�G�{�;|��H������w���HM3������T�G1���7�Q ��(�b��5��{rˉ-� Z�����uL�a����Փ��dY����(]N,�.Kt ��3�ґ~m�����coL�b >�{��jM=��_��x
g~C�.ј���#��Q1 �_��$F-֗S�d0<�N/r�H��B�?�f	=�Vh�?s�4��~,*=0viE����o=-��8���<r��'���~�W��9s�����E�MG7�(���C��;6�ߖm����͉[��9q�M���2W��"8���ZK�����'t� �l��]��x��rV�Ԇ\��v��*���C�炅�a����"�ȁ�ר�
N��[�\zd��q��B̿�l<��+�	���?Mo
�٪}��[�y�A��P�Y^*C��>{$n���}�#��eǅ�.4� ���2�qA�Z���XB�pC�/a�������A�xG�7�䋖NtK�J���5"��^�H���QҘ
O�p��H�K� �]�����W�|������NG��P����ˇZDL�}�L�4���[�9*f�e%�i�(!��<��=��`u__����IcL:f�&ݡ���!)�'�q�*L<k�)�^���XfA��ES��{9<�c�O8��*�ە�=Vv�(&J�p-�8�!)5Ľz��_o�Z|k9F)�O8>&'%����eO�o곚'�ſ�6��I��^!/�4�rL�F��8zz��������j�*�C��n�ռ���;���������-rB�*<�
Ltz'�/u�U꽿�V��Hc��^�����+ KCzv~�)�i�3�d�|���;v�]>Y�=�z.�R�y3h�f��%�%���������d���M$�f~�Wb���r����?���!�8A�\�"q�G8A�r"Yƽ��K�'j�/xt"F1Xt�ʡOo |��I2"���HDC�0[E�W�tY�	�2���3O�ݪj5*����M^�O��ձ��*_;뫜a.�(v�H�Ͼf��/'����2͌���0u��!?���<�Bc�w���5h�g��Dؕ"?�j�[yf�2F?�N]��CF�_�`��8M�P�K����d��Փ)��W�E'��p�S��[�|]���n.Z16�2T�<@�S��Kn��=�"���X�d+?�#��h��q&�U�$�P@�?��T4Jy���+k�oU9Yv���Ľn ����N9��*&:n��l�D����`+��|U̾L�;G>��W�����U���J��S�I/m4�Q��ww� ���A��SB+�[��
fY�iڴ��&1�d
T
�h
�U��b���	�:�c��5d14(��������ݼ-~	�k
�E`��.�{'[PR��S��ٯ]��K��:�����8�a���3I.)I�@8ML���#���b?��UJ��Cj�d=��y~�.^�l���Vr��\�8\g��|$_J��D�	Z��0�п�uO�ɹ�1%��D���S�Q��c��
9���|��?�1�����a�E�"sc�6tr+ �M� ����c�)����=���[V���E5��B��9��tO�Ǭ���`�,��[����2�[�_��]�A�ǭ��.�%�/yfk�uYI�!�$oɄ����V��aLqCV*K#��u
{�j���Y�G�g��`	קÍp�)��~��c�q}[(�+�pj��+�K�����ݒ;�1B���"-�q)��]K ~h�C=��}��[w��U�ݓRoy>	�5<5������n�
Ыp���<>q�.B>��F_(��c-����t�A�d�����	K���}��{��y�������u�l��@c��9��w�L�I��}ڇ�1
�i��9�X`R�U�K��V�ޞ��V�9� �J}�O+���(�l?7���:Vuh:onVmm5:[L��<��P�ű�&��W#�*o���S�1%��ԣb-67���	Y]��֬4ة��<N�L�i���ټ�L�O4�}�O�R��|;��C�:����Y�����J�����"RI轔�����GM��k������T�Bn�ku�Ӂ��g�j�;eN��j�T^Ԥ�-@��ji�5��;h�z����//�ǯv1� l��z��Ft�ݶm�ML���q�v�j��S����@�!,æ �2�cj���w�N�邯��?
zl{=�ț݆m>��o�kP�3F�~5'J��>y�{s���*u��S_M���WG?u���L�ΛR/�ׯ��`��g����E�֫������&���@�>3�d{����ۇ>��`��X�K.�����E��=���^���WW����`����ì��Ǹ��q��X�}�yq�5º�d��'~1>:z����a��=0mW�zteO�:����WQ���^>Pk����/@��#�G�t�"�U��i[�ܭ�'���τ��ɗ��2�	�k�G��5��r�&�#rN��y���w����zg��C�V�cs��>Huןi������/�i�����gg�1<"BNi�SJrb8�d0gZӔ��Yy#kz���n�t������QI���-X|X�����r!,�皳��BK���HH\+�@۠�)�����ݖ\��S��u��%����Nr�1��>�t4̍���B�����e������QZu;y#�q<x����p���LpYW�Mi���
��$�Ĝ#>�v]��Nqi�o���/!EEl7[�J�y�XCP*�	Io��*�'���?wؖ�18��S��(���UW����a�h"�խ��y�m�]���1��Dp>� �"�������������U$�Ʊ_�23B&�=ۀ�O/ӈ??�q�l� ��_���/4/B;e�uҾqP�\爬`�`��W5o�Ϊ���cHz��,��7*��s8�o�s����8�+��/��(�}hh(P�c�]��SGP�>��K���@�Xl܅n�z!��zE\tݝ.����mW�Z��j9�ۢ
˂��IU�j�	?�('`���}�)�z�+#"V$��f.�G�S@Q�x_�I�����QE�Y�T��<�Z��L�,�C<��]�.�/��F䮽.�D�g$m�"*��*��=�SZ���m�~'~�uyz����2V�sb��*���p^EX�XmHM�O�B%M�s�y��#(C�`�}!3�$�9�A_�h���FqFi*�PZJ2����4"��hA>k�M����O��Xh����*���Do�O6��w�$l�T��Y:K�ȉ��p8�-��g������������u�>���؄o�QsOߘ!`��Ȉ�Ob��1u��xs�a+��R,y~I�M���=� 4��)���&��Yo(�o݈���/���_c�U�?jg��H~�/N7�X�0� �������!hÒ��9��+q�*k��6qN�@a�;�.Ƕ�]^|��u��g��Z�.'b���K$1)��I��M���>q����$o[����|��y��ti8�.�������$)�f�̀���&�0�|�N�!��30u(F���Lu�f���Z^4��b5hZ����}�\Cػ��M�ˎ�w.Z���� T���fJX�d�(�8
 ߃DE58��D���q�d����
9�˟52p7�����w�.O�
\�I@����.��E����u���n��ک���ncCk^���#��K��	���ӕl�m��	1O�`�������T��[l�|����NZ�q����B^_��������y�K�w �?�(��Gb֬��pR���K՞vE�ڹ�4a��OX�r���콾�?x.��g&�N2;�w������i�����K��jGek���{����{�rS�qf�d�J�
��Ww��J��z��v�-�Z=��U�_±���J�G�<������}aFP��wXԥui�\;9-�q�1_-4������=�%�x�B�]+4������MVkn�@�q�̫��=6jI�b&���䊅kP�n�Ѥ�-$$���%�`��>m���.�n@=���������st�LC�g��6�=��O.FN��G�	u�d�t�oa�$��~D��h���aaz�UX\��f?�T��? ����ᚔz1�_��o2�ޗ~?1����D==�����B7�_lz{{V��^�U�#����~_��7;T�������k������(I��[C�H/��%�?X
��(u����v�М�
��V�3�XSLdM����01�!��-�)�Q�N���*����\���a��o�g��0%�L}���FګܚԔv�B��x^}h6���\����a2�a��	[� ���\��Օ}��7���U�C���h_�B��5����/4�)�4��~7�.X��ڏ�)X��s^FR�Lߊ����F0��i����(��=��L�bQ!s��\?m����!��:�6(��ns��t�N�]����B��wqE'�oω})"Mh�V�D��ռ��<�^q6�:#�ϱ�����H�ոUV���:}���0ݾO�8l�<\�6��:���P^�*�����=�~YHp��w����W"���&cJ�p���.T�fզ7kl��6��y��%<6�zS�784/�����9>�@�v�7"�=+^�G����E��N�mv�+k;E�I��������[
ڏlz���:��M���bO��ѕ 1�W�GG��	~l�{1x���o������@�~�Ň���6���+����k��wa�f��5���B��]�h���Tp�j���sYo<�Ȓ#�)�<2�w����mQ9��ᓇ"����ׂj+])k������e6oj+9���g@������Q��B[�u]������t�w����y�`��j�$� �'T��kd���PK   ���W|�߮�  ��  /   images/9c4d998a-0b1e-4d84-acc4-3fb4cfcfde1c.png���[�A�=�J�R��PJK[�8w(w��.Žh)��V��w^,��<���x??��5��Z���׬�{�?*I��R�b``���H�b`<����=�]`���EUZ�l�z�!+)��i�����T��ҭ�v�q��8�@}r���h��a
k������?�'�KG�
' ����"��N��[�m�<?:Һ̼)�r+�oß����Y:Z�3�\y�����
�A   �I�Z���� ���A�@ �z��VK�w������y҃A�xu�l��� R��'���o2",�� Ab!�����ygų�oA �)�!ZУu,=��5x��/��Q�'�������_����p�-���Z��?�ѣ� n&����������s��9��������i����؃����~����=�9M	��� '	n.[�E��չ
�c�g�j�-X�[<,M.�����ɓ4��O��^n��WR%���BB�9�o1R�-y0*T?��U���$Ae��sT[	ޑm:봥lI�o��d�ll��=�]��T^)�T�[7�	sn
��B��uH�8�G���>A��9r�N��>�G�]� Xwа(�
@mo���sW���tvϮ�&�#�����������IƩUF����b�6��GR��Yd�=�#zc�^�ş�����A`�\չ�����ڜ#b�?�l��{�1{�w�2�џ����z��2�X�uk0�x��Q�9��Ər,����%U$7����τY��I{O^s���eK �"[��%�YQzѭ�eȮ����Eo� �WQ̭����>�2�"�����?5�8��os�M�C����I�FICt��U<[��)7z��O��[��
�<��	�2T��;���I�*�:�Rs6~if�'\4���l��JԾ�nS�@�W"΍��CJ�)��֠��1���������竞!6�6�Տ�G�<C##���F��������N��(P�ss:>�Q�:G�����T@���q>���+�#���*�+KIr�߉>�xòx��������233�}d�e Ir���a�I�*$�3{Sŗ/hi���9��q�Sp���Ip����l	��扇d��G�|%q4辍Z��/�;�$�8mW���%}̙�����哑����6����е�/���"c�=���FLE��@cDR���In�,.�\-Y��$C���1]���:?�����l�?}Fr���6�m:���W~=�����a��T�p���Oj\��*@@���XM�_u�o�Z�r���%$�H��)K�t�D�gԥ���N_�ffR}\����q���L1�n�cr�N%}~qa��k�+@��ӝ��>�����s}�����9��ri��*��*���"p��4!���Xw�&����#��<1���2�x�ގ�wo;jw�~4�C�����M=Պ��
�������pt�����/u�g���5�6��.�,�����<|ó�]��FH������3�k����Su4��:'���!�<���PjY{��t�����Lzn����C�֞S�t����R�g�Z^w��Ь��f+٣V	�J�_��;���m�~�ݩ�Y�]����q�rss�v0��@AC�dlii�.�0����=��((6�.�"'��6���#�D�c���iq�3���̶m��c���̎�]�+�R7\�q�Y�f{�`�>;o�}Ȟ��7�e�:�A����Z�ˀ��𮱱1�M�kf�0�\�Y7���Xs*�jG;o�����Ų��yc
��ΐ!��~�+
ZuQ����:����M?�n�E׬���y+4ica�1`Z���t>��.�*����lnn_Y��АcF��.%��6js0��,�\K���@%�P
��5��� �At�6İ�V;M���򡫼j��zz>���_������45�L(�\{D�\�L��������|Q[ۧ"�$����0���V���k>��:��d=6�%8��e�[�M�H��������������i͂F��͓4ԛ�Y�r�t��Š��)ԭ��^���Ԩ��v��f�|h����~�"o@���󴗷�?^�XQ���d�����q�0���]�6bv~���D��n5�r�r�`y���Va�H��^���m^#�a����ݿk�d��`A9���ō\��`0�vw��_KkFB���0�qrr��Y�}����a�Xh�X�n�R���]8�s6`�֦����$�38b>�ŸSf��p.<�+L�s�\廬�<a玕@�`�3E�")�����/���N��\"���B&N/��.5�	q�T!o�E]�3��X�l�Ӳ=��
��Q�Ue�Jbe5��\���ăo��>۔s�w���o�(�7�'��Q)x�h׭Fj�쏶��"��n�O>�gh``�ѿ��.3h^�g����7q��m�E��v�ۧ�Z����U@�N�b�\����N��j4�4f`%旊hϏ�f�qm�p����MUC�\7,
qc��9G�^�t��K�l�K��n_�D�`~,6�&;<<�4�[�]�D��J�)�ݽ��t�9�G����dxˡ��8e�Ы�s�Ѯ��⫞�y�SR �|I	�iK�������C�ݵ�����N��v��?����G���k�=|~S�-��PU�<���7�x���c�*�1��]�R��CƖ�y:$�������.F>�
���=^�&����WY@>eT�>#d8�J�~>�a�����`d%������S�X���W&߬w�$��'zh������U���P`��x����0���@)Azղp赏r�/ �WA�P�Dc��(�VU��N��s��Tԯ5��G��H1�vˣ�h���FCA''��O�j�g��D�L��2��=l;r������E��>�Q��`�QwA���n�N�sc�2�X�I�XE Ɯc���u�3j����Z��}~A+�3L��f�� _���Q��f�d�Ip�~�wS(�yZ`
���dk�!	;"��;��e�s �B0NW�H;qiÄ�i��_;q�-OM�:�����bEo��,0�G/?U�����$�qX3q)��Y\jZ��s��UlqAH�Z,�dg����U�W���G�[��y�@n��s� �z�4�ߋ�yA��	Qn�Kmߦ�\��E�dOPڑ���9Ց->5���*���H���Lw�o�ͩ�G���	-�u�����[R�׶��?��~}����v�oo��Z��HR+���OdT�b6hZ+�gbn�����1��y�����?��x0":XPM�R���.��X��gd��8q�Hh۱��6Z�Do�|~޽E���n�ۏi.�5ݼ���L=��cߥ�vt2�=��3C7��x��؃j��Co��=�gԀ@��^�E�5y�f��t7����ׅC�M��F�HW_���]
����}8!�s�E��A�T�ʩ��^.�L�޺Ί`�Oa�w"��6>xR�4u�BSS�����`��SӨ�%���6y7=��������a/�ҏ��}�S��k6xů�eЇpX~Z��mÒ/rܟZ9�d|OP��[+O�r8�]��%�1��x?��6.{����L��>�`�djTB�-Ź��VS��;���e�kwPIh��ӭ���0|~�$ܟO�(A�ɫ�����ʧj�ie��rH�����<�E���m�g=/��F�>w2��s�\��J�0�j:ٮ�}n�}ۦ\���Ű����㲔u�v��\�:���q�W� ���P�P���-B��Mk�̯!������^����ƻ���e�h�"α'���&G�A.ॐ�������|�Ժ����XF��J�����A4>�����ĳߵE�,�I������t,K$�5_J��]��q�'���]hA���?5W�sO{�ǥT6�с����L�Mr�����H'��_R/T7T���˼�}C��m<�rU�u������[�(�*BJ����Ί����{:m4�ڮS��4�n��*AJ�W��jǵ�ǯٖiʏ�m<�}I��32���e����d]d!m��� ��	�
IYD�9�kyH�}J�&�	�� �Q��X�\`�}G�ū]��Z�m����H&əU�f��B���ڻ�A���H���Lt_�y�4��YK�_O���J@�FH5.jIf�8A���,�ԝ��pg� ǩ���r��pkW���A�EN��gFGF��N�a>�ǃ_�F$en��|#���$L���w�Hܜ������Q�X����A<���M����4L%>7�{:�S���; �(:�2XY�6ڋ�	�"�%t3���U�@Rx�}z#NN��v��&��v�Q��#��|��i�|ꠊм?��ط���b���"�E� �?��	�{���D����u��Ǣ,|>Y������ο��+N��n���R�by��N�:�fd���QqZ]�'D��:���|�j�j��r�v��n1�栚�o�s?1@`��}���_g��h��x�E��O���|y���[�3��%���#�d �{Ԡ����7˭�fw��k6�ALb��'������qptӗ�yC�R�tP����[�9j@h�"x�Ǎ���-q�ȸ�g����!�I��M�Z�����F�O�I�X�D]���*��o�Q���%��~�!=�����.z��;�ނW2�*�/ݬ|Q�����d�X��cGb�$,��V���Z�xX����4H���k��΍a��r��n��S�H�P���mg�>j`�yʝBPQ�����c�J�iUO������P>�zM�K(�}�W�&s7;;;�J�����|9W�?b���t�)�s?)��&���������ÃF�ې�ɛ4P@�� a���0/��&�
��j d��߿� ��߿�l���Wp�5���ɗׁF��ņeP�����B��,5泷3OW��o>8�;��
|E����G���|�9bva�[#'v�����*$����?E��[��)F�>�^	_X������I�����sՙ���r��C�e� p=ҥzW�ѡ���K�we7;_�-DM���e�\̊�%55�UD��*ق�a%���'-5Փ� S�[\��`i>1[��~�����=��=ɮ���3�ݓ��r��!�kƜ�I._J;z�CK��΢F�3a(�!��[M�C[y���5�����}����x�[��F-Rp_=+˅53�J}K��Q/.���J�Z���G�K�G1N� ������w��f������M�07b���Ց�$��0X�l�8o�b����z�O�t>����U�o��I�
��D��In'��4eZ�C(g��l#���Mvc���i�����_���s���i�t�7�,N�s��=	����ܗ;"���z�J_�Iʩ�EKG��n6���n��J�&Z��kyr�c	��:��K�����Jj$7���|�]�HY��w�:�S.6�]H��'���WF�}�i:S�Ԑ}3�IW���
�z��GT�t����-�W}���5xU��RrgfL.�W��E�,�i5a��XZ��TVV�~uK��!��t� E�٠�^���p��@�����=������8Yѫ���������ӳ���\�ዤf��v�z��!�f������������
I�j���&[.WհҤ�}�=
g���Ltċuyh��P-��u�x�QS���S�ɦY�T���hg��s�qQ�z�-��Vn6�]�:Z�]�t�$�#�J�N�M�٪:{=^�y��ŋ	t�����W!Q��dV�8oKKK�#� <<���U4���7ӠT�,bg*ֆ
�����q��8��N��~݋Jk�ܗ�{;�J����Y�۟��n��xmWv;�w�!E��v��K>qB؀�e�9�-���n<ZtF��&  ��q��Ï?scM�p��k��-���:�=W;���BO
"H��w\�X�I�g�]un)sY�?'(gʘ>E�� RsF����ޯH�k��ё蛈�Z�Օ�IhH��**���R�2�%\��3}oKςn���GY��Xm�<���ʊ��
Ү���3q��fB�nZ����@S�}�ǳo2L#%e�m��g�k��8A���������#����J����@�h������Q�j��,^|��+{�舯`�@��|o�2\dp:�Amex��u���8-�H1?Y�l�m:�W�u�J�������5�SD�;-ib��~��)Kb�kT���a�Ȏ�1�Kjkk��`�����K���@� zs�Q��|���� �dU7٬��2?�8�=x�C ��Oz����4-���S�V9�W?>��A=M�uF�u;&s��&�7�˱kB�����Ŧ{��W�8S��]��`§!#>\�����
5��ճ����ȧ���ۑI'�T=.�E���&�����븜GGR�$Ƶ�ޑ8�c_⥡����������`���I�o��)x����KyI�1oooyò-�$SPD2<�Z�I�v�Ot繳5�ޙ�t�~���6M���ͨ6����J�y�^ ;V=�?�2�
��a��P}ͨG��R��GV��^:�_��ָf.f����ɚe�𡝝�2�*�)����y�����Ac�0��Q��`r�OAF���Z�;�x�dr���z���Ҥ�&OH��#��/���t��Tw,����:��?�l\�Zxl����A�����m1<��d��Q����j. ቪ���[� ��!nC���}������$o��r�T=a�ÍR� �Xvr��mX����������t�"�3�V������ƞ��lD�v�۷�Z�K(/i���L?(.�d����'P��(�4.��s)?Z�
U�,�b9��+���2�7���C'�����;�Cd�?�P���9&�@c�=5 �6��a6��:p��fs�X��u�|
+��o��,^��m��8]b���6n�����	[�Sp�p�Ga�A��y��6�5"�U+3,x��a�t>�hmm��Q'b5��[�Ez;����{���W�.����p��XG|Th7�Ǫ��M�a�}:����h3kX�N�Z��c0o�?��D$C��X<RJ�5\�� �c��$���.�8�9o������5�).>��̤�VA�F�vRRR�����媲�/�PL��r:�62r����Nw@꾙�#-�</�7˫Y|�#�����v���]�:�՛+C�J-ЧU�G�qb�#>��s��S|�P���
�C�Xc;�4���RP�o��F����C;?�씄��`[Nc��p�'�oCK�)oe];�
4~E�_������r�/(n�ݵ~N��� 4;���xx�"�4����-�G����~,:��R�N�������P�ЩJ�&���f�tR}���Jc쯢��������v���Q�����'8�j����wʓ�(��7�1Ŷ��@~ �N�#k�����?6�������E���!�c򹝽^����A�D冭7�6�%�+?�u`Y}�"�sP�D��AQ�)��ďU���/��\1�ܐ�D&>1b5N��$� ��V_~�N��$�L�d7��=�����g^3�uŔ9�4hL	6�����$5J��:���4I*"���T
C��H_g�����<F��#Ge������aUEu'�aK[���ӽ�)�W�ĩ��w��|hx�«<�P�N��m�W�88�L��kfE+��}E���G�*$�a��A����{Ռ������Μ8L��{NE_\8k�)L+�|�O�q�G���U��0s�y����W]�V a^N��-�7��g��t7�.y����T�a��8*
	Ǹ���ĆQ�BF�]L�
��c��Ǝ��Z�LeX�%%M�����!s4�F���>��]y�ߜ�.��;G��ȱJ�CC��d�?
�3D��p�%4��ː!>����R6�(Ay��"`�ˋ���`�@	�Ib�������o�0�4VY�L�fy�B��T�}Y͹�d�h�}Z������e���������zZ�e�Tf�ȝ�f���R�J��q�f�-�[L�2�~l�W���ؼ�O��c�|�ͩ`'H�WQ���|����}�)"{Ĺ��@GN14J�@��%��+?_��y�'
7]�Ͳ1���zV-�<�θg�!`�8 � 3<�>�1~	�������v�H�H1Gl���z��M�8vӲJ�5�[aXx�-���_�'����N>=����/�q`�n�����&�}a�g� 9ϏnYW!��>h
 �R uލ��먵��X��Ax5���k�"�&��h��Oir�/]QD�T���s��3�&���'J�O��I�H;���-ʏ����,�;�#���q��đ��V%.�S�	'�ӣ�zP!��E˧�11V
�	��:V�8Z������%����c��hk����c��'>�U�~5 ����·a;xX3KcA(^�+����B��_�4��)��d�Ɔ�
R����B\��/걹���0!��ve_�W�Z�-����\��K��"@�c��������e��"E3��Y��'��w����Zd��	4��{���,�λ	����맾-Y�λ�_"�nN"oN�}D���+u���3M��T�A)�VlDɿC�Gi�KŲ��O�l����G�ׯ�d�'h��C�U����y����Q��~Jߏp���ʋb��i8%ɈplL�Ɋ���+�dd��?���5��	���R�݇?��}
e�[u �-&ˑ�T �qV��B�퉽 �W�=����/�����2����xDfĢ�8\��E5�����뇝����2~}U���;0q)�&}�n�xJ!�ٿ�<����RD��ΰ��R��,1h��Pm7UR�/��J0�|U80:d�f/��6g�EJ����.�#�^� r����,+����.N)�Fʾ�B[�ч�5oaX��/c�X��`�է�(~�-&�f�bbO�NVI�M���L��2��Y�8}@��Y�����Ã���FLd�|J�V�:�F���ޔ�Zg�+���kJ�2�by�k�[��\Նb�Y�|T������A��3z����"hỄ �v��p��@Ny�����y�@�h��ϟ�|�Ւ�1a](Fk���XjB�v�D���g��f�����:�]������/V�_)���_��I/S����\��_;�r��9ν���iO�
���+�:.*Y���Q�|AnJq�����8�O�a�)6�����4>^ê(ቆ)B�pFLdqb�E/��y��"��������L�\npΝ+�0p�ޙ�8��U�������������w�a��B+�J|�^��)�J)��Qƺ�<�w�=���$��/!m�Gaz��]F�;�ӗxU�I#>qS1 �h@����:��|/�p��1>�MԘ�� [��?�u{)��(�Q���{�-3,?>\F��#ɔ���E���-5RU�O�D/]����>~v��r�䰤������3�}�e̦�Ԉ��}s��h#�ǀ4�I��~?S^"��z[~��5�C�gK��+B��*#">���[jP 7.�Uص�s�_ ~c�q-?\�G�� ����� n�~m:��$�h<�V�e����'�b��^zz���j=��B�V��$=3����M\���P�%�ӯ��vM�=�y9��� ��n�e�Q��m;7΍-�e8A`l�{���~�7̈#і��n�^���C�p���C����'&��in�V����æ�lԮ��q���4M�W��'߆{�l�8�6�{b�x�^��Mܨ�,����O������v���)�}9�c�h��|�Rq|����͏|�m�*F�`��`0��g��P5^��fTuP'���8{��3�7�=��j�`8���7�cG���F�Ԥsv�.ڨ��%MeEf<)���U$U977�ɪ!Z���)~ǁ����L5�֍���r B��%n	m�+M^r����a��\�|�xb�f9?�iD�����AG��o�F����}Id�x3�#�~k��c�F�O)ۤ�������K����nn���^�[��E5QSc;�@�y������}F�|bL��J�gQ��e�QI�ڴ�|Z/��rY�MҎ1u�7'��·Ē�+����`^9���4�uMY����&�e��Ԗ���ѡ��3��<Aj��_�<qF�IG46�w���m��X"6U[�5�O�IK2E�|S��_��������I����B��6H�k�/�f��J�T���Y�Co1w�!Z����<�g����J���١(Pa�Y"��S~���ݛX"V?��>r��<5ΡDi����f��"}g�� <�jSmY�wC�E}>�W�w�3����R���Lˇ���'ߎ���F	���0>?��'�Y�4���S�������=fEg���'6�@tc��G�9#֬���X�9��
�1���`W�?���-O���Hp�JH�:�M��ksN��j�Q�_e��Ꝫ��e�f�`�o9tퟕ�[-/��x���u��8��*fZy(dd��mA(C--?�9.-���}�F�S}�\�"� +Խ�g�/w0����۳aq����|�8�����w{���΅�1�]�J;>3N�5�&�5��r��ZWt�J���\*��+L#Ag��H�@�c���Y�nC��B��]���N�W �}nqr�Ѯ�5:7�:����9��bĒ�_��eׂ��{�2j����)"��ȆX�������z��cp,��C�df�2�}���I.��l�󇰰����7���|��o��I���]��U{�"����v������;�w�oAo�>��)���Z�g�e�Ȕ�2^�ԋ�|�����[�B�ִja�T1�{���+B��Y�����D���e2�M�����������u�:pw�^1��y��ҠL# WV��F�xӣ}���p�e��ܱ+!��}�	k.��Ƕ�Ve�O
ĵ<f[��z��ۣ���gEj��W��ζ���<�cq�Sٸ�eϚ~��{��؛��y�IBz��g������rf�E�F]���ڲ�R̀�第"<�-�r���z�)�wfNQo�i��Bs���D*�|eN�)��Qx��5}A��\y�T{�-�y�$7���ef�l���߄��9T8���I���A� ��q����H�_^>$H�\�E�	��C���Q�&�f��n`áwi�V<���YHj��������և�+��WWg�2O�e��/4��Xp�K|'��5f�5��D�b���^���k؈�JTM��0t��z�$fG�^��Tm}���i�m�z�+�Z��i�l��)�.9{���t#z?!*��Z����V�X$?�&�� ^g8.�8�}�&�&U�Y��e��}�+X���:��ހޭ�yc?ق�?�k��	�������l����G��Sr�Y��-W��0{
b�A� ��=��x7d�uDy[�Yq"���кA,�M�Wؖ���jH�9�����H�'�?���� ����\N�H=�x��܇��&D�{0C8���qǑ- ���ˬǊoO[�U�v����"�xHX6�k������|�� ��H2��s����b��>U�َ*�ep��Jc�2
9~[�pnQc�M�]��V� ���{(u���8x/,���Ծ��ę�HBذ�AAP�_�tN9���N���	@Q��ܺ�2X&[;~����E��Ģ����X����khE��*�(�]̽�큇�[�9����
E�X��?`/��CE��d��Q�MEWS�=�˘�:R7��)�Y��E����)�8�`�%��Y�^M{{{^c����*���n�����:���(׺2²I��"����f�Ab���5m�ӓ}ӣ��[�˴�׳@9� � �nY�/�Ϧ���U�}�#�R�8nc��y.�Y��2<_���󏴦�&ρB< ���_u����v⪓8"އ)�u�Ql'<Zۉ1H���De(KL6�G�Y	���T��YY���$�K;;8��AJ?4�q
K��}�<��+�[�C��˵oa����y�8E��NO��c�G�~���䙸b�\���/����O��#����΂`1���G��~~�Yd��x'���f=�>�6�6s,9�N2�]t}�P<�P�'�$5<� 2����pB<~�$!���A��Lw�Z3�iIM���'���)�P��&�I~G.F�j
�,���W-'Q�� �l�pG@ܫ�	�EWTAQ�T�"4�O�Q��B�~�d@�S�*�"��� 1����ӄ 8e�{�;��g��d,��t������}��X���;�t�������U񎤬`�jI��/�������x��ۜ��<KpeI�>I	�EuT}g�F�����`^1��~�"�y���-�?:Gj
t��gt7ߘ�Tɕ�Čl!����OR��ßau�K�����љz�w���V�x��I��	����e=>x!���n���,Rnė�W��.>���l��c�SlA�:&�F�J17�m}�G�j���!,
f�}�~=</�I�b�pJ��ԾY�B@#q����t{{7	�J}�ӥz�wf���Ј����Xc�'%`2-�)5�?��˽�T�cЙ����d�����v���긑��qu��~��~,���&CbXe_rQ�d�%t�� .�l��J�A�͵=��5Ϧ��z?�,d ����V���$��]�����֜���ϒ��k�m
H�FP{��#� 6�M���p�d��3�鸨J��r�;c�Ɏ��`�7��g����W	<��k�^�";��p�aOz́�^�?�)"�KK�a�\H�X���|��'�	$R&�Љ_�*b	4�7P�����g������~��I��ր�K�2�=D ����N-����n�'Ϧy�mI�]H��vo��«�|��5v����-'捉盼��L��ߞ�2�)8$�=yȍ^��g�j@ⲤnT2<�6�Č���i��z�si@L��1w���7�-7k�y�4R�ﳜ�����r'(��^~���Qb�����ܣ���I�8�"�
܆�~��}���_9<<l���E����A�/Y���c�σr��U�7*	����~Y���#I&v�>Q�хq�a�pR,p@��9}F�I���8kp�RN5�G��H��R�I��"���x9��¸]ߛ��r�d���_D�;j��.UC��x$}\�2�4���'����p�3�^ھu��� ��D ˞���(�"�B'��E�{N������!އ����\�i��xc�8K�z.��7�`C>�0Tc^���-Id~���5e��u,V��xS��ڨ�����-Y�叉��yy�Ž>���D��<@�f�V¨e@̇��p��?̵��MjA�������rȊMy���1b,z�䎪4��Z-+��ORaL���d=�$θ�qJ���f,sFj�ir�¹��"�`i����N-czWf�W�6��0�7��=ƈ@.�$[T5L�c�|�G�s�T�~	� �Z���!�p?�ژ�H�0������:&#v���7����/�m�5A�>���բ���*�t���~&0
�гJ�����m9n�y�Ĉ���e��H>�Vl��3�k�U�s�o,��..�����Ի��_��tMװ���.$�a��z8�w�}����=�����Ӧ]���N7��.o8��n�v��d��a4�(=��C@�A�>�h%���Y�8��A�JAI�s��<�A�0��_�+!��<�|3]��J�F�](�+:�d|�������ǉbm�IW�F�;We�э6//¶����Go�/���O�}� ����E:�W�C��i�G���?�p���6���;�:0����F��2��|")aA�)^A�����bǁ-��Y�媇�L����Xl�NjW}/���,����7&}v������N*={}��<�_��d��%��I�QYI��\�蜾HPu�r�s�I�Cpt���%�r�t^�{���|�Wz�nDxۧ�z����b�0Ŕ{��_��V�.�ZWp r9"��{m/H$�����|F�HV�^�� ��f�6>�i��{/����5��ia�ū<�y[��q&B��,#��J�Ī�\+�-~v��!Z%��ḡ���~T`W���y{r/,k��ɽ�F���g�n�7"������'8Q�A��B"�pV��[C(�9fj
�6�Wbl�J �$���S�q;��a!��պ��>�P�硾���@�{�W'���޴=��̈́X!{���cW��U�+T�$0;�}���=����O�b��&j�zTP+�4�Qyj�ܤ�4�����i&
����Gd��*CWe��L�3JD�@Aa�?�i���xQ,^%u�F{��a�/_^͡;Ī(��S�~�)�����H"w�i��5������N��w)>���3w� 99��\��N���U�t8'n�r�='�����4��V=����W�~��G�ສh:6 ��cz��v���wAo��t�$���.y��������.	�XBp�I/�pz5Y�&�e�J��E
�n����b��z���|7S ��B��. ��^��͈d��|��-Xt��h������P�I�����X���}�� ��o��&���Z��7\TT6z.b��K�îrX0S �=26���1�$��&����Բ�]�����\/�i�u2�3$
HjP'����s���$׾��J_f�	���C8L.J�x|ب�r_E��n�x�Y�nߨ$V����Xd#B��L�A������T�>֠�2k��\Hm X+4���*�糝�����j��%���������f�A�'?/�A�<�y^E<$3uB����a\��4�a�������o�X��RHH�"f�O��`������5Z�,�k�#�]��'�A:@\Pm�{]�>_�#M�qH�����ڊS�(�}�ܛ���30U���"�  �A�Z�ש��[>�N�p��";rN�.���t�(�Oլ�;<#@�iN,�#}>��v��`���f��r�Z��a�ڳo�}�$�_5L*���"��zj�y�DJ

�o^� s�b�~=�k��w�������	���t��� D�20�}lqY������QV�J"�\��ǫ�]���;l�<M2D�sRV,5��v�l�.��쇧p���i֣xH��2�N0`�9Pֵ�#R\�O:��;%�����zB�EbMW���X�N�
貔� L	e�]Hӹ�D���0�ɢgB����þ�K�45��F�¡��D2o�qd��Ҿc`������d ���틾������jE����x�r�E^���`�c��'���H�M D���������v����|a��.Z)-zWB�L���-��\	�$�n�t�4��ٲvt~I�Q����/��&7��\�\��;F`��B��k$�0B����Y�~�J@bK�;!�t^a���Ġ���ʧ��� (8�B���;̵�`!�,���d��
fz]h���� �*ǋm��*�K�B��/����m^�An�B�n䴓��}�74�GB[���9��+�����(����$i	P˗mZ!s��+1KD^�����:x��)��SOLyŃ��)Bj�b1OG���f7�UX��a�W=)I��������|�-� ���S�;VDÙ(!��z��s ��c\��h���N0)7�?:(KD�Z4!�'�H��7�g�e�(z��G����ӥ�SV�����Q%��}a�~�O[��T͸�)���s��(�z/_xj�'ɑ��[(��B�M�xWP��Ͼ%�_7�q�Z�}�Բ��1�6%����ԉ������/w�R��Č��8��~Ѯ�N�\����~%둜��[ňSC}���*�]�	;�7����% Q.�':���͌>�%�د��`T�i�pWM?Qig@(�v�v *�KY���:oQg<��|���q���-��ÉL��d������ym|���{ק&����N}��	$��q9E�~8����^��O�����<>>>H��$-e ?��{�H�0"$w ���g�e�����o>�e�����j��ze������֑� ��9��.n��i~��f$�ӱ�`9	WVǑ��i�?���RQ�(,�L�6��'��b��'�!M���W4<Y�SDk�$�c.�s5�v���8ݯ{��wB�ٔ=,R�M�3�,9R@Uv�V���^�E����!@,r��)-��aT�-��}ľT�܉��LP��H~��s��SI����Z�v��f�2����+�j��Y��TT���߈A�i�U��m��4�yp7����il�5���]��1kS�B:3����,���5!@�o��b-n��ݥP
ť�)�^ܭ8�ݭP��Z��]O�o��7�=��=׽�g��_��hf�!]f�[|�����dXͷ�?�`Z�,>է?.�S�i��uSW2��hҒJ�ֶ��-�� �p�\��'�5��r	'h�"E*0��~pCp����	�?+�wv����EUx;�+�'"�yw8W�P��,�SL�s����W��w�d$�@&sW;�-�PyJ���r�����x��@��N�_��?��ĀC�2Xi���c��7���阘_�:�L�D"��[��Auλ��]lY�ǀ)O������r�6w�;1P����zAu�jG�3�C�q�1n����ă�
�9�)<6�[� 2���՛
q8w-�+�*{hl@� �tI�S�{	�#9��xW�C8�H8�Xˌ�!�SM�K?c�cS�C�O����pe}}}�/*�F�J��D�?������j����'�� 򮷫=�2�q۱����%9~�a�����)�緖��Z3�墩\��M������瓗���E[������1)<̕���苏g��,��yd9�60���76и7ᴂS��T��W�I�L��.�~���Q�P|�&��ᇛ�S>�����t0/H(�w,I�+��CT˕m��~~�A�oD1�S�Gn�+R����r�l:� Ã济��/e�Z��%�k2'KM
]��}��][cL�̥"4I��K�0Su�̋��5{p���1�@Y6&�o;j�K���FZ_�T�T�-k (#u����d�<�IT�(���gs�\�VL��'/i2����)������b'Dd�]6����0,�~�~��b8���n*@3�8�����dj�s�}u�-�,��S�M��M�E��@3a�fuT_%T�lv��"��)w�FBę��9R`�xr �K5P:O�7P�%Ӓ�g�X����K$���}�-T�GL�r�-�s	[�>@��F���bsFE�W�H��[���/�|&ley䄺�<�Y�6]:B��b�0�[��H� fi���~՘����E	���F���k�#B���O����~���#sI^cY���
��E�ȇ�E�]Q�P�QI�k�:�������N���u'ްX����)��]������21��&[ܙ����\b0�Q�;�H\~��cD#_5�0
���J+�)1�^�ǜ��H��BJ���t��C�o�G<l����>�ĩ89V�3���S���j"iCA3Ύ�PK�B��PN� k�~�{O��)|f��+���e����v����-�E�ϝ��:���Th��2�Z	�a�m4�݄�V�v��z�@��&ܔD�I�K�A(x C�EU���\�#-k���K�ٗs��4��r�`���q��,B'��*;�fn�RI<��KC|^�[�?���y���ʊ��P"�:���cqqI�cD[kk�����[�{�
C��y@z� ����-�ը�r����?�3GGu�e�E�1��n�ƬO��1#�s����B2FZ2�GӼ��R��>�2q(N�ݦ;�pAN��*^&"����leA̽m��\H?���sk�����B�Cy��c��Rk:Zs�Jд��!|?��1���O�U�g��|;g��
�7�+��%0�8��wm��đ�����$|0�r,�sa������9�]d��m������g<!o�e�
���6MMF:�2/������3Ӻ�J�i�3�����{Pnz�Ư�|��Ϭg#�-F�ĉ�8*̐5~"�Xm�V"�����8����b$�"'Ǭ�s΄����]R�]$�Ytgસی'����%/�BѬ����(���u}iu��S'��E�d�����'s���}_q&s�Z�+ڝ��5zs&��G&D�_��3l~�۹?*�L˿=�y~��g\2%�(޻�RG��g:��G//�IV��"��fcfJbՍ�҃��o���L���RFal�~pO�@������cs�r��x�ɟ�	mL�ϼ�	��/ OE�<�cF��5r7�^�m��N��ι��G��/>�FAG�'ծ���O�R��D�l���t�������A0�W��fo��o��@��#�&��)z�8pV�؊�����m�<���+\3d�G�y2�Z9��X� �8Ւ勸�߽s񭅐�}����L�6,Rg�����J����<�)�6 3s���ia�*BGtA�F��F�®��@��%��g���
�2��6#����YA����Ԯ�5�Td�rA	u�%V��g<����e�z.��Z�")����Ӗ����G�v�3Mo���R3��/TMQ��|�U�]�8�*\�cu����}����
&iG�7_�r��t܌ޡ�&�u��(@��_΂n9��.}���0-��/����AIN����l9��R8>l��A�B�u�7N	��:?�Wm��\�k/�<��С�3d{�����u��t���*�8�"f���]���5�h�d����*π��+@IɅ@�� ������Ë����'�Q�/+���TL�v�0��ɿ.�+�_��]̑�v�7y�jcs؁�ka�d�U-�����=�R�J+�4p��
���t��1C6"�}S��Ƽ���|�M@��������<SI���Vo$[����l��Pʩ�|�ѽC
H>8j,w=ui��isq|d��1f�/��!ߔ2������-D�����0
�S@Œ�u�Ш$��Ӷ�W9�?lhQ)�"�t st{�	�h���7vNw���Q.�;�@����|�>�ԟ�JBO�a�۷}�e��S-k4(ңK��	����(((,�7�c&��}��#�UI4	|�:��c)(��͵I"p��b$����x;e���*���θ���BQ���a;��y^[k��s1���J�cQ(\���ϧO-��4©-G�u���H-'�P+�#�Z�]̳�c�x�E�`X��'R���F���0�\H��QC�^��<W!?�ccɬ<��	4�t�A%	k��g� 6���<��������y���x<�}�n�Q/I�	+��������Ι���Pe�qp�5�`0�~���}8���(gzT|\�Q�\�m��<=�1��,��B���� `�F������_f_ө��Nߧa�X�녇��֟<����-��-�l�]B�����Fhs��,���/��p�"�$�<!eGԸ��}���s�b�%��?�ʠV_J��%��p����"7F6����:uS�.���ְ}�)�'��فUX�B���s�����Ё�8%`��_z�y��ȲdJ7�c"%�����mx�9�$tQ���f�.k���?����J����{s��rW*M�,�{O ���<l�!� ��Ag�'�Q�N��Q�9�����c7d���o��Ql��]M����D��J
P��Z�ϧtE��#yٿ�qV��RS»Ӂ7�ؒ�K���Lvm����Q��I���_���<.�S�/�B3�|:��٩ (]E��!����愰�� ��)|�����u��(�IU*��>F$����K��p�nDQ��d��Mc������Q����g�T��'Y��1�:��T� -�^zܛ
�$e��q�R%
�!���D��
�!I��5��T��O�hDBq�*مc�>BR��/���#���LIL��u��#���O�'E�ݥ��9�l��&&��N��hsonHw_a��c�C���mmTa5c>�&�|���ɻ��f�f$'ߔ{��s�2�
q$	����Y8=����k]�L�+�]i3v�3���m0�����	�����]��Jƒ,�yw��g��|��o�Cps���=��m2D:)�������<e*. >��4����9�S�[jtײ`���n_�g��ᯠ���p��+����* �B���x �h�������Y������Ԇ��0�kY/�zK� g�H\�_���S�+�ȝW�F���� �\� *[C����ZS��Y���4b�d�M��A@,i}��Oh2�-��W.�T<���I�2�����l��^q�o6���?@D��i7���CE��V����Q�� ��������ގH�+�us#�f͉0u����i=O��NB���Եy4S�
�im6��s�0C^�q��O�=�GBh]�S����ЀT����*{B��{'}��|�۪%�r��9���ɳ�qm��Ԉ���E#07����9`y8|� �;=���i�<�U�7�D�Ȍ�C���MH
���I��~^�nO��pe
�I�q�=�Eə�prW�o��%�`�!�*v��(���WR�k���N=2���]_haf^Üe����E�����s�� �}q&��A��ϐ�IT�H�c��Z���]�:/��gF�r�hѝ,�G��G�ӕ�)���Exu�������T� ������h��O���WlD/�33.���6s�C������)���5�����Z;�� 2rꐶ4�'T ��^�-�1H �`K����"�L��+��N�	=��!����[�u�WG�o4��fM�����s�Bt�!�F�� �r�V�*M�,�/:��Uh�m��h�i���[�O��U�}�9Q��j��~W��ġǾ�D �O�;���WUe�QU�$����[�� �pf�6�+D�?+}�*����KHU����`�+����%�~�U��m�_=�e���QQ��C����Ӆ��!0=�C���PM =Om(�$�md���N��8���@9N*�@M� ��NboL�(����:@J��/F�߿��$��� �Y?l��?dTK���pŉ�6��	}� � ��+�c����N���ֿ�U�N�:O��}�ޫLَ(��
��Ib�<��v����O|��ʇQ��X�`ПǴ�Ii�5�FN���J��Z����,�T��.4.���#��L�m�M*��Xs�ÇY'u���p� �G�C�� ~�|Ǽ^�W�U7�ɵ����}���ƬM�.�������C��kFaA�>�z�eb�m�4��B�fM��~��]M��e#�[B.�A��7Jc��W���%g�D@��Ӱ��0B����g�huX�Zv�L/%q��gVH�P���q&���=�cr��)�g�h�w����,��ͅs��#���DSG�9�Xd�>�x�7>Ј0��3x��Z�c�b;p���@������!5Z��fԑ>]�KՉ��l�T�WLC�ޮs(�@q�����X!����-6N3J�c�P_����l�V���_��޿��+jl�{϶N���R"�c+��y��ݲ�?j��ؠ��kّh�^/��3��7���7�{�V�lG��F?��f퇘7P��Q�%��677���c���<~�GjV����'KvG�H�n��!"��
E��C���}ʮ�4�1R�fПӖ��Zd��mvo��}�N]ɔ��41��=�Z'�Y�!u:�ա� [%*Y���(�����d9`E��c���9Ş�(�N庍V!�"����m��M-�%�0]���$�YOƊ_�:Kqm�#�A
������:̫����ԞTZ��<g���o�褰�;��s����$�t�X�� ��wc&�¼��lL�鵙h�RP!��8�(<�Y���{q��8��/�ϕMK�9�����˭�j59�X�S��e�N#ʻ%�����#����9��jÖ󚑑��Cq��	<�X�j�)�v 7Y���>{���:|&k���̜#QUߊ��OZ�J�.��K!{*����{���q�h���J�1CI�?��>l�i#S�O�J��,�����xJʏ���� Y�e�`�c��$�3� �eY`�Ikmj�^�#��p���d"Ũ]�Е��BRb`��s��D��лO/`У� !���a���#�o�(p��{��q�q���^VH2YKn�M��Ob |�!l�2�:d��/�D~¾y������=��5�$��曷��)�1�J!���wK��
����c``Pq�B�*����K�g\6������=�Vf2�?�c'����9x�f�#_��{����#8l�
⺩&׾NC�Mᔆ��u �K�$
e�Lxa�I����O�1�b�-V�#���m��������
m`k�jDSJغ�b�
^�t�6��@5�fT�u$�GitU
3t�[t	����E��e1�sǔʮ�۸�� ��.�G�s��e���Ƅm���Z��d��1X4���kz<�]�L5"6��R��2�JI�9	Ѷ�"���.��ѷ��c�;R�(#�8U�\�̎Y����̮��L�.e��ց�����>�$1OR��W���D
��R�!����uBz�!��0�W��P��u�e�������L�0e�_��Rt��7�pO�O��t+�``�,�cB��f)6���"���P,��t��8��{"y������~C!KP�QLp��y���H�5ʤ�1Z��%vV�֝��ƕ�u�߅/p����I�^���o�T*ͨv�����胲��ŉE؀;CD�T �/Щ2��F�f�!\����k�TD �H�Ɂ��B����b���R<iϨR���1�I�c��߃]/Jo:�����6�hƂ�	��&�4G$
�]uM��I֡ͫ�<����AF��\٥�S4����̽t�g%�%�h7�����~ֵˠ�r�1N�aJ4�uU��i][	�E��B^:ݞ�1��6`�ǚE��U|܅���D�a�<��i�S��8嗔vU�^�e
�77�!Nt]v��I�m|B��-�z�e�k��] �v��s���?�T��u?a�O{�ɔ����a�e������Y�^w�6]���_���Y_f��`������Ck[�������G���E�.뚄�.	L�-��{8o�U��ck���k6��_V$�?o~�[մ��=)~�9o�[�vP�U��' ��&Dݖ\|RIg]b*Hό� O��|=�ΐ_ԥ�<��6�@�d���	i�t�k%ԕ��"-z������� R��Ņ�4+8lGU�Ct���F��l-t�Ȓhs��Wt
 <�}61�1�����a'������Q�6���8q�߆�W���V?�*(��$�HP���Ϟ=XƹY.�f)�E�AJ�g�H���7���c��}K�nlkSPTT�Hf	�)�M�NF����'�}p����]�B�����P�������fo����H�6>{��2nyk��(�B����ƯEEyx_��S.wϻ���H���vK1��� ͹ `�I�3��f0ћ��t�*��u��w"t��(�s�K޺?�NR�{�d��w3�o�0��q��\Z���S��ygN�65$��Ӕ�B��Qa;�,c�]1%�q��0GVlO(c����>|÷3����!f{����4��SKС����[<�2�

ܞ�q=�9-aUf����T�y������q(�^III�|��N� �'�f�bcz{?eKt��oi�WeU�,yX�P��+�o	�'����V�����ѱ�9}�R��� ����(�r������!v�l~�,q�^uO_��Y�o��)�i]�#V�zλQ�f�:=�3T-5��Y��a9�ҝk�!�(�{��ŉIW#�R>�
]�����qŒM3��:���g��p%�����)����Ź���I�*��ML��$$)e��+|d� U��PC2L3Z/�wd�����K��rӧ&�Z���z��o޵�j�z
8Ew]@@��!Q�o��&��NܼF*�my}�]T� rz�qN*�	� ��{�s*�W�ِaD�����|�[����X�w�s,�Q��ɭ�)r��Tߗ�VK��ؼ����2tÄ�(mC�������@�S�z�� '<u���z��G�^�;:���Gtf�.Izl6�3Jص�W����rt��a���p�-S ������,c���)#��R+y����b ��6?C�'O�����A#?�2aq$9(���8�i	(�p�M̮����������z�����'I��sl��Q�8����(^��e����a{!8��5Y��3���01�9 �D ⺎����W+�gF��iCd��a0��1��&o�M�9�y+���H����{g���7��r��F�3�b��q��(Px�
��x�����9Z��-���'�a�*k�:5�L��*[w�I!L �b ����=�V�  ���#�x�'0
-D�#i��7����F(��v���g���>z{�~��)ߨ�����7�h�{9�s�<s�r��W�`����.��O0l�p�=I�w+P��$"���a+O���d7��="6�����l�c�E�;D���y��P �DE��uo�3^ش�bxм�̝�eK�w~d�(��DR�N��y}IQƘv:'�A���P	
�ő�7��	+U�Ui�2��^�� ��A3�e}��|B�M/�aP+����T�s���NK[��Uh� 6�#��S� �4��_w��(Y�c������"@qi�h�i�fǏ���r6/��	^�4��&���N�y�Wy�.N��EN��Q������L(:37�fT�a��S<"��o��x�h�ԫdD_��X2�%HMJ��\7�3�׃�j�m��*d�����iwN4	C߭d�0�6��w*�{۴Bm䭏v_�����@Mn�=�� vn�<r���Ɯ\�i�n����ya�4$ETC~Jd�V����<��>�F 6���\e�^���r/5�{�(�#/!�$o2�{�c�h�q�/�Z�!H�M%��D����nr�����&���	���`�c~��U��sT		m��4�-�5��j>���}V�����N�`�޴x�)�1�)��s�����ca4�D�IlO����6��HR��G�����.RV�'�Z�Z^u�a�Eh{�1���}��eW�B�{�H�Z�L��&��Ͼ^���>����&�KQ������\�J���c7�`�,%5�31�I1�.�D_<�S�]<K�gje?�o�,?^E�+��ݻR����"����3�X���.T����<9�$�Di�f���_��w-�2}>���UJӾYX��>Z���LV�F��(E�]���]@z�X��v�|2 V�{A��I�]'��	@���H�HHᷛ�U�-^Q޸ *� I���/_�5H;P =�t��ԏ�	��-c_W]���R1W�а���Ϫ-�i����c���B��V��1�oL�ῘY��6kˁ��mE�I@�HP4L�`�GX+_�r���ç�<�y?
S�/��D�<E�An�ә�����f�AO�TcK������UZf3���[긋IQC��s�.H���Q��p�:����/�qą��>EA�$�	:�x��D!��YqӮa����`%L5�F��??n;a�P"~e�=_��Kp��o]i��aF���P�U����/	u�%�4Z˺��,A2\Z���~?����mq����ns� ��,w�QV#���a���|۸ �hȭtWNƏ��1�Ԥ����qi�d�xc�I �������c/ul��]o�#Gf*}MKNҍ�LT/Z�h�����@��L�eݮ���b|.'���d��1 =z�i����=�ˎ�ᕆ��L�Kj�X��&T��~D������c���l�y4h���C�kJ���X�ơ��@;a}�J,�)4�^����֛	��Z�	�3����$
�.U���W�Q�^�vŜ��q�xad��h� �ܝD�����O�tN�^�u#D�4�Zp���# l�����sun.�<�g�y��j�,��G�+��pӺOb���&7�%Ϛ�W�|���*��?�pC����� �γh�%�>�jVX~��;tiIh)%��;X�.h�5	��/l��a���E<q�tyھ��$Oh{�44��c_j��GZ��\P*�Aď�Q������gZ*i�}P���f�C�̢����|�UUU�����4x]~�S)S�{KZ_t٫l
{7�'aO|>� u��^I^�׊��[�`$PT��n�����l���"�;J�Wږ82 �9V��F�#1���;Fe��HR־�d����'4�}�n�i=)q>^����b9k��U�O+�3ı�{C�ȝ��w��
��S��[��z(u�,OOH����
�$�{9pךl����L0��b�`X̕kQ���������X�H�Va���b�m��@�A;�3*�Vfo�d�C�:��A?j},q��|��&d�UU�U�`��l?`|S���{6:ƞE����-VW�\&��c�P6��A�<nhX}���ab��U 9�cD��J�8���D���̬��$�J���v���ʹH���p����Eʞ�n��ϼ��;Ih��n0Ğ�8bk�Yw������X��W{�N��Sv�q��'�So{�3r��h�i lM��-��Ų=QI֗o���v�8)�	jf2	k�2ʪF>�6aj[n,�����F>�!�4|\��[!�V�A���z���pzB1�>R��q��=	�H�엍H�R�ݓ1	��	���k)``�E�rQͮ�ױ �9����a�7E֯L���_]8p�*AC�7��Z;H�D��Z*844T� �'Wi�5��5�|��k�ٹd̕Dx�~�l��e�i+_��AB�h�A1&@�Dڡ4V�������S����/�6�~qΖV~�^M|Pp�,o▴<ZF�w�E^�����M��u}$��,��P��Ϲ�&E[�󭡑bp�a�J�,�橪�^A�(d[i��TTR���<q3�n�&���f�ÿ��`����IND=��u9�T��o�L�	��ш�@ٞ�-˵�]����^���t��}�}�\-|
B-�m���%K)�&?��I� wbO0�8w.y9mW�B���b���bo����(�3�]s��GR����?�q��	��������yP0C(��*���Z����Odh�4P����h6�!Ԅ;�����"t@Ϯ���3�N����7���Y�82:I��f`Ɇ"T�J�����9�~b�bN����Q8��
��� 8���v<�Z@u�I��>BN�=��;��Me�\q����[��K�?;���F%[���W����r��SgB��丯���:l�U�t9��<.��6��m�r���w�-�d[	������G�#�n|=cf��FjG(i���CS�LDU� �)���`�o������J�s3�s��qv�i��h���1��IǞ�I�r��i{��jkͷ,�0A�ˌ&�*�f�0,6�M����U�LP*0�A7�:Q���.��_I�2��~)�t�s,�ߐ�x��&�#��9�_�����R7�>H��`�W8�P�cd6kVtA�5Л#�*�:�M��d7�mk�����f�(r@霧5=�#���j��#�@2	��ƨ�r!j��A)!a�y�&�Nō�9 p�������!�N����$����d�+>��=a����>�k:9E�"�dw  >^��~���fa��n��͸;���O`TR�7�?����z�y�r�!k2��,{l=�u݅|��P�(Cu���F⶷���Xw>ǲw
e�a��S2m����Q+@.D�.���a��g}jg�X���B_��N��(���B�$����|�\���G���p(��1�.��L�/��������� j��E���_Ә�z�3{�R���P���
���;�m�!@���F�J����h��dQ�j}��-�������I��s���O��?�X����{��$y��c�#[F�YO�XQ��2�0CD	�`�����;�q������~�Cg�{V�V�˳������JWA �`��j�MxA��8>H9>+�0������?x���op�u���]J��d'�����@���~��}�.���l��z�>���F�Μ��e�P%@��B�C����꘮��BP<���$4���W}
̢G&}����/J"|��_�x�E�	z�_Wh~� �y=0��^��lSeR��wA�<�p��L0���S�y���^����g�6����\�3�[序�M]&w�f����(�	�i����=H�*]DE_�n�fBϷ��\�?y��9�9��f{��۵�A����k�-T��0[:��{UIqhq��0M���`(�I� A�
����w����&
�o�DÝxއq:䪴#���|�\��z����l`��KJPϥ�
���u]$����!�u�~n��!6��I4z� 8>#񇳒�12��%P�KO,w��υ

9�7�M}ӈ)p"��Bw�Yu������[?)�����m�L����N��Oh0*** �N��^�������J�֛�	�9��w�r��Ϗ��{���zEujK�(�ݝ+�k�������p�r���~-Z�?-5i��!�?!���]D_�;���C��>[���8XY |���jW�,3n�gj����7sZ4E������7݉�*�2��-`�8�]j��}Y��x�zGHV�6&$q�6�ؙ��#Q
[��9L��O�|N��/dM����·�֩�I����F�vWZ4��C�	��ŮN�]�(ե�O���RUG؇/�D��]�[e�6���$�x7�Lf(;H�X=���*I�-`��*�aVR��G�=iZ�;�|w�?1��6L���)gg��@�?��b-�b��>�޳��ݗ܏%�0��^5wv��Nr(��:$2��{հ��\�vg��z΅����?��i)w>�����ڰ�|@i��ɀ�0��B�U��	�5{������e�<��c���1!������X�j��b,��~A@�ʂN�p��f�M�k����`d$	�r��}�\1 �����ή�*�!�T���ff=��:䦆t���&+e�Jx��tN(�u�����#��cgf�y��:�K<��|�~Y~���v����ȉ�Q�WU1>pH�J܁_���1���X8�US�� �X���C��PH��8�α�i6��Tb�_����|.ZZ�D:�q�O��z��b�%V+ٝ�.�V�'��W6�k�.���*9��O����_Զ �1@@[�F���:x7����NF�A� �UCu6�� 8�(�k2�]�aD�1!��K���T��lKB�ƍt3�!��\q:���l���;�����v1m�G�	ᥞ�v��ȑ�u^N^�V�����o��"����HSi�^�n��~	Q���/e���j����ꞢL`����X<p�8�R��)s?6�v�2D6B*}��L��،%�$:�d��p�띙U^� 
ҍ�<��*�v����I���>�rQ����p���N:����d�
dɃ�P�8{|-4@?�g�j��#-�@ @ÿ܁|/����a��T�?M�+����EZ�����9�b��-�+��5�?<�S�?��1��?I�����첛���G#�?0�)x�`�y��ظc���D��"�{���/�Ҍ�1�kW �2R4��d�������(5R��ؾ�����([Cc<Hbf���.��z���894�(�ξ&Cz4]���K����y�X�;.��BC��t��Io��}%�-��Ȳk���E��2q��/�����ۨ�0{�-k5n��0]qq��3و�q��j/V���,�V�f��b�N��T����J��
3 �eɹ ��[^������P�H8fOj�H�m����L����a5��[O��~閻��<ĀJ���]��8M�^?��Q.���_��e�5` <�����i[&x��O�b��ֆ�i�F�P�4ʻCf�݆/%1�c5��
��8�)�i�A�	�45�g����Ė�I6C�?H���z�߾��{���~�ds5��v��t�1�E�ؘ�4����5p9�����m=���7t��rU��_�,�Ǘ�����f�[>16s�H��,�y����H�?C�[A�7' �T��b
��"�u }5�D��Bz��v&���#���P���U�ݹ��P%�"���^�(n������G:Yڹ�����v�~�S�"�"5��m���v�~�5H�@k"�9�m�+��8�㻡 m�S�z(5���D;Vm9n=J* �KШ�-+T��}���Bs鍃wgA�����-��<;fO�a�]�͸�+*[�ޢ�GR��i����1�@k89n�в#ا(�I��Z���*i��Af��������B�ȹ���:k]�PV23C�w��e��� ��Q��#*���y��& ����X
:��MЃ��"���"D����p>�y���p`l�=��E0~F��a��z�����������D6����&���?��1�3�V0b����,�~�,ʶ漰�U�a���(�?�J��nƈ�/e�lȸ���
ƃH� �Ig�p>���z7s��ɼv���|�\��������4+Ε)�.����������p79����.W� 7�G�,��k�;�ް��{�
 �lU�#��-�>�.93l�a�hP��^.H��^���?�#��$]�%Wl��0GL�x�I)Wf��A6��/*��9�L>����Ї��QX��Y�/��>n�WC�WSM�W��޺������:H�ӌvh�	��شh������~A
 d��OY\���&N�������{����(E��IXj��zx�SKIӚW����p"�6'�eϬ�^0x��6S�ө��|� �Q�z��b|�9�6!O\�m�1��Luc��,���h�@1#�H�T��6lЌ굲�ˤ�ډ��F��9��/@#P,� ���� G�Ǎ�1�wO:?+"�I�@��@���������ݾ�e�$OZ
��DgR����v8�!ϯ�+���y�s�G��:��ɍ����j}�,�$��8et��&儫�q���[�NȖč���0���luү��4U;|o�9H�4��	,��'�B�"��ű��M��S|ltX�t�l���~�(m���m���C'	<�bٷ�[Z�f`!�8A�y���m����A��]/I��p+d��Ԭ��rwK���G�K'䂚�T���!ʕ�| 
��N�+Bn��G�'�B_���S��sD�%��rH2c����ݐؐ�Q d,y�:��;��3��,�@,��L��8�v&���	��`���~���W����S�'o
�~/'�����4�9��ֽ�$J!�{��]b�m�K\����i�B�.s#����R��߿��&�3ҭ?�ʨ���������[�ѷ���Q7��a��v�G�Z��89�e`}���۳w�07	����Q�%�볹p*�����:9�R?N�D���nY�QO(5�ȤjG7�=��8�R�c~	�'Ӧ��m���l"��k��|%2l������R�߀ލg\�ٻ�5��8ٯ`|����Ex����q��ߎ��U\���Ϫ8L��D��R4����L쒦�Y1���������.F��2�O �z}Ϳ���5ے�\��離�g�ܥX�������x�D��|�ND [��`'�wR��Wf��[�$��?dqt�
���g�lReZ �&�,��>/a�*	K�r���o�<��sWA���o'�Bk��"��Ti%m)�y����,Կ]	9z��^��0�uiY�g����s_b���*�FD���/&��o��v�۫(i���"jo5Sן��^ŮWS�2I��mT~��cV��!�V��G.��p�S�Ϥ޷*[z6\g���T������Ij{$k�v����N��JK���T�Y���B���/_1q}K��%3c`�^����T-�� U�K�������U�6��0�ˌ����~=��/=b���oRk�M��V�DT,U���`O���p�/���_jrȀ�C��k@��B��a��@x��+v���K��"�΄�� ���҂���d*,���w�HOq��v�O�d�2�� ����
5�����n��{��P��bԼ4+ˎ�%��Ta=�k�I�7�z�>�T�@�*�0Ҍ���%Pd�j �&�G�%��H�8[�q�u+��'ԙ:φ�lH�W��&0HmA�` ]��Wk��M&���`V�tz�?�n��R��Wo�a�Gl{\,%�^���}��k>]�Z�6���b����Q�(��}
���?�%��k�@l^��y��F�D�>e�*�r��c�ʺ�~��8����K5y��Z;�f����O 
Wm\�?��މݝߙ[V٢��*#$����}b�pՀEP707����)�b� ��n�9�=��j�2Y�|�[<�Ð�n�N8d|I�e�L�^k`��wJZ;_S�^=*���.�đ�^x��Ħ%�4o���׾W?E�}�ò�.!KHǒ�
H#�tw�R"),)���"� ���!KKJw� -� _^������ܙ;sf�3�{�s�̽�B:��Ԡ�\��mC;�	�x�˂��3Í�@�&�HA{y�6��?7:�
 vp���ٜTZ���O6{�m�j�۝����8�:84쒒�W��>>^ys+IMk�����bk[v��}lU#zB;+ń�m�6��)�C�cl�c�&EJ�Hz��#�B��.�bą2ӱ)��Ķ��S�m���J���.}�"�Zp���
n2b1rU�<;O6T��d����t��;m���`o�o�D��(����]P)&e)��C�1�����9X�i:�k]���c	��-y\o�'_�ۮ����i@��7���fB���)ŵ����Fԥ��-�,�"%Mԥ����&�5_y���&$ro�m�e}v�PL{a!D�N\s\uӥj6���J��1����BO7�a*ժ���]%~�mQ
f(O�����Ƞf����p�Q�?�!�
��[n�X�䝀ʺ_ ����hg�I�K�~k'��z���r�狒� �d�J4�_<�X"�JȮ����7��"O��Ne��+�k���C��=� +Z����A��s�]��Z\$R�A�{6�	ɟz��)jGV���������ۓ92�!D�T�*�a�~4��odl���G�
vʹ3C\b(�qY�~%��3��!�Qgb����X.�Ck�)�@��"��b�w�]�Ȧ��}����d.�?2���:��S~lu38������[�aV.���1Ip�y�w~茅�~����$�AN,��Oy�Ȕ8!-g�2z+����.�u�.��h�l��K���0�%�����{;ND��?j�'�,��k�F+�u=WA\6\��8
Ca��ix�w�cn���l��V����P���9�)Hnq�_�j:mҖ$�40S9v,�a��>�>�3�/��O�T����$9#bB�K$+y�[UHϘ�=���ZMբ����i .�5>.3�Y�J�������(� �0%W�{G�N7���bɊ��>CJ�3r�LQ[X*vh�}X�s�[�d3�t��X'��в���ذG�Fl�T�Ϙ�xd�s�^{e����){n�\��&F�����^\J�Z�]�X6�y��(�}��6s�xT�7��Q���b8��J����|6V��sV��k~b d�]�Ȅ���/��\�x�3
H#(�5�)�_�ô26����ſK%����C����v��߱?� u!�	b����.[��&�[���DV֭���6l{/XC{��M奣���dߖ�ۡ�ٕ��.�6�`9��/$��a/����mj^z`�Iq�-�K;%��v�ʖzې?%qN�O=�t�!G�m�
�._�Hۼ-�D&)�F����s����G���M�SL�t͚>�|,��(fV�!(=��z�\��u�ٳ:�Z�e�ٿ� �H�~J�=U#U|w�^�3�����)�b}>�����EKH�O/H��h�Y@]���)3E��%��zIԅ��3Fd�F`N)�3�XӺL	+�az��i͏����ӾR�5�j0��x�����Ҕ,�j�8��������~]�uh�F��Kjd�s�"+����̨�������㣯~�*����B�a{e[��0�=6I_B"��gf8�ʲ��i�Gl�z�����f��������O�9b��[���	%u&驸I���ْO��.ĴU����'�~"Z������<�?��!q;#��?sJ����G��D�'��ͺ�1�q��<�HP8_�y
�kPl�Ǩץn����l��"S����G{L��@kH\#���g+�{��65��8�n��>�Vs*��m�� jy��d�~�{8�q9��*�φ����ƪ׮7)ǆ�v����]O�qbT�q�����p��Վ�k��'h eՓ��>>���N�@��3n�;�b��� ����ܵ��ע�e��/T�E{]��Q�#���oYij�*/���p{���߉
8S��s�N�!��i]z�.�7L�Z.�u��}�|�%��v�BL�ϏM� '0�$�J�V�S����+��.��w���W�iC�f&��8d{V���X!�%Q�� ��~��(� ؎�� �L�g/���|l}��BZ��c�b��Zr�ϑ_NEZv:x&�p�ޙ�;&�51ЪcE�}v��i�1G�|TL�o5%뽄���.$?�4�<P�ׅ�l�>d�9ك��Eh���Z�z�X�C�"��^�(��Oys��)�:Z��>��Z�/nvn��;�:g�~���Sc�89��R4����hI�-3��_}��G���0�<��}/�������f�i^�;�5���[999K�ľ㴽��.�(�\��p�N�K���Nۇ�+��i2��+����V��Hz ���։y!�]��T[�d�I�z�CZ���-��Ʒ(-���̃�����U��߉_���q9r�!$�4u��}����n~Oć�z9C�I:f�g�X��E-��g�ۆ2m�|Ay/�u�ln��C����� !/:�-��Y���UV.+5�K��d�u�I�w�x]����!ma��=��[^���� 0))�L�17ZF0� �/ӚN�f�����OH����Ȕ礲�tV���v���yZ�s�%Z�ǹPޚ��V	"޼o�٣�]]]���x������`}�z���b��ğU;#� ����7�Є�B��i��7��{���6�-�[9�g�}�jC:������\y��dWڒ�5��-�/@p��?���&ۮ�q��1oDC�d�?|b���f]����ϩ�lg�Z�#kNy8�[c�{t�>��!��񋭵������Mݫ�S�#�d�17֍����坬���ؒp kj�K���1N���J淢�c��g��{z�b"h[a��<������	Gই>� �O�$|����oޯε�~?a�:�{"4~�A&t��Ί��.��;>-ƞz-X=�����4}�� ��_P�o�g�+�E�m�^X��P�����w��ǒw����DƑ��#S�O|�
v���L-=?���F���M����t*��̔�Qz/�����Ɲ�}��h@�<��z���f� �E�I���|�]\��~�����]>�L9���R+
5�jLA���������*c�׵oHl�������ϵ���K�Q�JX8n݉8,)
��iܹ櫌Yr⛌�r��Q���7���3�`�o��
bGD�RK�����4��4�E���.�S�>_B���4��P���2�+*غ5�5آ�� ����B,W��|F+HS2ь)p��5hJ�K(�΅!.�?^=�΍b�t��}��Ol2�����]B䅊���"[���]�q�΋�Bﬂ��|���� dsu��B��������s�[����W�',��u�L���Ɗ���ȋ�<�0�J1{�~Ӧ�T�+cD���	���9�Ig|��tOꖨg�=7���^�����߿;���k� �t��V�d9bF+�:&�*�?z��9���Z]�]�Ҥ�Uk�A"�D1�y�:M�=$;��̋I����ؚ�$-쇋�A1bbb��JP%+��X\��Ӹ���@4)*��Ӥ���Ļ)sfY -?�7��,������;��oi	�yę#�ǹ0�D�Y��9/A�|�0R�d5����~P�������Ь#��Y��I@�_�~x@ve� �k=�E+�%�v�^t�%���_��1y���)�ʑ$˶�\����=Q�N�����=-� Z@͈V� '�M��9��Ț��������\(�B�Np5sޮ�|�;�B������[����T���ݓ��e�?gR��lݖ�=~�������k<F�b�lr�T'�9�=��R*ӆ�V�6:oRH�<��ǒ�s�3��O[�k�jg�w�������Y7��=e4o�gw��+��m4,I�z��
�g��c'��㻙z�6wL<���uq�k����KcTYW!��V Z��VQcn�L�"s��=:Y���Z�{�v�A�HIJ{K�~�(�{��^=�kf� �=�$�'q��,�E� =f���@G�EN�(�����T��%���s(���f��
�-�$0��ԤT��jrNH��V���Te?y�_^y�_$2|#�;�}f��K۫R�޹�=p��t��^�^����%�h}�"���Q�x�k뀕�HΓ_�H
&��w<+ׄ��323��HD�{��|۝���l~.
�Sy2��
}�-?�l(�ȡ�=���]�`�?�r�&�[EB3�\�`���'��߇����H!�0�����<���2b��)�u��氾q��ʪӞ�O��j�JP��ai�D�M�e�cc$����F���^��Qa�R����)��d-;�I[|r|*ͧ��?������DOM�a�������|��Ԁ��P+���HX=����N�%�:�����W�*��_m# +�)H�^Ő�κ�o��Ƒ���̎�ew��M'�K!Ui���/��}�'h�O�<p�$�'r�����"if����ʌ�S�ˀ��֠RzZ�`Ɖ�������� ��e�\�K��w���g��j8�t::�xS�)�.1")���ʵ��(NTt�{�T_�k�?ϛ���-��P����&y�џw�����V8���E��A(W�T�D��F�+��P`n�*���Z
xH~����"�]��=v����9�>�G.Is��;[��Y�f�xO���9��ܝ5�
��u�������>>2���A	�5g�H4�������E2%sI��ѿ�`��Ǌ�.:�{������_ZZ
F��͇�Sa�`��f
�}?~9��󕋜I�N��#��3����>e1�Fj�I-P}>���T�l��)h{k���1���l [h��Ù�k�0 � $���Q��JpjӉ�m��P���1�
1���oD;-�t���
������!� 7i��B���� ��r9�$��;�0�Op��2�ÍD�^O��K���E*�\��7U�������G���TQ��a�B:A���t�謵p���ƙ�~��q�w����=�v�E?n���l ~�̵�K��^c\��^�:x��wc]��������t1����<K��������{������z�)u�@�s��6��o�\y�c'�Ճ�� ����κ�����ُ���yr��~��Ҩ��W�cA�r�����'�6�U�E��C��,K��mM2+6��J��m��墦v�4ʕ�;f��Q- �8D�sJ��O�㽂�_|���>e_d=̈́S�3.��&p?��'�E�٫��z=�B���Bh ���r�M����=C���]K����5�3��Z��_*��4!ͪ��������C�6z��%���e/Pnj���d �{�O3��
(�ӳ���gm��˓�8;h/�P��{yl	�H�y[�r0���L��r�YwR�N.�;�V=E�{a@N�[��{�&9%���	*p���� ���+��˪9&��٧|ߝ�����������ɀb��֍���A�k������a�H��0��q|
yN�D�Y豐j�����B=�y~����>M�!G��K ,�*��4zF��l�Q~2�]G��tųW�g�+��oXP����՛���a�L��.e}�Ƿi�^����l���/a��n�M·X/{(6�`;���Izޓ���^��XK^�r�	;�����Y����"BV����K0�c��yM��sKII2�T��nz?!4(,��2I���*�R�.��K�����N$�`fJ"��c;s1��o;��Be�3u��F�z�y�"N5��	���e�	��,ēLeM���ZkY�J����[[?R$z�x�q'��mi�J"���
�4X�r��߿Ǘ�"��@�߳H0��3NV�90��U�8��O-+�aL���uX�l��~�NA�{���}�O����OZ��W���u��>�$|�d�ĆB+O̘u��AZH&(�93� ^ ��u���0����Ҫ457_']���R�ǐ/p�3�a��P{:^�nXʸd���}[�0����<L��evx]M��(�����_pje?�/on���_��ٱ;�x��@9�SU�e3aU����OC��Ab��D����.�_��=w�$A{ku<	k�2��/`0�g�`.}�cwe����e�y���x�~Y�f��wj���`&��\{l�a�:ݗ��}e-(e�<9�a��FiA�Ee�Mj]{ނrK�����g�X!�����ҕE���)���i�& F[���V��$����#��	ﲜ����v�s�W,p�z�G�������5��� _�#G�"5,�韩�z�BYU�ϵ�����Ԕ��ͧ���1go�׶ġ��i������*V��=K8�C�+j&��(&���\��N�q�KZ���9��V��SM�n�v鋙�bE����f��Xk��ȅJ��j9��'nA�T�.�G��h��]0��`���H<�,�\1!�����{�1W�J�� �U	�|�]�ݟoݾI!��%�N":���ğ�����vԻ���Q�ʨIo-O���ㅝ�=2PMx��;/���5���7T{�͕�ZY����$�jɬn:ۗبJ���8A���u��Ď;�<L�eQ�.s��K�o�W���mr �,�֐���#�-w�6ī+���H�ı{!� f���"�;\X7���9 ��_ݢ���-Nߌ������d��Z29�_��_���5�(���v�ֿ��$3jl/��n`�< �8��"�e*�Sj/v,�
�}g�5��;��\�o=`$_�����:���%$�_ΩG[��vvvRg��A+'''��Ք�y��iBN�&k�>V�H����ۡ�<.$o���L�mNS�4��|T��rMT����ghQ��\F^�&��S�Q��=g���[�T(�m9d{����L���f�������5�Շ�������w�g�iy�h��,W��١�W7��Wr&z�K��Ηt4 �V���'��������`4؎��<��	:�@M,U����=���}�E��4�(��_HS��r�`��W�6z�1�1U!�!krl.a9 �~c���t�J�]�$����V���ls- S$D��+��q�=<�j���l�p8t!B[}��;�س+�r��a\�Sk������ʡ�fj��TD]"}ǒ������Ynԍix��\ʟj�F�Sp:���w������}#˸}Fw����PP�0���k��g�|�䇦���o`rO����>+��>5-m}�ƮNU�G	�/<���t!���ޥ���58V,{E��C��Dd�&�H�WHgTG�\r�5Z�xxbNg2�\"��ٮz��6r��M�T1�-�1<ƙ<7�k��ip=\�-��4K�h���c�Q�����u�$�Z�3\�5Q4�`��2̓noę�M�ґ�B�9+�І:�糢I�z��͗&6d�m{��Qp�)F���H�3��_� �Js%y��,�ٰ���(�)�j���6nE����vu\>�E��&�(�?���쳴{�mo�������<�A$ �}-��@7������e�f���b[KC�p�u�-D�y(N�Y�<�(���n	!�щ�i�|�X=�rc�s���撬mbJz�lwp��G�o�e�,ޠ��<<�b��Jpއ��X�E�3��#9�k	C�aGG���"�w�~�:�G�Z_R�Ǔ.3*E�'vG]�'wg���{
,+Q(\&hR� �3[�3#.'��9_},����C* ������L��X�\�V
��������T >��2+ �;R�k�{kd8�
��	��K>��r�vWjp�xo��4�q!v���?������MpD?����������P.g�� PK   V��W�vh� `� /   images/d74878c5-97d0-42cc-abc5-9bd8c586a2df.png�zUO\�%Z���kq9+��R��
wwwwww;8)��]��;�d�?L��Nv�œ�%��� ��@� �,-%�m�����n� B�_\T$E�jg�N��Ƞ�ńՀ��=p�v����by�u}.|�ǥ�Dzh��YщScǐI)+	3�!�xu�(�� �S�aPZю�X\�����]�?��I�����}��u�fW�<��̰m�x���'�����_|�~/���H�eB���KzpBZ����#4��
<T�Yį��Qy�?��S��t������Sم�i��[�s��$��պ�v/�r���.Y��˳&��G�����Dԧe�9��ܽ�����&W+K���wU�6��*�#��iə|,/����/2�2�ɥ�:n:���-}��e�[^H��"��o���
$�3�Ɛ���[�����@�!���7w��9��%��YlC�Ah�5�r/BP}��Q�Ӷ�ʁH/i �%��7]T�Ǿ��� �3�C5Li�7!N��"?�O�w���.W��Ƶŏ�x�p>���VH��}�}[W~gO~��~s�;�>`��c����V��;W�z���Գ`#�'"ɖ�Y�r�:&>y��]��M�l�'tk�&�v���m��w�g�:	e�<JZ����%u��n�o����R��" �nz�I`�t"���S;����2����kI�l@�r�-�[q��%b����Ԭ��r$K� <�R����;e���t�zm��i�xX[���E���Է]�t4R�U�Ӆ���-c:�pź9oO�,Y��KV$��M���,�?3�7#�lcU=�%F�����,Q1�� #���%~��[�X�Z�Q�X'��?����I�5*i	PzA�[�8���x���C�6:8�a��xvc��k��Ne!�����9Ϥ��V_,
�	GU�S�Mt�F�2�����db�zN�Hf`J�O�Bw��g���5�����m(20�í�Tp6އ��a܍��!+W�q�/4�܀?J��nd���̯f���MvX�.��l��Yh�z[�������ja. �ߤ���ρ�^s��Y)c��Kg����B�]��)Fu݊E�"�g¸�X�h���x={z��Y����-��_*m��pRq��w �vΫ����}��ʜ���F�f�/K�!:ę����U��x6�l�2�&���*��Z��r�X�xE:*���b� �"�RJe�D�j~!�Nb�\�Td��*��v����Y�� D3�X��xJY�z�{�LaG{�4��c�H-�Nn"Uϳ���"��O���j�a�AtO���M�?C&�5�4��dǃ��������Gk����z��>/\+
6�R�C���@+Gt`ɣ�6x��3�3]��w����8/d�[yAh�L)ٿy�5.Q`��]��?ߜ}��l��{�;0a�BT��K���Q�8ɑ�c��z}��S��w�%�Ʊv�Aş�խ��m��$t�0�B��OPp�ϗC!;Ҹ��I�����z#-���(�À�W&�J2�|� ��k���tO����{�h�w���F[W�ݜ������MW���$�KϽ�T�G�UF���V_,�n�\
�lJ�r�zڦKOCb�40z�4a���e�1g/V~��r��+���	ή �k�\ʆ�w�ښ�M������h};�?C0�S��W*�����461ށ�q�����2�(?Z�ݾ.;!�<��N���Қ6��RS��7�}���/V�B��̬-�l�M���ի�i�|v���D�B�c�g��\Ĝ�%fݴ�\��&�2�
.)%-��i���"bq�] �m�q�M��V�EtueБ(�$�w��8�X;#?���ώuf?��U���0[�E�b͛l�*�^��>��/($$ԾM���
�4����0�eg���d�l�s�i29�J3��9����d&M+w���:T~��Ѻ�;Ӎ�*2L���EX�9�$�5�$f�����VI)fs�.º%
m��'o�H��'o(�w�'~iSYZ�}�A]s�H����3�6��Z o��gf��vr0�O�pK!`8��狝_�ӝ��-@x ��J2�|��s�x�E �c�i*'#k�������ƺ��e�����,����֊z2��w�V�_�Q���rxUn���.RrÒ:���;Ǆ� ����$����d�St�JǴ^ޏG���`"���� �崗�Y�t2D�2L��p�S��6���{�d�HF�2Bn�V2���5����~�N�+�Ѻ:�����`#"�A��OS'$�]X����^޽�.�`�����=��|Z���j��5��Ș��͙�c��|����1�$���|v-�rc6��.\7Y����&D�����5��z��%����?9�n�kg�.|8qA�P����Xդo�2���;�%��*+�Zw�;��r��$�Z�qu�C�5�c�-<RӉ"������C���B���Љ�A�b�'t˃��GZ$�jl�G�V;����v�-�RH��$�x��6��<���a��4l �VgT�DU�3˰�"�p_�^K���w2�8�#��*�IJVv�[B�B�|��A��W�M�fA���*V)�K)�q�)�Mn]��(�X�C���2U�G�?�Z3�24B�+� �K�ǚ�О6K�K�:�g�@�	�����?�/'� � /4hިHv����HR
(�w�M�	���xfS�Ya��w��vo9�l�hh���޺{�S�X�^`�3��X���0���\�3��&a�Z����cFPC_'��iI��c�#��%p&û�B$���]mr;�{�˃�%K���#z���̃y8O�������v�Z���u^A�&m7��ݮ��ܻ7Ыn�g�vp^�a,ƻ.>>�m.�0�r"�9,3V^n.#������_��o�2+��BV�ΎIc�ن���!� ل2|C��ڠ�;�`A�v
�G\�5�e0d�sz��'�G�ɾ
�-x(΅h���O��9V����N�,��@D���ʸ��vdQ��[m�l|p`�;�~&]O|�8�~��z�{N!t�t'� a�6O-f�d� f���Á�.;�ĸ![&©���J	��G�'��`�(�]��تp�S4�e;a���腝�0��ITT1�4��� �Ȫ=Rخ%5e���V��6��E_�C�Z�{�n�����}ͣ�����@�ΏDF�-� �k�
N["Iח��=�?�pa��]--faCVm��:�Tk�����U�n`�(d0C��+b@2��Bm5KXj��qjM�ۄ���"���Ā����"Z��W��bI��5Ty���˗����F\�3� !�{�V��JϢ�[�sn�No1Zi�Rs�[��j�ҥ���(<�T�ģ/$mQ�ۄ?�������f�'_uI���2�::�=G
#�bݼ+%p��LPI#�W]v�Q}��8�<J�7��=K	�0i�C�1�� ��^E�I��a�������� �-
Q�������~����I��/]袵�A5
�D��5��z�{��Є?1�S@�d���d
/�e�'��C�:���+�w=�42�3�`]�95��2�@�[:�s4��
�f��2c���t/�'��i��>S�X�	�ً� �l��f'=�8�iJh��bl�G�8�j����r�'�����f2�j.9_��B���P��M*Wh�s��j��K��	���,�2%c� Ͻ Ve�f�*�?�x�?3Xo8������3����$���uj�ЗL5%S��fԴ;�y��
0�j��-U���Dt�ȣma�F�1n��r��tɶ\UQh������뻰��%Z���=c$&�̊!M��R�U�DQ@�a2�;Z*�0b^Vuxx�Rbu��y�h�z�y�><7����h�	�|�FWWwecC,�l� NF��1L���9�-��Cg�v����e��~���2D�5��VOR
�]�As�����@Q�_\�EA8��g���Fp�2<�3��"�KVV���%T����+b��wO4M��
Ǟ@��J2���9*�B�� �׬C�e���>I
��A\x�>E��NA<&��@�$}��u��i���>/�i��9��?rI�Ye�l�o�,�Y
��mf����{�t	��GT
�Ϗ$r�tGF�ʣ�/ڦ��4Ԣ�N�Eq����[�P��ɲmqN����q��EN�W���z�A�ȯ���_Nh:u�-�i7�6�Fŭ�^%����~J���,�ĸ�|�!<#�z-n�%���zx����*�c<Z���?堮[C�C��r�hȍ7�ڿ�I�ĳ�S�(0�k���"DC�M���[���M�x*��w�m���,�!���l8�@;L��0�D��W����ӅKx� ��u*U�
&Ѿmɞ�v�Wg��9<��e.��,�����J
�8gJ4���rnS�\�ɗK �g��^|W��3gM�/�6��w��yL9¤,(HA�V��Ƥ�6LTs�l�K�X#�b�yM�ٌj*9��gӃ������ۆf�~[Zֈ?�_SU�r����O��:8L���o�3V��j}�,9jJ��P�5V"=ת���9���%��s(0�ˇ�>��9 `7��e?���p�c'�D��O޴�1���1!�l��F��8D
D�,Z�%�3R�tˁ�ʪ���	Xi�;ۙ��.8�q�?�m'(�2҃ㅩ�fp�g��k�vB�m>B����'T���sȦ)�q�|#�i��*H"JZ�T��J�_#�J��h��L>�V��)1҉��X�x���t�֔�/21��r
���aYU��
>�_�`� �8�<q4��1�����-��]jPЏ7d�`ۜ�1���i!���u�5�\�8�F��|�����9m�Ƒ����iݒ��j���� ������!��htT�uۍ���<<a^W=�ד���ב3ʤ��H�.(΢�
`W�v�F����8|������~�,�82<�4ڈ����m*jh��V�
�_Q��\r�.�s� ��k�q'o����R��8T��۲�Z�J�TJz���,�Ue;�W�מH���u�5���Sɡ��� ���͊�$���_5�����6g��Y��3Y���э斴 '&k�#�R����LN�\y�h����q��d�� �!�ܚ���ex�٠�2�y�/xuU[��묝Uj�R�����.]�7N0�#��ؤ÷e���6Wc�̓����*�f��(7�H�L&�m޾AB7���C,bف8��݆G�\#��yT(֦�:#�㙢{�te�`�߶�"@�����g�?���X�k�0����w��R>]~	ޝ�ɼ��R~����B�F���˦y�7��e"�F�	�XO�l�\�s�ks���4�j�4��U��"¥�#�=�R�}����G��[���A�n�T?��B|t�11�7c��׾&�\8�����m�֮c�N+B,�eݏI���<��C�Sz�"��%]����cޡ��n4IB��z�Q�ط�,3�H3�F��%)h���}����n��ĕ�'ѕ��]Ӊo=�JHR�/���C�r�sF�����7��>�ߑcX�P����-��
�L۲ �ݗÌx��
5v�pI#���n�l�I�sO'�xi*շ^\��+L≱ԇ�qy�ҷ�x�j{`a����`Qc�� :��S�1�7X�y���*��&m�X�o�p�f��K�aP<b-��a�^g�1��M!��pm��b�f���|\�0P��l�2��;�*mj/��nm�U{��TOM�CZ����q��:�t4�ZD�lf�p�]KE��B�-k��Em���h�\������HN��=� �вG:Ά�]��~��qa�+ʡ1��D�%��_�ٔ�K��#�Q8�t(l�d�4X��Gn��Ƞ�`u�%:I@�ؐ6#i�8jh]i�
6ONӯ��Kw�O���Ȼv����<�Uu:�튼S>�0a����T,靟@?���ֵsĩ��j�+.f&t�n˦�9�S��a�qy��߂�:vKD	IOx���� ��A8~�F0qs#@�;�������@��XoVV��Bdn���3�����J���w��7��{
d3�It������RCIc�P<�
�/�HLP��Ԥ����ꨌ�����{2#�Kt	�,
!�H���$�p���i�IR�%+�<9zG#��̯o���!<�u�Fx��>���JD� J�oB6�mێ^�o@�7����!"��Dϡ�[J�����/��������c�5x���<+�ceV�6�`�_U؅�ȍ�Q�o�o�g��eb��-��,�pu ~�x	������E��e��e�Ob��i�3�yi�����Z����`�_�/�.qj$odXa�h�%S%D������N�����JZ��
�":��
t�չb�������i�k��|����Rq�N��9fI���.<��Boy��`"l�����8�$�%kC�*ш�'Jh�"��TI!S��cVX�"\���~�}�ŕJiT!�"�ڨ��}76� ���p.A���H��j�Ă���J��*���FcI̟1����Ijf33Rm��촡���#u0$Ǽ(��I���q���L�4���̂x�'�j6�l�T�M-4$�j]s��5�ʸ�=����n�����he��߰BU�F��c�K��*S����+� ����y�odK���-�;�X�����L���V�/�"�vKv_�H�~̡j2\��PAm�l.�eG{��N���^��v�0�j�~�ֲ�$�������J�p��d#d���#���L5��ܸQ�� �C{�ZU��+x�t����H�7�%��i��C6j.���k��r�;zC�,���4�JN��b��F��_o��"E�$��˓�9 n+{4�J���̀G���$ry�t-����+^��햎�RM�Ğ;�ud!I
��kU�H�
������5�e����QCGo�n9b��/�PS�v��R��u�7#�O2��ӛ�F�$2��n�;��{�/4tx�qg�D�W�&OO,��_(�	�����#���9_��54o��	PN&�g�'��j	ߐ�zf�J8��р�{f�?��]���Od��Yd��g���}�Z�F\%��9�wM%zF�E!�A�߮�=w��]gP�Gn&��ݭ� �.G4�P�Sq<�z�� ����Y�#�w�MnR������h�k[�G�d�0Ե��pK��d��X#UQ��\v���k��E9���Py7ۺsTW�>�ֆ��#�ԭ�7��-NVE�6&�-G��.ɑ!��X����,Ǘ&��z��s�Kd>��U�|Wa���z��~�ǧ+����θΞ�X�7sf3G�I~7k�\ :�D�eP�rm����PD�V�6pY�u��(Q
DG�Va�qS� A��~��U�~�O�~d��h��}��j�}_�2�a�K�d��lt�iD�F�_�����T��}�������(l95U�����c�L��˸�5���	�g_�]���q�P��������nd� Q{�����I$�cJ�z���l���x���ӎ�p떐Fg�48+�����V��o���{�����Xp�73#��͕@��\;ڈ��sd*
GZ�͊����|�!�Aa`�ڴ(�Q�|�[������AY�%�z��a�@[U��:�ퟥ:P�
9��*N�#�Dr�M!F�,��Y�h�1�@S��J�c���R<�K�&�!-���/�c��H_�X�m"+=GX�x�](��:���L��A"U-PC�pN�AG�ūR���{�)G�P�H�g5S�m=+�5��� ���x3��7��3�9��J��0x�
Z��D�2j͡��TήqBX�b��d�����,�(�q? 6��n�5� �f��z�$ފj���L��z��H�9;:�}M�G�Y���G��af�\����	�X�F�DN )!6�Z-�u����PbWZ�)k��/V�8?V�&f�'��3^�݄~ZŏO!/����n�(�u�M�9+�d#�ȵ�b�t%>S�w�M��(�Ķ�8������+k��y��f��ȯ?3���[9�]T�(f@�
����U(%^��P�oJ,C����	��s<꺃������p�le�����4�H����i	졁�j������O=�?Z�<�(� B9��f�=�C3+k,���&�Ǳ}-�|�>)-%�&�D[L��Qy[��ΐ2V����5�j
��/�.ѥ?p�� 
~��Y-T;%!Dqw�u'��N�
k^�14��/���7R��9�����=�����	C��RىX��"g����'�0�*�&u<�53�9dHu��:Kr�A�:�����jٕ�H��"Z���W?b��.Y����zkhD�p��Ӛ�[�*s��R�[4�W�DZzZ�-*o1�౟�+(3%\��\6�"1T�&TFs�I�!S�k��R����r����E�7~>��ϏjEA�XFȆj��d�BI��_3Q�,7pU���N
1�90ڨV͑.�Y��ۯ�������R2��/`ȥ��n'y�S(dTS\�A��MK1�^	�l%kfpo����ЃDNdH�$��VF0]�y�s�\�pqV�i��ްR��q+h�'��vTh���&
����ྡྷ�gM���8ntKh�X����b�5&�[�	Ϭ����R���@y�fg���Z�Q�AS�
s��Ja�Ei}W^��$e�.K/��k�{��K_`[�F����R�O��0VV�o�&�^�/>?�ե(�X٢�i�.�#i�0�SÍ�_���3���CC��5�|y+h',VН5�`Z��pw�&h�ݿo���Ck�݋�WE��=N)f�^��x��#78/���qQ���	g�����MEO�s7Uq଑�G������}��k�{Â@7�ՅՊ�)�|�h��
ʾ�D�$�!.����'�;�5�\R?PF�ʟ���uf�c��ɻ(�t�K�g_��z�y&_z������$���H]�k����ѭ�McMx4�'����j�յ��;�z�W�uW����B�ý�vO`�r�Q�� 4�q���!Gg���}^	������,����~�5�Xm~�BhN�/���,�/���ù�!T�	���S�՞Ō��@�W �������i�̇P4,�t�KC��؅�����|T��jML{@*�we�ҊM�e��#���+PX�������Z鿱F\g��7�'��V탳�}<�l�X�^����S�w���D)���?\� ǆ�A���$���~s_Ys%o4)8`��P��_�~���4�R�7*?�7���&��5��FߔӞr'�=mz��L��� \�"����0��L]�m�L"ށ�X�jU���E��6ku��Y`p�C���X5V�x��<<��",)�V"7���$�ʰY� �
���{�zdb±���MM%DK��(%\��Yێ��cxvZ�F+��(:�c$�y��Gr�Ĝ�t7E�ӈʧ���STC����~��0��ص9�B��B˩x���lw
�7Y�5V�L�6՟F�X 0W�C�N��5���%2�6�&�u��|4r�h��M�L5�ғ�e|iD��L�ר�S�"y'���k����u���{HF�	
7���ɍ�{͍��?Hd�	�D1%����'��{i�$�jYx:m����]?�MJ<K|���ٖl��ۚ�CW��b�z�3 �b��4�����E��FZC�^�~`����6�_����o���!�h�ד���)��+����u��Y�P8�+�_F�Ѕ?���`������C����0�a]-���/���s���d��]rc�6�<���Z�$���y��(�yH��1�����p`�f�(/j��p�d�Z*����5頣c+�|�GC%'W��&�ۊ�k���j*���d~�<L��%=Ή_��}Ζ0�"�s/��i�Ti��"��6u���V�3Y��\! 7ä0����6�S1q�4��Fg7pAa�k�!
�U�ѣ�%�^a��t=v��W�Ik�`/f��xt)�r�k~�I�_,B���T���FR6&ALnd�50w@=NY$�eɲ���I�����cQ�'�Ln`W���(\7���[e��[+���/�����VϤE�A���+yJ>Z&k����M��1>�� n5�}�g�d"h��SW�Rp��m�z���~�*�5Ud��;d���4Ǜ{���.�.�̀4��ڶt�"�Mz5���q�j��m&ln�f�OɘP�~ZHu�_z�ݠ�&�g|�����]m�)J>6�$�}2u�.\�^O���*�z�(�����l��q�l�}�;�:�����T�a�`{2`pwt�N���5釐�|[�jv��بF�:�Z��~�đK�h/����K���W�7��(�8Y��4���T1�3��c���|��R�sx���uK!�.ϙY�o⤚���PC~��K��l@���cE�&(q�=6��C�������?L�H׮�S���E3���_�.�s����O2S��;���NMP�N�ܶ�qT�5��8��K�@���%�B��:<�k��	�{"�Ѫ�k0�k�����p
�C��6���,��w7ȝLI�v 2�(ˎ�ݥ8҈v�X{mh^
ѵ"��r��N����+b�` �T�˒���HW��"7�-�1 W;���=?�
��]	��������������o�^���7��]���&�dZ�"Ő�:�e+�^s� s+'[K'�~��.�֜�4`���믢բ�5�״:�ѝ�@�����St嘼�����:?�ˎ8C�s�ij:~���U���:����jAtL֢�o5��T��Yr"O�dr��|�?z�ݐ��B���z���j~�Dh�&�{����RѺ�tnM,*���N<a��4�v������0��R�uW�y��)uc���%eyp��zb����#�f�_� +M�s[��.���K#�F�U����fUzbդj�Ld�*��2����q�	W�z�4��(xUA��e�ȂbKS��K}~��Z��a�Q�CF����wքO�(��̊d�Ǔ8����`�.K�*9o��39��1�pf�I4��F�!?ڕ+���kZ.�d5x,._R=L1*Ui]Nû��֐N���
����ݡ��KO�_�Rn8�����ҳOe��Zͫ�K����4B�JoG��sF�}�V]�T|Yh��`��4'e�_���W�^h6��!�p��r��2r�ӌ��-<���n�����}z%^&�=��z9�j�[�3���7/�b���wIpo�q���Y�Ƹ�G��Te�(��|�?��#%I����w%���4�N2���~t�y�e��u���b{��Eõpb�E\�ߛ`d�2�F��f����QNAd9,���S47G���HU�I��������Y -��`����z�b6�:Ka��fV5\�T}咛��黃y;��0�]�c�Ǧ0-t������u�ֿI�~lz�ܫ5�g�%z�b3]
⏦jޤ�������f}�`�����9
!���z+�,�������/ܴ{� dt�>������]y����)��:��%��?��|>��C�@��,~�2φ-�*�B��\������Ⱦ�N�z���E��ՆDm~ *���)U�CB[�0��[ԋ��<��eN�c$
�J�wu�r��k'rM�9�M�
�Q�+�#�X�[���Ԩ�W&_�=��#ͭw�lU���I�Rȿ���Q�1/�Pi�.�e����l�ɎA~ ̙����X.>���`�zk¾�W��3�nPΈ�TK;��Ң-���a|��A�&,�˧�.L[Le��f[[^׀���s�v��iD�
q����jJYL�M䥳=y�W�l�K�B�F<
���|!���w�>������7���W�T��_J)�bk��b�I�(7��}�׫�E(q[�6Μ��:-�C@�z�'��a�O�e��.-�u�
cO�/�8�?5�5�58���ۏ��8u����3y�dƏ�=��,헹��o~h�����\)i�it6{$��o]t7IA�K�Ύj���j�"����.@�۶�dx�q�Vi���MN��vU1���pd�W�Y�4�6��y�'''˗	CT�L�`�GUĚ[Z",��ѓ,}D��h��r����#�[߯�(�gL��q�	�E%K�
�쀅�������4�vF�n�y�c����$f��n��j�l���@]�A8%GCռ�^P�ww�����fJ��/��M$jdb�ѷ��c���,��o�9;-/-!�%WP�~�W��ɇ^����sg>��ݜ�U���	Rk�XPXu9��Xf�:-�k���3���t9�nxZ
�s{!}��C:�Ak@��ѺH'm� ���it��sJr�S~�D:�\R%�3Fb���$Fn0j�a��������m�7�'��8������1���dOwG�i�
�DlRA�L��veJ�F�7���8��pi�.�����,��`��g�!9/.;rͶ�ך�:#���xZ�e�0�2T�u��ʿ\j~" �S�����߽��Ǌ��˖�/����+�^�@WCkCl��h����Tl�������n��F��Ô!��Rl���*Tݿ\�(�^���oiLI	���~g[�	j���p�f;�7mNT={��z:L*�9��yT?|������r���h5*O��2	�?6�7ky���-��S�jT��4���U����S��L����#��)ᚯ�7=���|~�Osć���	�;4���G�i/���U��W�ڃn`�����EK����E b��7��y��X��i���;7q�x�6sW�&���e���2��?��7}���/����L�$��գ4��f��|f</�@ߺbI��lIS���v("�3 ���߷{N�,����ɲb��k.i�[y�i��x�mJU�9/=�����ޕ�?��!��ݐ���t-b��	�+�!�	��cD���Ά�������&kuD=� �Q�V�>\�Q��n���D�Ig��w�`ϑ������e
�"��c;{�{<�������Տ�\-�O�Wq�<���b��T�Uj��j�H^OS�Y��nvLɁha��#"b��֏6H�AɨFk|�z	��?����J�v�������qw*-� $�7�9o���F'))?��f37#�F_�W�>��'8�'�O�x�����9��Y�A�z�d�$]�"�սѣ�މ�g�y!���/}���}�+J�\*/��C, ⧍��t��!G��%k����}�^=7]�Z4�6�B0q�T�U��9�c��ʐ�q�.	mz���sBL�`�D
w[������V���H�Q^Ĳ���q��{G�>��*��q�S;��'+��>BT����	֗�N�ڦ���R��4�[�#5�C�vr_l�����b"���r���ݍ1��*+n��(1�#����a��_"���7�;]�py�2��^�P�)��Qɳ�Ž�U�d1�J��S���xXԵ�7g.��h�3v9H*�),�׸��z���G�C��8����4 �y�w��@���aȏ�>#c����W���>�r5/�O&�Q��Ņ��zwH����G��6��I���\\����#��܎���������-����.�#�y�4U�V�y ֜{��k�%����/5��������h߮Xx���Vz��+��`��rL�e����q4\�9���2�O0�H8ЄI}Q��{��D*C�$G��_���B����/#��������lc���W��q�O8EC�������<F�S�'�ѳ���Ѫ7�W��=��&5'8��(�q��M��(�7Z>��8�n�����2v8����X�2$��s8��T�#wyT��D�ܗEڈN�;_ؠ��*x�v�qy�������z��
�_��+��[����c�n�%s�o����7�={��}Ki�� pR���ĵ���濹~2�0BږFϔ�~�͍��?�>v_Bk��S��"��H�'Y*�چ�u�:x���W�Wࡀ��|���ǀ�`�D	p�� ������Zk#�W��p�e�i��i��v1���OT<+)GZ��?�=3�Qp�%6����*�
y���ۛ4��S�����hi#��4r��×׫�&�	���
�	*����8���l����x���G�{��^0�?��b�f2��������"(��Z�T�KT�҆`�c�Iz�օ����%RȒg}3ŕB�#�FJPG��7��ܦ�џCQ����^��9r��<�@(���{5}�|� k���$����p�B%Gg:��l�ⶖ�<��Z`��h[a�ffJ֑���gn�<}.�ݔ����d��:�Pf�;�K+BA�G9��s�95��"fA���M�u�V���[�0�+:ҎP�H���Ӯ�o(�_fx���2A�$�t���^O9��ݍ!^O�v��E�-��#˽0���DM���	`X�R-`y\�����g����t5q�)��!��]��]W�=3aV�"??3f�݄ ��$��d�8���@��w*�W|�);S�D�:���P��5<�?�&��P��s1a0̈́��*~!KV�f�����\qz)]��/��9\�s�����E(�M�!�&-���&[P{y��9��}w�s�{v��W���\��H�i�0u1x�d�}݈R�Z��icD˿�^Ml �IS�
���fv�/�hE*6�-z��Y�������C!֖,ҾG��D�P��i��C��X��'ix�$��9J�"l�	1
#���m8v�tz[IxŸls�-!�"���I��M�&t���`�a~VQ�<la�fXR��e�~Q����镮�^�^�gK��Y�K��罢����譤X+�cD߶�����2)�{��xzDA���0�hh��\�p�ʥ���ͅ����g���+17�A���`q�Mq^:����������Y����͛�O��������f��ָ�]�����������ޫ�sd.DnS,<�x>�Wl���p��I�7k��9r�GZ^���EL"HH�2yU�U�-q�4�~zD�	٠��Ϭ7a�}<��SV���\��11_���۽o��?=DH]^�wFw�9r������y7/��	�aӉAH�O�7� ,^��q$8�g|�,�J�N��M_G���ސ�@>�u-g���es��Mƥ)�S�$LT�';��Y�Q�cj�tT�uI�N`��]�m��e��R#b�!��9:�������Q��5�N���޴5$8��˖#C��3�^���m1ӃZӭ-��'݂�;V�z��={#����t�e���/�����z���wq�n��r�>F2�{�%kŒN��c��}�>4o��<8W�ıh.�?�᩸�E��~;�*Hd��,|���}g�'�Cr:wy^l��n�F)��W����b`����v����#4���׽촊$�O8CLjE]�O�-����=��t@��%�SL؆M�vCr��?o�ύ|C�c ��Bޛ�ۛ���'�<K�"�O��2�{���Q:��]�δ�'�/�=���"��Ё-^wJ�4��ԇ-+iR欨wP��>8��PM��Kɪp1}�����	Z$���y*ݾ8�1�>��؋��7�X�G�f�N��n���Bc2u���}��~��NG����%��p�w��$^�vb~7!�='����?�{��m��hk�JzY�,o�"������H���ů�9F��6���|��}Y��K�͋yH�yb�_W��4fTB8{��o�h?ϛXm�"%��SE����TPnJ
�3�YA��SYk��>Y&)�*y�QoY0�͝�負j{��6&�G��W�S���cY}!v9~hC(	�6�όn ���L�a�D��y6��V��˃������
��5��=3�Re����<��nD�������(�M�i��Q>��	�D��)$@�!��ř��k�^7U~����D����é��X���[�ц�[=p�zw�NՇ8�{�W��1��CF�p�a������t�UW�JʶY��st~��	s�o��P;v��\㦬je[�4*T�T5��Q�����C,�k|n��B��p6����{�M�0`��HH�(`�o�Ѻ�~0�*���k���N��A���|�_�mw������;�d��S(4�w�︳>ȍ?���� �E�C`�w��w�� 8�A��*Y{M��*��q�T�0��/�3@̿��q߶�	z�k)$���U�t򞢧�&Dl�tIxofܮv����Ԋ�bzْӚ�RMb��H�$q��BZ]L��&Oa㽢*��Hr��X���l���#u� ����b��]�< ���ţs��2�M�!�ٹ�?x�{p�u_��}�å�x�o�c��<:����^��kpxy��,i\Q6�%��jJ��s��4���Was}Ip]�A��>
*�JEE~�K��~��H�*��!��	k��Ih�B���\�׿�����kaV��K^�K�|�f�i��ڏ���mPAC6'�^`��h���CxN��S��?[�+�G���=xSB��E]�Ʒo¯��{эr	xHcV�U��\*؞��'	9�gA�Z�P�CG{s\����F2�A�G�4��W>e�I�@ᡗ����+�|d<�~"�/U�"�����8�x�/��Xc�o�^0��
W�����=3x�{ފ����Y=�OW`L��T<=�9SS���� �u�-PG�Lz�<�l����yO{^� O�R,���</��i�$��38t��w������
D9$�|�s�`�x��/�����r���� Y�38r�0��7О]�8Q��y*����ā�M�,���=��D�nU},�]|����ݬ!���&fg���azj'����_�>������a�CTCv�ca�.D�ԓwH�S�'��rL����VV�p�Y����ߊO�K�>�s�?�Ԫ�#s�r���=��ؽ0��s:�𚫡L����j;�q�ͷ�s_�2��4��v�w#�7Ǩ�v������X���׼�x�%gbm�t[g�bE���D�jxASHا?w-��� ����<�9W�wށ����ҫ������H��w������n�T�����}G���t������}�tԏ{=<�iW��\���҈ti�:�-d�XH�8�Ts_���?�����+G�+o��	��`.�����Dz�h)`{�_9�t�^[��8���`��"/
��u�>]bۙ��"K��Y����o�e�^������Е�2m;�|b��!���W^�*\��K�k�\�Po�HO<Ε��6VWW�~s�;���;�#�7p��p�=ǰg��t�?�!}d�輳q�ݷ!`u��g7��ɾ�	�� ���Q�Qi<yV$�-*�ҳ�( �wf�ZE{���@�IՓ��6%�M'��}�������_�⏖��c9��߳�0%���9x�o|���8�"�4���PɈ�1���<���Ϲ��ӏ���.��������1���#>��a�Q)<)n����R���I� ʻ|�%n�t�1'_�d�jG������ ����L�^'�>���'���H�B�&���_L�u�їi+����cN{�`Q���+���*�%|�JڐP�PM���� ��t�����y���Nރw��\���������,Ӈ��zߪz+Ǯ��=ӓ�$#"�d
�aqŀHte�+" Ie�i�a��a�����9U�9|\��5�����s��;�uΜ�����繞���S�����+�+�L��"�Պx�)6;����`6�����4�4�Y&�R&��?q�>�ti��t��~3s�QO*W�$w�?�{��z;��������A���]1��M��u�Ν���B0��
���ŧ�d�L��O_�Ԛ���EVmh�ZA.��e��?�|�1>2�]�4��q:�x�#��3/�����#DI�2Y�8�#Dbl[ЇZ%��9���K1:��!��>ik���)���������+���*l�6d�9XL*�f3���<�����嫯���0�V�}��*�٢;� �bY|�+�"Ul ��A�����)�<��]>��-�#>3	���Z]Z�V3�T<Cux�Y�����K5���c.^�#+��Mh��U.��98��'
��4V��$���dsоÂ@������{Rٚ�H
�6[Sz��pډ�/};wl���ť�aE4A�TA[G'2����r�w�*PfF�ho-�b��7�����MȤ�P�Ee2��葪�t&'F�K��?�Ͽ�*� JM�)��.�7�s����<�6U�Y��X�Hg280|�X}#��[o��t��/�T�'l
,�>*�4ڼv����a��W�`�Xomۊ�y�z�_x	^۶O��IZ�* ��Z�j-����^�i�v �3è4˰�58�n��n�43�2N��Ͼ���ۈ���l���Ʉ3�9����LJ*7m�N��O�e�D�H�@���C"���O\���I�R9�%Kbj|J��e�����HE�p�-7ḣ���E�GO4.05�*����A% �����K-�������p	�D=��f�U�JE�z��O�`ppX�2v29�M��f�1��% }Bv~V�"�b� �+����Ypɥ��އx<"���s!�s0i�����|�+���߃�k��I��_'��sp84�Y�w��A������?�D&�EKWO��Y�N,T'�	nfSV/��=��� �S�Cf�Y��2���&ǹ%�*�2���J��r�o�g�����R]�	��`"���x�s�_�b�M�|�r���E����=a��1���x�������r([_MJ�Q�b��@�j�Wt᪫�#��q�Fl��&���(�<N��Y�J�V�8!K>����[o�%en^�����!�I�i�.�&,]���Edȕ�a�`2���WX��Pd4b���R�T��!��yr~�ԮC=���
	=�Z�1��,��$~�V�}���������J]"n���XTi#P�W�&�$؆���}L��b��=X�|��̜r���0�B�B	�~������0[Pj4�t�0�!f��|���e8��c�<1���u���t�ֳ����÷p�T�Zt2���F1��G��Q,��c��>�S����@��cG���#'Csz126�+�����ɯ1[4���ZU�7�8>{�'p�E����ZL���e��'6=�������܊d��B�w��l>�$�d363�8�$\}��L��a5�E����<U=\�N�.�T?|��m�(I�6
�9���J�s��.����E&ഛeb�d@��d�����ŗ��]Ĳ%(� �X1А�b� 趠�̓[n�6�ٔ���E�>�h��f��=���w�m���X�$���3��NM������g�x,RɈ���4��$W�m�J�p;^�H����G�E&/=S��'�}���W��o|���Lό#D�QUA{g���|����r�R9jMXliQ�4��dH5�5�v�(f�P)&�
lV�R��]�,P�%,^�����x��-�w��H>E4�
�a�?���S�RiI�齵s�nd29Bmp�=��n�	���
f;���4B��p�L8��c���X�d	�� ���p?��ߋd:���?k�:
������+���On�]lrq�ԋp(E|���qĪ~L��IS``K٤����*�V3"�.�?�3�4�g��������NC4�k[ސ���f��QR�"����пd	4
#
�t�[z\_f�	d�)�;b%&FG�0�8\HNO���N�wѨ��/&`R갻(*����h4j7�Zh�?��ؾ}+���?��s�@<2%���_-�/����*�Z�n������M����܌T��Ϧ���/�c�X�̛t�qP&�
E[�4C.�]�x�B�v�͈DfDQ�򁥂���`�vy�n��O?�ˊ+>s%������鲉����5�f28��S�4Z14:�]{����6mޅ���fW�0ȵ+
۳s,�9�4��b>奷�6o8�/�b��e>Dk����I
xl(t�}&���My����:���yԑ?����g0��W�?���_�����^>�_=򫚣{]SuI&]�\��4# t���9	�j'��4	�1l~s�yg7�V-]��"��瓀����9�R���z_����� :;;�͚1>\��f�"o��+��b\1��{;��'�ZNb�a�R� @'�]W7->١�Fވ����,�K6o.�{X���Q*���`�I�U�Й�V���G����CH5��g���سg�������(�
0Jխ�[���?!]��dhb.��j5�n��Nj����o��k��f2�j�8��u��X"բ���Ï=�ǟ��^L�b��6m�XAG��r+-º5+��������+���8����969����:<���Ū!��J4���@jv~�C8��ㄟA�*F�0���u��/���Ex慍���?C[{�'g`��(0]���A�����_��χ���y��d*.ו+�G�d�����܂h�(�M��!��B&s�
I�~�Q��ӗ"��fѣ��nwz�v��^+����(����1�Ȣ��D:Oo#fC�M�\*\f����J��xə�Մ4\���D0D�^÷o��o}Վ���x�R�{v� �����N:�t�}�(�Y,��V��sz���q��.��S�B$桭�C�uk7���r�]ai_S�<;3��'�/�L߸�;88=�t�,VM��B���'ׅ�b���$�լx���q'�-+��%��/��w3v�E����B��˪E�u�p��7©���
��wb&���q�TE"Q1.%������dM&EX݀I��d6��X�ש�K��,���ѨT�=�,��{Q(�hG�]��[~�c�ص6w���z�4E�Om��PJ��U����09y�z��M��%�+�}�ٗ�y�u�)x�����+���۠q!�4�ae%�X���{�r��Y���n�OK��nu���x*oȇl*�ngL�:��(��|��?F{Ь��T����|P�o2+����n������kW�������0�%v��S�s�#���L����8�g��RQ����%���OEz[�yi���O�E)�6��633�B.+����z#V�Y�d2.ti��"�&|0	r�ؾ�-<���غu#>�����H̔���D/�*�R�V�=�don{w��w(PT�Рj��n�^�4�\��0�����I`<;�e/�y/Kɘ���GQ��`r<�����\��ML��oc�F��\�����Th��<���Gu�/>�я�����]X�?�����������;����ŭ��%��)lE��`���x)K	C��Q,eu�&ۉ��:,ZżT�����Y�� ��:��c�1=N��lQr�S����&�31�c�5W՜Jt_1r��Z�����!Fy&E�D��9p�l�u�1�Zѵ2%�+�o<褼����~�/[�lU���T��j�Q� V��RR�Yl��v�Cx���f����=������+���pz�󆄃��177#Ys/n~F�T�f�Q��%(���D����5������E�������_��K/���{p?:bxv
����\���-�r*�(Ԭ�[ԋ��~�]>QFq�E�mh�b�a���ظi3�:�����B��D���炎�s#8b�r�v� ���h!�8%�]Ni9p����Ͽ�;����,�u���9dJ%x�~x\.4*�݇E���w���a��2�J�:s �4�����Dd
�˖c��}px��O�Fq���M!���e�~�ȴL&��n?��6�61Sn��>Dcq<��'P3���и(/g��Jy,�	
8)&��K/�Iҵ���@0��]�w������`hr�7 հZ]A�-�R;6m�?~�b�~�Q��k��*�ZKLYP�bEWg/��x>�(���4(�ç�mh�����|�:=!�+E�Rq9�իVb�%�}`�s�02A�~\�����4j5��'���W������t�y.������Ũ��YT������,��V���
�F��$�,ďn�~�^�W��2��p��q�f��O�X�e��C#�/B�\0��R=�M"�L^-�7ވO8�\QE��=��m(�s�l��7�s��N���@"U�jrIԙJ ^+�e��_���W`rjF�*٨t�ؔ����l��D$��~�S��163��HT@�����s��]i@m4�ؐ�D����ty����G$�G�\;�O:�d�RI�ϰ�U���@a�Q�*����>'-�
0[u~R��\H�?���xD���+8��c%-!�NH|۸�\Z*�l�3�H��I���)LNF015�s�4�Nϋ�T�4?���V[���U�8�G�IPF��F�r9D�MS�K/� ��!LM��N�tׯ3*�,�cl���Dd.�'"��O(|�����d�*Rc�.}�
�:֮?�	O<�<�Fg�e�nT�53�g�:�D%�ıG�]ۥ=�2��J ���p���r����,Wv5,L)!�����mN��p����R&ubhpX����O�Z�B��(Jk�{�ؚ5k�����X�oEI�ܡ�N��ـ�@�����'��������GG�a��ȝUch-}��%���0�)���a/clr>s����`��0��|C�+yTT�ɼ�[I��$��8��:����yr.t4-.Z�j�gt��O�b��?���/c��%�g��
o��M�=��d1n��ӄ� �~*
�#8�?�+!�J�C�|�$M�$��zF
�=D�K�l��iZ-î����h�28q�*���R�!�����~_X���2cll���7<�{��g�.���i؊����aL�aQ{�g�t����I����w(���n<��G165������XX��n�g�1��#���.��,BG�v�&����iX5��Kv��>	k ��h����
p38z�*XN��]�k؝~�Z�1_U���	毻v��;0��">opI��b.���ņ\4�훶�^d��J���?�M��+�db�\�~�lX�^�M�upT��d�{��2�76�C����S�
Vt��(5
��lh��b��r%Ŋ'_ވ��(��24�
�f��\D>��lX�v�Ua%�,i����m^���5��Ï�l4"S����l.7�+fzn�"�8v�2��,X���=�rI��"����@_g7�ڵ[�ٍT���x�r�LnՌ����a�+��w`��H�38묳��݁�}{;��(��Q����8��p Ŏ�a!;G#QE�w��O��1,X"��Y�� ��b��A��'��"�Na.�Tb�F3��T�Հ�������v.��B�>1������]Ӱc����������De^�F �{Ӯ�r��G'�ሣпh	��LV�L��r	�3#�z�	�ׁ^{Ǟ�A�B�̥Qa��YEOЋ��A|�����k��KO,�����"�U� ���q(>n��n�32&�V���z�	��~�Ϳ�5��D.�B1���G�l��ɹ�F*��Ҷ�F�6�Ţ�T6���+�[��s��������f�z�@sZP.���+ƙ�{߃���3?���6��$bs�ڶ�U�9}�\��5E�����q���f�]��LC���-H�x>����)i�	 ��    IDATk�jGnA
��L&�ˎ�������W㳟��9�T�J ��?�� >�����G�Ú�+�l�2q��������1
��/�s/o�+�m���,,���H��p�"i�&����rx��'`|d��TJ��E2C�u�����j���&�l�Ì�"o��t��l�.]�T�k����)������AYdF�����q��>U5׎;�ـ��m���x�Rux�)��RW���$TM��UiZK�Ҩ�MMk#�N�N��T*Ս|m�RQfs�^/�v{�Ag2&_�[�'�F��.Ws9S��l�G��hԋ�f�b�4�0�J�����4�ah�s
���5�:M������&���z�D����Z12zt���\�Z�9��܆�_����1������ͳhm�A������6��4����(�g0���݁��4E�00����b�RFz5���k�߿o�p�	�W�D��J+^���Rf��۪�	��]����3���V�jW�� ��A�]�5s�׍`uR=�Ѹb20̻�O$ �Wڇ�y�1Nz>�|�p�$��Υ<��z.�~�Q8a�Z��0IUВe�������

��	x�Nl{{'���,]�-C��p@�e�i�6�q(%����փ�`���M�A�sM8x� �ٳ��Q���r�\#���b϶-8���$j�iw�+<���x�!Q�ky4�i�mF�*y���p�����Ř˕��ghfQ�ۏ֯A��}���tv��
��g[�16n��c��xu�v<������a*G"2�ٌN�s#cX��3~G�э@�B�N�J��P���0�;�����g6���͌Y&.0�\�5�F�ڀ�PŢ��l������`CG��zn/�1�F<��M��Ʈ�����Uh&l�p��R��jvlX��p���駖e�t�۹�
�.�3/��{�!W�#N�����6ܦ&6,]����y���FA��<^�R�C}&��={1�Ic_lV����l�5[��b@)]��7���h�Ca�٦!S����R+�g�ú#V���~[�F���Ͱrl@)�����M�ؼ�SQ	F����wc�X�܏l&!�.�Ê��2�}pf3Idyx�v�L��NX�F�|�Ix��g���K�![��	Xc�9����^D�T��|��J/.���*;��V-^�O⓸�a��ې� ��4�.��ls3;q�E@��NOO![����������^xUvoق�N;������d�PE�X;��M*�ۇ��؎m�)��+Uᴻ�d���DC�� 6=�*2�I�bI���>�Q�v�iȤ���/���l5��Q�����ֱdɑ�OG`*�a{Wp@sc��  ���#�z��4� 1
��b������������1�z�ih�]��$E�^)t�:�Wv%Lp����x}�V�wt!2G�.�� �@��	�K�}�X��gP�.��:M�s�m�J�d�BZ�(����v|�+��e�*+Jt�V�#�
��� `�1��=X�n5V,_.9�m�����)����</��&^z�M�?8�/��hRڪ���{Z.d%2��������#�bjL%� ���SRh��J��b�8.����U��!z�#@����6M���"R񔼗�E~;+�6�Q,��͆!U�5Vkը�����y�:�6�5�N
��7�Z�ڴ;�uL��]�dR<Y�)��Q�������V�J,�uvu��O��}b|t���x�����Z�f�UEI�2�Q�4�=߬Ռ&��D$��LuEU�&��>$UU��z��(JU1�r�јI�Ӿj�����Zk�5��X7�u�jm4�ED�(��X�F��o�~M�M�(Ĉu�d��mZY�9l�b6Vmk����d�9���A����=a7���;TG�Z*��$�J['�\x2�#ظ�yd9L�#(20W@#W�R*I�US�y�a�<L��:�-B��o����/i;�Z�K8�T�Zٕ������RŃ��t�'	J���b��$����@}�juqK&kE.�յ�m-'x>x��F���M��(T�.j���L�]��s�]��}x�����wvb�E���Cgg/��61�c������c�~�𓟣k�잜B��\.��e�E�����-�O>�ݽ��Z�z]W�9�����R����K/��?<���OD���l�TpҺu8������/!�/�-Ѝ�ݫ�پ &ig1<����P ���.<����\��$a��5
����1t:V���E�	����b1aA;*���>�:��я�y�t�X��d�l�TBZ��a͢���[�R�؉JM������j���߻���Ka����7a��FFQ��d�����A,q�X���TB^á%p�07T����s�H�N!�I��'���}C.\�%)�42�z<nh���a,Y�\@t*[+�}>N�Y$�	�=r��~��/�o�
D�ii��+t85��%���X�h5�{VCsxQ5U������B�O�Ӊ{gg0W��P��b�o�P����Et2�W7����~�5I(��apd?ڂ�LLO���?��e���������
�h�9��A1������0T���.攼g�^榦�ey�E���߁�_x
�"�v>���T�@{:�lX�'�x"��U� ;�98vP��Ӊ$�y�y�u�.XN$�i��%�6�lW�b}�N�}�Y�����Z��#,r�S-P4�&&�tQ7zB\y�%ؼ}��"���Qs�T�C�^c�ZS�㌓O�� �l�z���J��,�jMX�|9���{�7�F��/�k&���
YTi����`r��7�;q�qG#�aA�b�w��18�ֿ�EӬ��ލQVr,~�M�r%Բ1�<�vQMe��g7cْN�1@0��<*V�lvu�f�1������#N9�,���0��<jբ,H�.�MR���Z&lڲ���fw#���g��A�Xli��C "�w���.�t;�z����y^��f��Ԥ�0v86�;;�/_�rٌ�0]�N��n�MO-fSҴwbb��Al8b-V�X&�_�=e�5*���p���M;�e�.O̡�w�DI��=�d�(��>�'�Ã����HQ�o�����_��N'�<�(Ip9��0|p�X}}=���A�T�N�4<&:��e�N�����(9�5;;�bA4g�@�P(4�n���h�Nb;�5�<Jj���f�J�mXkcvv�Ȫ���0�<�:�ĉh�U�Sn��t��tVk��!
�gff�.���i6!Ɣ��F�Tj&H�)a�ۛ}���Z�f��4�FV<(�oԉ���J�^*kF��f0LV��ȿQ��h4j�L���ɳ\*4M���J$e�Xo6
�mL\�iH�Uq���'���M�T�Y�՛&�������_�y][�N�t0�h��=�3&������fO��ՅL:�1�fmW�2�,��-�`��l>�<E��&J��2le�� Kk�IꔼF#�Z�20R��������fP��HM���_b�:o-q�26��%���t���S&��a�Xh���M�M��{�Aɘ	
gK����JWt�/���:Ʋu&/7(�[T��\vi���]���OCk6����o��0��;�'�JQG�_�흝xk�>|��[1��!�S�p;P�����GXk%LA)����Ux풁h�����z	�Ͼ�2~�ǇX��3r�\f��Y��{�cn�~����X�l1,V':������� I�i�����ٝw��o#�x9vOL�rLͬ�TH�����G0z`��������KVN��S�{�J�=�<��_ۄ�L���qxl������cd�<�g�m�.LOӣ��H�8ܳ2N��#�Z����1��C�뉿��׃�\A�\��B�5k������ϼ�B�x}�pj>��L��Zn���R�=�4{�u��bxbZH�~��n�ǬX�#�.��/��+����=m�܏��6Q�y~t,���݆��wcņ���B>�9p��sO>�r��,�6mK�	��d3"����mX3=�v������;a����Ć�T� =2�sN9�8�x�/�Oo7��/�Y��fa�cø���w~q�����Ȍn��u�NY~j�2����0�*.]�|�*����m�F�X�_y9^��6��1X�^�~"��?ԁ�lao �}.��"�lQI�V)�=��~ϥ3�5߽Nb}���1x}n�#Qs94et��0z`H�k�׸�!$�X�.X�i��.���v�ڎx���3�H��d*��@���\vdg���م�/��RE wGOL�*�8<F@SL�9<��[���Î
��	8vp̠k�M2��Bp)tzC(2a�����g�yF����ǣ��G��L�/v�=��&2(���S�Ș3s?���X�v@��[{��&j�T��#�I�P,W�����ׇT|V��0.M+4w��X�н_��Ͻ"a�Ӄt:���i�Hլ��=��39�4�=�_�,Ւ����02:(����6�]�����`vfZ�� �yFD�#��t�'��ދ��b���bDA��0�P,��`�����۰gp���`��U�����w�IȷD-���z�"L�"��q�mGZ���h�H�v8E0�r�!�}��طo�p]�~O����&�b�%�Nr}�2?�x�81ܼ����ف�^݄��aa�$����ţD��k^	����Ӭ��^Oz����b4�	�#&���'Ȑ�155���zaA8��&�Ê3�#�-�[�������sF`��iu}X픶s]��lYE��X|mk?���Z�F�oa��]Oy?�l�r�\��utt5�^o�\��A-����b~��#���s��a��������Ѣ���x�.��km:W��*030"��7?	X�x�퍘��)d�Ԭ�N�%ch�J0���^��Y�#� �dZ�rTh@�E.��29�g�yo�݈A�S�}��?�w���j$��H�9a����e���7Eyɪ�j6��Y��>o2�E�ȿ�(K0�4�,4*=ߒ���/8��4]I�m�d��\i������_��ͮᬓއ�_��!K�GhC���r��9L0;-2@��}n��vh� b�,l��+�N���_��Obr,.�=2�@2�C�j��@ς~=�X����om�W��m�V.�h|Z�1~�����xǝ(M�`h�nx�>��XM~��mpK�
M�ʱ.j�{~�;���m�:��s|UC>���~s�wQ��C"R��D� ɯ4���/-&��n������{�m�����0�0S��"��o]�b*��;�A9o�֭{18C���i�݃�� ֬�������ˣx��7alk�D&+m�Z"	���;��W���3(�+b�	��������B�X��m�ӡ �n�<��N��އ�dsS�hw۱�Ç��y���p��V �3 ��������
��:��%�;��0В�b�կMQ������K���A%��K����	v�� SH
 �����d�G���{�@�c���+.�ꂷ��럿
/=��ܼ;�"�n�a74�3��XV\����O�57\��͂�Ɉh$+~j�^+�}��/�׷��>�=��tw�C<a.\����O?߽�\��/�`���M#����&V.\�뮹!_�L�SڵL`ӂ����q�8TU<��Sxg�nX6��S�`@��1U�Ҿ~|��	{�����uR{w&�t�]�(���Z����/}Z(��rM���Cc�h�����.��چmon�ş��$C��0��\�M�p�X�Lf���ް9�;�b2��&-u
�*�^7Fw��綺a��Oe��X�d�6�{W�\��~�'��
��04�04i0�@���Ҭ�Y.����۾�#7,��T�	��d��!��*+f�Ia�����=�9�\x]NTK9�LO�uI��y�*�o�F�5�1�x�����$Y0�mu1K6�&���B����!�"����Aݺx��H��������d� N=�D�s���@�W[�� �����q1����އu��`��ŰS,d���6���n�ҕk��o`r.��^z����2�U�Mrcs�,J��H'gQ̥��OMc�E�(�NXq����%8��0>>*�d��~�o���GPF(�o%����H#1'�"�ڵo���|�����ݻ���) �6D|�OL�(݇M��b1d���~�wdL'���t;'���^Q�r�h@�y�s�� �ń.x�:����y�F�%ݛBA���U���Z��sz�$������^;��-�@Ҥ����YsW�>3L]��Vk�bն�x�I���,�m0��=x�g �w[G����G~ݴ��O�2��F<����ð�ˈ槰gri�y��p�ٌ�5�T�������t����.�V��1b!����h]8�^��E(��I����U���	�*�aR�ʠ���#���O{���� �m�V�?���l&鞬�@Uƪ"�:��ס�a6J��=�F9�ۆ��x}l�Dd5��A����RP1����=����X �3�fF"U�jQ�6.EE5W@��D.OՔM�Fl�ɪ�d�L��C�x���^�3����N4�b�����179���4�*�P6��n�>�K�ϼ�
������hT@]�m��_���9�
r�Rɢ(1��Y?�ǎޞ�ܜ�t
/oފ�،�j� �\2�JvK	���]=.�Y�+&LL�1:�ƾ}����>��6;�.#���p�-�1��ލ}SS��Q���_1�_܎r*�h2!-����L���ݭ"���Z��_���ضoe��3����'g��=w���`vb�T�����)m^�Ƙ��݅�ـ��	����ʛ[PWU$�9}N;z~��/Ǟ77�ި���C���*�h1�\%/� ��C�<�{��(Fqt/_���R�[��f����|��w7��z�Ξ���+q;����*��;��|_�Q<�⳸��ua�����9���]��<�|<pǽh4M�=x s�T�"�(ڼ~�"q������]���)<����{j
���b,\�
0�ŇN?���7�u���de�Aa�ö7���������(���R�-U+�eG�V�N?�\����76art���1�<~x!�(>���	��/^���6|��_���¾X��]*����O�����P�\���P¡3,v\63����d:��doL�c�R�D��9z�զ![)"�s���A-���m��J�l��k֬����ݍ���;l޲Ꭵ�7���N���^i�Z̡��yEA_O�z��jE?,f��e��K�R��P�R���}�(���~����BD��W@�La@;�h��1�e��u�Nlڼ�]0**���c8'��WOf��L�-��&��*q.�o;fH���d�b\t�G�j�2�R�Ѣ�4���
A��Y1��{p�1Ga��X5�Z�
�&�n�,���oB*[ų/n�T
f�����9lva��i
Y�RL�\.Hh������JHVwI#��sq�m ��~,D!���p��b+�yFDe�@�������Slp��P���'���b��(�"�R���Ֆ{��m�&`j�5)���id1���糲Պ����.�V����@|A?������yO8X�/�$���E�C>����V���XE���hJ~&�F��G����Ԉ�^�l#�fv��jR՝�w�W�����mޛ�{�6������j�<�����,���m��c�?5���)���j�t*/��z�~��V
�'X��wK���[���Oš��yPt8\��-�恗�j���9h:�(ת�&�B4�y��
��V.��F]T�U.e��;ɜ;���ml�1ԍ��I��1�A��WD�W�Nn�RQ�XI��n���le%�4��TQ�.���YDShU���~��;To�<�ͬH��r�,��Tff��y:B��-�5�Hr��fU3�C#�4b�Y�6�.�%�xFQJ.��Jе    IDATZ������dr�a+%엪4�j@zbn[*�U��2��&O���"jMp��ךh����ؔ8�+���:��h�
(�rPV�{�T/�EF�7���
T��tb
�U�Ն=�2�u�<��amo�1P�]J���R�!�#��@��B��"�kl�R�ˏ�XRV�����֭��&��h,��AE�ebZ+!򣣫S�_ټ	�����y0�����p�/܆?�df�ao�P*T��1�PU�/��ݮ�e���I��G�gbM��LJ�!�p��]��-ߺ���S؝LN�adt�R={q�1GC�Ꜯ�|�{�a����
��:̌�QKX�݉k��3C�0�V�Q�MN�
�+܎s?�A���pZ,����_�OLe�((N$s%8�6!g�t��������m���N�.�e�;�$#� m����3_�w��n�o���(�Ę�{߸���a���H%38p`O>�j��N�ڧ>y	�����q����bV1M ��6>����K�~Q?^~�1,^� ��3���A!]���gޢ�d�îapt�fg��ix���$f;�f &@ٿ�2�4�m6!h��ؕk�s����>��6��`����`㫻�G�B04 �=���Y�ý�inLMLˢ�@��raْ|���`ْnh���i*�]����М�H�2��{�����>�f�"�	��S�4�ۊ��rt�O�J���߉���F�X����[�-%��x��c��9Kd�(�LV��4;�SY�K,Z4���
��fT�eIB��F�ƱYr[[�l���W_}g�q�K�UBF��9<Z<X�z=�{i�fSغc?̚�SQ��*Uia�i��f�.a��y�-�ɺ�O+���rH%� �ݑ6�F�f[v� lŲ凪F<>$R5���|u��$V�v���6�n�*`��� ��cJA+g�W[���#��Z~�Oڅ�<&`"�XEaL�Ŀe�`�!�V���[�|=?�e�K����VRLyy��l�� �;����-m0Hu��Q��>��lM��#��~�3�^V�@e����9�Y�{�q��z0~���J�=������x讦�s}��^sF����lqg���ѽ��
���B>�B6�hA1���	i5��T^-'D٢Pc��[?������ٍ����­>����d�VU��@=p��(ݒB�^z&�>�-���:�#�b�ɬ8��, ��S�����tT��萹�\�ͻ�Pd�w06��88YŦ"���N�Ь� _Y�N���J����LA���H���HR��݈ժ��4��5'ʕ<f�s�8��6�~d��X4�*�u��Hw8�B�-J�0�j�#�l����:�9��+�9xl6�2qx��Є�bU8t௕3"u�wU�^C&��1	�ND���� ��*
���E���/+F?1��JV��&�E_[���p�f�i���BV���YȠ\���a�8�-"[����OT�ss�@�C�����8]�d�kV<�N7|f�=d�b������`&`�s��D���f1bvjn�
B}��.�0���f^�j��\|>�*L���Vm(P�=6�]�v�Y3#�/�Rg�x�ͺL�BʵZd�eLu-��ɞʴ@�G�R�|Z�{_ �d,	O[�B��>TU��+c֬K�46;:�N�
$2���]�R��c���y�|�"d�N���� �/ �ʢ��`���#C8i��(er�����2�/	��2���������d�}�����8[��QC��F�*���;	�xo��Y D�j�_7U�~�1�;���lzi�4�Þ�k�U�f�2|��VҚ�4V*�D0ԎSO>Y��G�bbj?��p���&`�h�@�L������*�ڼ۷nE�G��P� O�U5�\��$76=�s�(x��6:��fC�Zժ���B@Sa�'�n`��<��h��
��B8�>���;h[�ZÎ\�Q�Q���,B�-���IXM&�Z� W]�1�[�����T�:&!��5���bG:��7��-���G�ū���>%����y6�I�(˰9�������ƛ~(�/��+�C:��牀��YN�<_[��,Ǉ/��gt|&�����E��W��7��/�� �gj���Z(���w�q��atvzq���b�>��p{\B�z�:�JŀO� ^ym6m}�����oG$�G$��jۑa~�M�1��4ʥ�XyHA����v���r8��81;;%^�|p���+�j��C��_�I#�C�gEj.[p�{���H���XB��R�CI�'�=��)�I��L&5|A՘3�-�9�1#CÇ���-�X�-	 YijEM�M0���'_�"�����(��Tӳ�������(�;[���;~���"(㢄`SVL)��u�/�#��u�
�;�09��iRL�ׯ?���C潩��-���	�n��w�������*�����:�p:��
hԒ(g�ⷣ6�[>W�����4��ר��V#%��?I�?��*]����'��?߻n)��А�z*9GT���f�F��mW|����gT5�PhԑCCZ�TB.N?9��u�O�-��Br�PI�g�
+e�MȅɕC*��k�TK�*f�5��ج�bQ8�f	��:�����x����Fdj�ha��y� �V ��4�����)~ a�p`pbma�<�PA�[�ٌVɄc[�QI>�G&Lz����$󏼞"e�F�ҖD#_r�h�jU!�3���p���XD���������Ѵ��'��ٞ��a��rx�\A��(�p�5�.������xdp������(M�����/8���֔����@��[
�y��tJȽ�JY=��U���.'l���t �se�EH��	�������� ��ܺZ�j]��R�E��/�о}B�R�����p�F����v��	K3���}��M�Uq��`���'�6K�`�"�rV2����1)Go&&K "�`u�F��b	
��D�8.�M%�E�:3��cg*�	�fi�y�Uԋx�&��������
vee�Qhq`D���Ea�	�79��+(W�	e*�v�6�UxdҢPu��SC��h]���L1;yc0 �ʄ��C�)�$+�O�J�>�`���C��[���Ǌ C�"rc|fMՀR��t��l�$����Oxc�J�r��8x`/�߇������@"���{�t`�K��~�� iV��ƗakcT����މE�~�,��C)ců�|��a�\X�f5��y [�@[h�����nڬ`�i�8=05UQ�QC(��w��E�p�:�ky�v�#	��S�d��j��i�*"�\Í��,H&b����cnv&�|�d�����[a�8�\�����O���>��"�c\��D�!و��Klё��q�-���K��_���Zؾ����u�@Ӧ�!��/Ɔ#����|�R���xٚc�E�Oy=g�Uy��xi�رk[���\4Us	���c|�+y���t�09:�Z5��"U{����?���b�
�^�[��Dt�����P� (
	��?v	fgY)$Q��I�EI��qBO|�[�����{9��ļ��Q��J����A~f����8ɘc4��Z1S���a���'?��	kq�Z-�Ýd>=,��uZƽl���ժ��:Z��_�&S	���}�}lUЄ�'���Y]��t��v�}ς�K�b�Z��_	���4����[�z�w��a�[�����(�h��PN��i �7,F�^��g��j=*J�h��[t�:����ɉ<��OY�[̇�][���ۘD�<��R�K�4]mɥ���`��/!���̠H�]�U1�e����1���ި�ź���]���d\��b��qN0�	�$%�@ �X\J�JU"S�*�OGs�	�I�+ex�NL����*�*T��s�X�a����K1���0kȣ�B� A��ME� ("�����,���"�bA&���a�y=����� +�C5 �H�Y.�i���/JLN�h�d9d?�
B媌�:���f�c!�9rN���������g�J4J;�i��$�JE@��5�r4��"RmUo0s�%�g%�FU�Q'wt�K����V��`�v�L;��\EӤ�P�i.�̬�1��>KM�:���<IX@?�&:���(2~�50E�N��D��F���l� ֽ�j��^}2�B�yr�^��.�(V��S�Ҁ'��j����B�lF����U�U5M*jeV58ț�b��$f��=^9�'�`�9���,��X���{�(;��JtW�U�n��s�э@$� �$R")�
$�d[z�9'�����~3��z3�Ҳ�h�T6M��42m���T�HR#@��@#4:w��s��}���mj��֚g�P�E�}Cݪ�η�9�썼O].����ZmD8��*k�_G��E�"Qէ
�+F�CF�)�q[6��j]
�L�x��FD<Ez�IC@b�����w l�_Z�C�I�Fӊ��x�m�kI~[���ґ#��/�d�ޟ�	�ဉ�@�̪b	ղ�|V�m�)8fW�ۅ�ʢ��O Z�K��|��s�琌��x���NO��qL,��ɦ�C��<��E��p��ݸd�i;��Ϟ���
2�>��ana�x�;HgG�89�w���>*��l�L���,�uE�O�,�w������hV^��b1R7�K�.�IH+�>�q:t��6��?��p��	�q��Ɍ�v,�F�E��n�w��8��կ���z'JS�·��tb����'����]�`��1�אI�M��\�[o�E��x화p�ׁ�IO����ǕW^��C�8"��1���%3�M\��J<��O09�ǃ��!񞥴���| ��"��bx�3��V�y�$f2�L��x<�s=J�B��@VI�̴���D��TO�~�; �9t�Z��#�#��6�Mo�EZw|A�{4��5%ӕG��(b����^�۝�ץۺa�5?s=[?_��������S��䗂?y���\\�����'�sDPK\��t�����!����=���ݶ��P�W�������>tǽ_��F��k�~Z��.V��� ��]d��0�G�e����M��N�XVܔ,h�ؚ-A��;JB4�X��#��T�?O�U`?^�:#�!�Y4U��:]T�g�^&3����  �:�ʶ�&N�����4�mX=Y��/I&K����nS	���?��p:�)6�-7�v$}$*�.��>���₌�W)�hX*q��r�XLDX�Y��9!�jh��1��yů�f�Qw\�,�?:��Aq
p|����i�du(n�8r�J�K�Kf�!�n�,��Rï�0��Ь�|"5P�s��Mc~i^Z�I�C��@��G޹�[0�m���O�ԫ�>�
�`�<:}�2P�հR*"�d��E�r7*\���&13?'�45�FCM�pf�t��Y�'%&��obi%�����dˈv4��#�*�C�X�1p�@N�ҽ@�˱vE奀Qh�&]7�k�U
Q����$��Qo�I@����<�\`���D�s(ϖ.̈)�
h()r^D �ڮ��j�ZWU6�'�Y�c�@f1��U��E����j��s"Ry�Ģ0\K�t�xZ�"3��*41�8����-��,W�arB@�D)�͟W��rE�	��B�Rpˉ[�DV���@Nm�|?A-uM�Z�k���t亱rN�>��몷c�����&�}����ٙF���{3pQ������	�Ù��pZ�
R	�K�b�M���T���
��TԹa�>4]ӕ"�t^6+V:�Fej��G��݈�ҌLY>t���j�%�8}Cè�|�z7�R~��SXZ.H��r,Ij���6l��&$n������Fo6����(ҷZ�7p�ЋY"�Z�лՓU�'�'Ҧ�x����'�t�9��rj��+�2	᭼�\F�����5|������y�YiO���?އ�q�� �Ds�X�`2D
��ܴ(���[���9��*;z`J*2����ż ��ø�˰RXƞ�w	 $��/EQ	�H�#�5����S��ґ�xv�a,�KH�{�_.��V�/�Y����N��Plh�'6w�"�֢�E����)B�
��?�x0�;�oX�WU#z��$	��9���m��E�[�l�iR�"JW�cPU������y�I���Y��.�Q�1�ʗF�
�������+e��V�`���3���y͸���|�Z�D�)���^���d���%($�@�A�\9/�f� ��a�_����'��_��;���Xz�b���H�P,̡'kb|�Bܚ�U;cx��!��C�XFy�&���B8oJ��/�.e���c�ր��hzi��/����	��F���u��b��f툉�ǖ�2�%�j!��j�y�Y<v�|��MC�ؒ�3ӧ���S*�1�-�Z���B{Ʒ��k�Ŏ�[�Ph�DcӉ ;؃CgN�C/���CܸA��TZx�^�������gظaT6���?	)��o=�-�q4Ѳ=t�.�4F7���?�z��r��do��"�H}�L<���3���>_ī/�S��k�)��z�0�����Ml�|�k5�;uT�6�Te���iF`�L�_�/�(�ԛ�\����dЪ+�@�bL�#�(n��xF�7�����c[��ɠ ji �\!�%*��s��\s<���6�?G%�-����{Q셣�q�� �t:�J����i�!��Y��\j���rXy_��	mi;�V5����H�t�MX�I���K���f]@���X.�l�� �u�ֽ���Y��z�?< �|�:�������@�NM��	7�Lׂ����i��J3���:�� \�'n]��ևGN+�l���'�%>\߆��/�@i� U&��=�vh�E.��+z$"�~n���$׏߻T�J5��l�1�9�)Y~ �ɿS�X���Wc���0Z��5�B�J,�V���`�r#�W+�V�b쾰��64"^^���8��f��LD��M0�N$Q-�Ѣ�!5#������A,��ߨ�+��]\>2�kv]���i\��l݁��!�׏�>�(.�d6m�.�Hr�>����Vz�8j�&f�q������mv�zߗ�JD�ϓ7���Bi�]�HTt��j�������A��NNH�`%� ��rr(g�*�+C3^���:1��'@��&�lقk��V�9��,�������t�r�jk�jr^���J���oŖ�MR-a�����+��,�V�8�^S��O~�3��w��.�&�p��;��#f�QkvQ��x�g�q��94Z�=�����/� ��QT
�رe�zI�#+N���`��Q��#A�M4��wA���J���'-ٖ���ѫ��#B��" �b9�����'{TTU����ꀄe ��ii]����z`v`|�
��i�����W.�k��0��1�=��y����31�{<����$�g^��P�Uڥ��p���i��aF��B�G������#�쎯|�N�^V��p�Ģ�Y��������wrVt��X$��5�p����jԪ/�^��S���lDx����~\�\�*��6�GBQX%C��^�}3�m��'U�QX2�,x��?5����	�g�0GAZ*�Seɨ�j�p��1Q���	�,����2�����)~sS���O~�TOc�8v�4�9��gOcx|�S�hj��W�}�z��}Z���ʙ�s����zS�� �ʎÌy����q��Qky�1�(Vh�n"�b����־aL�������ב_Z�K�ݰ�Eo��^���8I��P����>�es�5L4uN�v�����Ͷ�G�yaN��y~ԍ'�&�%���*2�h�REla�6|�6�����Z�M3��˸����gP��e% 2�1V#ӵ�l"�ސv�C��4j�p���H+1��cn9�Vց8���BkU��L}t�����6I�\��D�䜰r��$U �	�`]+��>ߗ�b����,+    IDAT[AI�W�], ��R�2j�����El�C1���sP%��)19��z�Z�!t��k��Rԑ ���Z+i��<6�RGu*%)�@�Q:Af�-|��y�{d��-�@��l Ae/`|��/����a"������ے�g�XJ���z��E��K'�P\A�\
Z�Tr	���pW����Z�R��6����J>7\ݶ���ڳ�a&$�6'&0�p�E;��G1:�����+�v^|1��6�?���MX�06�I���T�������?��H'�1;5���>����p��l�g��O�ѱ!�;U��Y6
yU����WKےհx"���,�+��Q�nD�g���1��h��RיN?}�g����S�Oc���ry��J0��(�r��5��w��W���kC�"^��t{��ӛ�<擒������9/<$Ur�{<�{{���?$C�<w@Z�����rF?-����T SC�ݨk ��Kq��!4���l!��+����^l���	�=��٪lR ��� ���
�`1f��ʎ�,�-7�ғ�R	
*S��&�.���nG�����iФ����{�a��~�z F��A���i�&�RN�v�~̪�~��UV;AeQ�j���Ϛ�}�a���(H}�+֎$����Ȏ�4LDZ-��@�:���6Ɔ;p�3�����`����S�kb�J�8G^� ,\���0�E�.�/�j�+$�*z_�h+˿��H�^��J���mײe�IqJ+0��um��c�k�K�'~�g�O�O�D�� L�A�â��ioD ��]l�-���[ކ�R�jS��sg�"�����iL�q��ǹ�E�s)�&{p��p��d�It�m4;���'��~U���".[�I��6l߈�p˵%�/j���S��5\�����Gp��f8�&�x���d��vb�MO!�/�I��sR�x��1�����M��Q%p���>��2�Npnjͅ�Ԅ�Ҁ_oK�GԦ	��ob�l9��-SAݶ���	R�n�\c��+��ӏ�������w�M��M�) �6�^;�\W�ۜVm��#A�b�Z ��B~��>���*"�_ge�a)6���IJ`80���<��Q�+
�T�*�*ۢO %�d���l=q8E�虵��C���3$�
��0K.��0_�6ڰ�轕�F۵С�AD7u�"��&X9㄃A�$^�`5;���*���mN�s����[��3"mN��XU��gU�g�B L��!��k��������E�̫|�d� �5�*�T �d&8W��Ȼ��7�+��	�`#�ː�D�[�k+�4�.O[���#����-�9�����B����jŐ]؈8��a�L�Qn�m�\#1��Yx�x?b�,6��q}tOhw��T�U`�P,����E��V�J同�b��<��ܽ@7�N����[�ۿ��q�e���=�Pŋ/��?|L@ضc(�PX�����|�>��o����P��G:��0;b���l{lp�"�ĨҒX�E2�Ȫ<[�������7�R,�95c�Cy���z�}�v\q�صk�PT[������҃�`�'g�kK�L�TF��?�/�?z�)g1�i��vVXb�4��.b�2��:;�7��0-���13��ޞ!I�L���\W�ݍ�gN�c*m/N-J��SrZ�B�*�3�}��(�'���"�+>�B]����G�כ^w�|F:�Z%��LM�'S�Eо�n=Jbh�I|
8��A����w��F��qkB�/��Z{l=�{j�ǿk��S�z�N��z��`(�U��5�� �L�k�m��g�P㙯��+¾���+>r��>��l��J�l�'�A�>��t	�7u1�i�������t������w�(Ljm�X^[$q�?�ףp}�UFppX�W�iE|��RD3a�٪��:h٤Zu��@�A��`EP�d�?���8�f*���P�3�.����c)iBSH�
��H4L\2�;����;hkHEc�W꨷��t��w���JfV2&�P2�;��ؘ�o�ӧ&�s�b8~���ǱP)��b2�H2�'��#H�fPh-��K4Θ�u�&̎���N>��F� Y��w|��JG7�j�\@������/,`���%��tL�����0h��u�k!��^�����kđ�\�ȡ�;U(�V�t7:�t]jVs��4���QQ8��d�b�5��-��+��䉙t\+L�C`�ydƮ����?}:e�HPb��15 ���g<fV(^+�F[�IO�������H��{���	�KJsuU��!�&�#��G�������è5$�H)�2()	��!y:Ғ`;Vއ���2r%	0��q&?�2AX� ��{�Rzs�|��ڎ϶�k�mg˹Ձ��@W@[tі	�҆Ul�k[0���B*��1����9R�40�5�c{Tt�h`��S��>���ҲU�M��.�W5L"\PVjİBm~jc�yQ�Q����D���u��$d��^oz�dc	B�%�W�S�4���h���Lǵ��[^�$̱ܩ�f�f�1���,5W��1�M`��`{"�]c���'1�q+�GFQ�T102,�m���x,'�K�)�d�)�͉���E|�λQ��H'������=;1:6��><����JNd_6�
����q�W���߄驳HR�,�b~aJ*}���\��i��X�k�|T��S99O��Ze+�ׇ���ɓb��*��\�$es2�v:�pC^%���*�X���t,V'�X ?��Tet8u�<���/cjjF�^:���v��I������˯�W^���q����(k�\R<J� 9�a�/#ڄ�	��'G	�C�Dx�;U4 i?�W�=�: ��<h	��4c&�#�G�m����Fyo�3^�U�� +պ�0�U��	�&��1 3��0���3~��Tk '�ڗA�-��@l=�
�N�6F��	�Z�sm�Wq[���/�FQZ#�w�Yی�c���a�����+���wR�.�5,8aq�U9�L<���"�9Żo���s�1�H�Z���ͬ�^��2��r���E��S�Ot	2��+�G�������"��O7خF{�JwF/V�H���ږR�oY��u��M����(�{�	��0�j,�*���A��w8��(��Of�vd��h�;�FP��ǀ�?;�����^Aͨ#9܃�y	f6��i�����M`$�B"��S'N��R���iU1p�^X@�ZG�M��e���0�k��)�k0�&��6��q+���Y�~�E�ݸ���/��\v9���z��
�:NNN���s��d�Lǐo�`x6��P(�c@�⃱(�Ti�,/א�F�i��vY��['�M\G�d)�J��^NE��#�\�l�VC�.l�C�݁A^J�%Y�O� ���E��rn�܈�)&]Bg�����a剭�B3p����V��mEԆ�b���(�'^�%k���j)���ilK�F�:(��ARG�i��&��vb(qb(���>���*�����Qi����ϊ��B��(���~xT�-`%���Ҭ��tqzv
�nC,�Fb�C���Ꞷ)]N�%<�>lue�Zl��@�T����X�&b�*5ݺ2��|+VH��X��ԛr�b�T^�'�&����J�$��*�iV�r�Q�UQ��d��*�:�K�3���*e`l͂��Է����̜����H�T�p�Z�GH?$@sh��B�r�l�$�zk�ZpMQ���̘����Ly񴅸�F��1b;x�uo���+ߎD*'�+�Hr�	Q�cY!�g3=��>/f��6���J�c����_B��E�7������st13?ǋ�Ҩ��:�LcqaJl��9����M������#�ɒ�MP�	J7W$.�)*�ј��X4!�Z�f��ϰ�zt+����X)k�@���hN>[���(�򹬈r��1�nK�I@V��Z�a>�P�$�#���u�ؾ�E�R���Ż����	\{�x�����{�C���zS��E�[$&ٞc`�@M��b��SH}.�8���w)�����*ykkDvE�WR6����yn�/(S�J���b6��@U��[o{s�<�P誖Aʸ[�'y�9U�s������ LW�t�"��N��V�Zh��w���;W��5��g�=������$��Z�a*��I�
1L_Ρk�c�Ν�a�{���+��}�������G.ow�8Z�)�\:���6�m�`SO���oFm��r"�ӆ�FQgFJ�ۘ�F�.�$Y��Y2ce�&!4�]
�BK@6�i��}�ѼZ`��yI��1�4G��Ѣ1`�J3g���N
�ꏟ��zը�z�a4��X��P�E��ْb�հ=#��],bk����۱85�N�)���(�s�~ّ>w��>�/q\���jSn I�EO.+��r	�~�;8s�,�XB��K$�'�������َ�hE��r��B�*���r&:KUL<s;�FQ>3��o{~��_Gai�l�s3`���?���p�=������8={]�TP +�ɀA.׃\,�Ak���\Y��ϑL�u%�K�%����n;]%���Qo!�ʉ�%T�J�U@�9�P�+S}lq��-����r�6����0��Njs8��.������=I�>; �jT`��Z���[Q$'hip�\�
((�揪����C8P<���eyd���j��*�$�ӕ�j��f�Μ��c21�xD��m�&osnⴜ�2!��5[B�O���H��]�Q��X�!Z�$d`�L��$�Z9GM.���>?;'4�7��� �3��I�LJ�R����kIYI�دV��L��:�El�]]?��i�</Ș4��H�v>����
���*���ͪ7��I )�͖��
tt\�V�е���FS��lC�IJ%�o`�JC@:�^�b��cR��/sʐ�5�D1�X���~:tG�@o?r�^93��pbQ,��Qi��a|HD��eN&�D���{;��k���Ԅxq�"����P�K�S@ 'ߊ�J�������¢�&rC�@"%���+��QO
H!F1�چ�ROW@�*<yi�H���uq�r��ۆ�1=qw���9=���Qi/�-,���;��KW}���8u�vIYpU\����L�Z0:u����8��S"n��\�!@I��$�25�����Vabkޗ���:���&�9Z�tp`XX�ۼev��&@,�!�R1��x)�F��Ɂ!NY�'��F��	���0�-�o�<�Z|A�C�NW�t��{0��Е2�N�N�����C�Ĉ�	��R+�!z�|�����5��5�g̛��v�/f%���^�_��ϵ���kM1�� 6o �2-��_~�K���\tV��B�O�C��Oښl�)���w�ۑ>��u�M��`��*��	o*)iR{����R-)_��7	�Rʥ��`���<�T�I��d�3L4�f�5<v�E���Q��y����l!��Y�V�FjSd��@l��Fs6���pn}�kq��q�y�!�Y����0_^F���=#��e���p2����(.-�%K��s���ѓx���Pl�P�(�M�qWT����"9��r�#�a���ɭV�!����K8��1l�c�I�ݷ��x��p��I��n�J��|����&���G`%��q��-���H�X���'C�M�]i!�v�\��-���D����3;�s�j5v���D�E���f.���4���d!BM��R�ΠF�ZQW�ށjA	�����-r�9d���֎�Q�*�+�v�Q��&KH�4[_�WO�[���$"X/�8����������-MYڱM�dT#'�2��n��"ZU��i�E��luYyyn� U��m���l��C�M�U��o�UT�#�&�RG�	D��|�H�M�i�Ͽ�n��Rb$E�D��rMΥߡn5�q�4gO6� �{�ɚ�®�0}�x��qe���������Y
,ȵ�8 � k��ڰ��M�9~f��p`���Ӆ�vql���PO�������M�Plv�؈�ͻ�ƒ24�%H��E�d/���P�V00؃V�����U�&�zǏ��J�(mi/��Ra	n*3F�,�|�b��]h�J8z��.Л�p�MW��8+�]E�D~a^�n��Ғg�,�0f;��/x��*�����d��Z�-�0�B����*���*�H��׃�``��S������覍�|	_����Y��v�B��B�2>���"'w�Ң���+$�M$�)(L��ģ���?����s���O~(@� �֠�RY�h<7�c��`
��s����Aα��A>��cǎatt��7��^��kQ,����Z��ga�2�$x��F1b��TEL�0!>\W��W�I�Z����5�0�X8~��KM��a}:.3��*����$�F��6��-���U¾����|�������kvl$��|�P-��� 0>�ŶA��~���;�^'��(mӔ�{�Y|�{��N�� �ܶ��eA���ߋ����� 3��2o� ,A<����m��/�^�Z���B�g����հ`!=���
�:r�f���Pg����HUo�<��AuD�İ(ӅKF����c��p��=0[\�>ʭ�o����#����=�/��i�.���Zq4�E���7#??'��?8��^�#�~K�"��@Y툻H�eK'0�mn���jf�C�ے� ��Jb��<��P,��o����|�0[*Q�^��񩻾�G���1ԭ.2�YDc��H�],7KB��X���uKڑ��*��#�d��.e;���x|+��"%`I�^����^V��3�_�0GȺB �ꈪn�:R���>	�z\Zs��`a-�
@ͺ�\�W�
��0j�I�MG�d)h�AҚ��,gy�����X8����j�I�j��
��(��LL͜�<�`�D�I���qӴ]J��qt��ك��	��%<��sj�^L6͖i�深���%pzMչ%Dچ�hк:T�h���V��7��X`���Uૅ@�*��+��NU+��0wD��5�vT�W�@o�:>�E�VUS�)�s��@oJ�N}O�j�D�6XpHn	�:�|^�$w��S��K�H
���m���9���G"݇��;����T��LE���Z3s+ro��m���i�A"5������Ph���3��6]d29ikF.�Q�F�C=��˰8;�C/���C�����^��A������݋�������T�X�f;�\1���Fm�F���#��B���k'D�%��D"(����(R%� '�4�)�T�:AK���r����������ܬ豝;?�r��E}��q$�ēYL���*+�MQ��Q0[o�@� ���b5��;����⮅���G���8/@�q$�/~�LX�桍�uB����`J�K��;�5�,����'b��Rl�2�M�8uꄴg��!	���]�L�*�E��*1T����/Zuz�(�a��wpi��r0u��I����[s���(�x?�{�JD-�p�3�����<���P�`�2�{M���a�x �·~v������"ٽ��%zB��@�2���&F��x�����7�p���Q��0�(��"������
:4����A/4yA��KK��-�+�W<3P�a2�)0��(t/2A=M+�kI fu%�RSjl:O��(�K�\~��(������c�
��d�M]�)�U]��T��ڛ�m�Fٰ�y��@2�C����ch�R���#(/�׾��E���_A!�kNF�o���������P.�������=$�2H�f�q�FI3�yd��i�V�<s'���װ��&�0�1O��W�W�܉�Ǥ�À�c��?>��>�|7��P?��m`�)�+"�l��I����'1�GΏ��PD�񂍊�Q�xT�.'���P��@􋣈�˴�7�N�+G��Ցpucvڪ䭕�}��%�TS������H��ɲ�V�A�bt�[[k7�
n'i�    IDAT�ɼ@���L�<c%,6�;�$��	�0�6X�4[mG�+&O�X�6eMV��� �c�j(��ݗ�֛nB*{�k��F���ߏ����r�V��ǥUtbr-����Z�YFܰ�W���p� ��Ť�A�@O�����(��,���<�6��kch�[ORj��>��L] o��@M�o4ј�-gG�2[��u�s��k+��*�l��NPh��F>c�R>��&����h;]�g�	ǯ!i�xӫ���@/^8t�A*5������⑚��E,�A�H>��H��N�O�0�V�����pLG��l��k���\�п���]�뮻3���]w`����b���3���r�_؏={v�-oy�x�*Ζ�V�*�	;T�'���V��U��_UH��G�ir�(����x]Xq�-<V�hU��|@̺99ȵ822"zd\\��5�n	�r��D2���`%��d~��x,-y]�`3E߲]�Ky}�a��05=�{��?��UG�B�"�N�f[j�Q���:��� )ҽN���\Ǔ���7�N|{z���+�*����FM�'V�U�K�0*�ў>ˁ @��^�z�K�,h��c��׃ǟ����F�W\/��h@�?_�3��iR�+͋��$� ��p��_���0-3r�iڟ���}��^�?<�׭�Х�bf���C2�26orЛXƎ��WnF��qdIF������L�#��^,TQ�=P�!�ޘ�X-]� �����-b�bm����]�¾ 32C�Pm���A-"NQQI�^���噪��`�%D�+��.'��+E"��ǉ���x�/rZ��N�0S���u���g�Tf�[��޻��&��4/�h���o>����
�΢Ш�޾�۱kd���cj�,"�+FT���g����<'�b|�1$�3�璢�x�0�c�'�_~;��N?%���#g�|bR�3������l���y�, �I��𩿹O>�� ���m݈�@
��'w��n�*B��zͺ��/��pj�nv�G e1��m~ s�l�I�$���L[�"�#����r͆�li���!��E�?�y���)5i*v+Xk�D�lNo����S5��4��ƫC��0����ᠣr�O?���t!�[e�h b��͎�9 �ӑ���u���4c"�J����-���1zY���I�q��q��ΞG�� |�[x������Mb�]��\��:��^;.�|U6#�xh�ōJ�D�Q�>gP����¬���`]k���[��ҩ2q>_on��u��#�A�^s��9cՁ��c#a��_��jAN�����ޘܑ�ɇ(�L���0�;�v��d~
��0�U��p��K�}|�wn���fg��,4�L� ��yzY�J���^$�e˽�$��ơqL�����GP(����I�n�tE��i�\/c�U����Ȁ���xm9�/bc�`~�.�;i�Q=��_4o����b��u��J�$�M�聾^9wuZ��G�#��xBp���y�����u�ʿn29�Պ����Q�����K��ĉرc��(�_�0L�SQ݃O�쎅L�_\N�>-#�3`lqݘ�5)OF��ߤC����߇�z&'��������̴j��ղ�N*��ou_��_8iZ��\��j���i�]c[5���k�~R.�s�v��w)��4�ł�މ���?d���h���9֜��P���=�Z}o��AR8���kF$g5�j�?��ߩʠ�h�X��=��t��9}>�݂�1�m�}�4��8k����<�����X;��>y�������mؾ�X�è��Y-t�s�:Eþ�~��7�x�0r,a�2EΏe��<���ĩ���J�bYZ$�4Z�ie�Y���J��-H~+A�Wʤ���m���Đ8�J�BЈ������F�}k�fbPbLB������b��2t�m�1<�8`�RJ�~[6
�P[i��8Z�~������0��%Y���#���v?}�1t�"���h鸵6~����W��VL����xf������{�ԧ�T-��V^�E$E���c'̈�JX�.ڳK�X�ϞG�O����M�b8��[o�Wlنv�����{��񩿹/>�n,��M#ذcќ�j��l����>��ګ�|������߃�M`Cfv͂_l"iFE��c��m�! ��Q�w���p+�2�!]	ܙ�ʍ�j�oDnҺ$..|)�Sm[��A9�ן�e"�|>.�A��U�&�+����Ѭ�CmE´B�5��
5Y* a���]GJ]��na�nu`�W՟�a��֑�;��r	G��v=83�4���n}����4�C8�.�Vq|�$��:~��qzn��^��	�(�Q:7�,\i�i�+�Z�'�}K6A����$"��?��������w������3��� �����z�)�hhJM��x<<>'7F]�����uxAE6�_�AO1b���gk�����&�B0{f���
�햛���*홳�[D�\����GǱ�ҫ08��Tۻ�TJHg�P�Jx���3_��P-7��j��eQI8Yi���1�u\�w/�x ��q��T�ї^¶�c(�,��+�[ȁJ�r�\��R�`Q&A��)��*'�k5i��1>�LBR~���h���Ǥ�M�_N["�kU$D(JlZ�:��"�ʪ�p��\.'�8t�b���Y^�l.����u�'�O~i�V���1��
STڐ�o�-	jܨ�:m�ȭ�pM<��71��� ���~3s��FȎ�{��*�����0����EJ5^�	y�^")�K)�w12<����}B�+��ĶG�5��q�E}�h-1݆���w(���� �J 5E'\�^�� 3�dtB+�5d ������
����.��\�<Jz�����0�D��S�� ,�i��j՗J�k�P��æ)wW�������G��V�z]ׅ���ǿt&}�gdB�7�i��Ҧ���I�Ȅ�gMRj���d_����|(M@im�7	..~��2���%�FL^�L�b�_OMV��䉨��m#���Y.�5Z�@T��J"���p&��U֬*�Vz
�"�J��y�Q����#h:���M���:�s��0?=% ��j1��SO=�O~�3X��ъ�J[,�!7ԇ�z	��킝t��-��Ql�P��L����I;r��)&����܆=���E�X(�Rm⁇�O�yV*���/���A�-Mcd(�7��
d�&6cf�����=X.���-����ʦDoQ���Q�$E:��D�f�kf;
Y�V�=I���a��Wi��q�4�Z)N���U�@N��NI��-�6�hEi	-5-�2��^UT���j�*�%�Bb>'p��W������"m�sBO�[��������0��}�EeՑ���ʤ�m�	��i`|`P�#n�CCC��� J����"2�,N�?���`�{�"�#!���Y��0mۢ+��<nݎ���\����Q�p�_?	�!	���ZѢY n�`WO���i�9����c�V��I<U%0$��w<.��3�pPD�V�������F ��-�WUp�0�0A���Ȕb�V@�T�;o����ɥ����C=���{��ah�(��E�/RѝB�Q5�I[,��ce���bn�W<;5��j(�a��7l��K/��cG������#���*�Jn&��ȥ�ur,�&N �I#�bg����v��&����k;u!���%«"�JAW�1���xG�s9�妨�3c��M���J����E��l�6�㙧�����5ת���ZYQ뵖X+y^BZk��ʲ���Q�@���徧���m�]�FQ��'�|C}I<��G�innF*t�ލ�`�\B���T�+Bdw^+�yݒ�)������0������I����?<��4i?��Z
C�3]_�:� L'���.z=��y��^��{8�]x���#��{�S�H�{O?{�zLKrmPJE}��w�X�Z]���0
�L��g�7��u���c�?7�����+V	�럟�<rGlhǞb�T�h2=��ƣ�YSxՎ~�-עp�z9V��(6:�(��L��w߇y���3�1;;+ecV���j3#%�����f�A�L��"�����	�͖�FɺԯO��q�J[-���u�
-W:��1����h�dq������3#���Y�o���<o߄��Jf7,��/�#}X^\B�T�L����ķ��=�4��ˢ$U��M[q�u�������~�)���g��'>�)!�[}i�,�Ev�3�9\rե�21�4��RQL�?7�Q�!���I%l0�vd�z��x��{�tnZ��33?����8p訴�����<��_��O�Po
�|Í�����fF�<�Hx��v��V�k ��,u�,F�K8ۅ�^GGU�x#���`�*�g��)�#���Q-z7�U�*b�dҶ�DZ.�5�D�*5k]�WՔ5�ka/3٨�[y���-�<D��AL�p5�4��uA4M�]�-��^��S�Q��r��5OZ�g&���:�w�er.�g�����HzQQ#g���I�*ed�{Q���&'ӓ�l���k�@��T
~�&��v��
��s�t��$�iv�XX	�ky]�-��y�ޙီ�l>����k����H��U[ym�Rg�|ݞ={�8�'%Sj
t���Z19N���nB������Tq�L(����cc�Z�=Lm��2�N��Щt����Y!�w�8�c''q����ܲcu�H�^Z,"��G;b�R��ǣk��W�l�X7��<��'��a���_ݤeP����쏯T�1���Ȟ��\�6�;LTԴX�/+,z�CA4�.�M[��t����㵔X΄K�QU�� ������E�B�ť<<7&\U�vEʈ2�+K0�tB]j׹	����-�N�jCZ�̻8I�Z�-����z�V�)��*2�����ї�#�3y.�P��!1� �b���p�R>סN�=��i�G�.����]�e�4��?�AD�B�&�K�A�Zl5��\����~�����z�N�nGj���Q8AZ�>�7�צ��DU���?���X�x>4mD�N��V�ց��� *���������1� �_���_��+����_���3�q�%+ņi5؎l�R���6��<�ؚ�o�vO�p"�I���x���#�%#����߸@�-n֦�Qp��Q}x VZ��X�j�Q�II\qJd�c�1�Ҳ��f��L� (��dܺ���fE���q��ͤѓL�]k	H#�#H���(�YZM��
�nَn����?��lV�tQjb~nN���|���wÈX�,�[B_<�[���}�����#B�\��E�v���~�����a$=L7j�h��k6y��6FwlB<�@�UA�]����[]��1����s�ۀ�������!�A�X�f�������qd��t�M�oȢw� �"��<^{ťx��W�U������gav�����U��j*�&�&
Zl�z�=UcSg�b��C���?.\��q���6\�L���2�0�' "�i���#��SMܖKU���=W2R�\�>���T�jm:�\��l�RZW�n�6�ݵ�W��A-\I���[�)��iaCM�@���z2\������]y�G��t�H�?7EQ�.�E���K��W�t.ٹC86y_�Z"���S?��}zqV"��@f�%Xv�N��ed��xK�~V`�cԛ��6J?zd]&r����ɴ��0x�b!T����т���zc�A��4E+C�4(�㜚e�k�"���l���ߵ��J����5yL �
U?��@OMr���(�NN _\F�Q�+�R
�Z��]ģq4�6|��ۍ�p�hw\4�`8���(�B�qCt�8n:J]��숍��"z�br���16>���i�-�+jB��J��D,)k����W_#k���9lٲ'O���s�i)�NO�^aŗ��m���ާ� )|M�B^^�2��?��Hȭ l��FP��&��@�׉��H
)�H�|�CZ"�+�e�tQ�^a������F$�oR�,�����J�<��Ka��乎�o7��ɏ��4+��\<�y��l^9	��ӜG�Y��TX��U�"_Λz?�+�Vk(Cuzi�����������`q <���c���6���u>��`T�C�n�y:��v%��[���c��:>��O��`�R���t�4cC��>��X�&1e%<��W����aX�� �o�s�՟���r�7_Z��aԪ�9,	�bӨ��3�}[��7_���)���T Oe�\k O�s�O�:�Kˢc�- �7P|�d&�*s�LI*b�L�i��`�y�,.ѲQ�tU9Y2�1j!�븨���X��Dc_2&�0V�,G�:���T�M���~��FM��,//NOcfb^����b�g _��gP\��#G��c��j�����<�XOF2.���[�؎����[p��qQ%��^,㙟=�'~�St�6
���͛�����"��&�9Db�[e����&F#Qt�u����p�.ݴ^���o{.�	�T�v�r�����G?�q�sL�'��@=�1�k�V	��Y��`г91�/c!_C���{���:Dȓ��)J��\�E�=湈G]Ѭ�&��lH;(G�\���ii	�A��E��	� 9����e��M0^����
�9"k`! �]�z��O�Fٔ�6�C�i����:V!ۭ�ٞ�O�㔪���+�	ω�����.�B�V��j�k�J�#�i����Kϥ%��]��g>���S��/!�K�߱�i�ŗ^wމ��d�F'�8U#�:�*x�����$Y;���X<��^�;��K�����H�-V��8\���H��56xA%���L�-j�����>���|?W�aFV���|\�t�g5����AWp,��s�c;|�V��b	��[���#aE�n����M^2D..W��7�d�_�pҺ2u�"`�*���h�vI8Q�%z:�%^0^u:�:v��a5Yg�H�S���>}W^w�9V||,��I{,��$dq~gv�hV�<�9#�l5�h5��Wk�aF� �+m���r��iR�"�n���I�5Rm����	iJi�
��'�7���H�'�$E�`Չ�TNB&E#�2M\�Nf�튀�;6cin
�"f��7Ծ�q�x�΋E��
�G�`�?����@�j1���v<ה�!p� �`_?~�Wuu�
��wޟ��$1N�>�Z�$PO#�{���a ~<�������	o����±Iǫp�_���{
��S��x�����:h:~�dU���%D~ه�Ϧi}�q���p��{y�O��������Z݊a��s�����R�ͷ\��"Qau����������x���'\Ю��hG#��u��u���H��̌���J��h�L\��:cPb��pvn
}Z�����ۍ���b����X���$��H$�B�fI�7���[� ���[T���������XZ̮?��O�?��ق�͵+5!B�ŧ>����y�P�5���[���W�{.چri�޴�������<�T8��L�gl6l�,@�X/��,9�j�*�|yE6-u�Rչ"J��f��o�����7^v=N;*��ʝ8{�������#H�"�eHF�[-�K�V�#�B���m}a5lX^��6���h�����[Ҳ�E=x����*u5���#��	�y$7M��0+���/h���]�6�a�>���	��� ��^#��Bc�E^�D��,���R���`�2�@Keh����T��~|t�Z-	H��f���� T�4(ԙ�� �毞/L(EM�\%�@B�~[8a�g�L��7F�?�o�7�x�M�����(csC&�;ڏ�8�;��,�=�n:��A��*�5�P�c��Y�k.}���9������w�m�^��3E�D��בHΌ�L$0�W��,�BN��yJ���e�|}�V ��T2#mGm�"����뫕�An~    IDAT�/�/�����e�>h7i@΄,X�ꏐ�A�(U8&N�9�B)ä(d2�c��eM�#�an<7����
��O��:�ǥnE9vR���ʼ kgV�%1�eZ�A_/ZuN5Vts*�	�T{mGbB��{.݋��Y������qͳ-���zc��6��Z)�#1��,Ȩ0ONW%�u���|ip"�oHŋ�I��@��L%5�ʽ����rurY���S�4��B0Z����;�t-t}��i���"bG�|Jy=ms��*��!�0r�FF�ѬḦ ,����z����K�y[�r�z�*Y<&��0�&�bx�ʬ�U�Z�*��{��^-�y�=N6�}h�I[اX�(��kT�<��m���r`�����h�0��kܛ�D��$��d�~���k�Z]	ӕ/��+���ۧ�O����5?�F���ݿ�?_�v����;���wu�{�m��RD�b�]��񘀰�vd�7��ɣ荘dB����J�\��^t㞴��,n��l5!��"J�)VP䂅$5y��Ѧ��K��ʼ�*�R��L����1(���3G����SXa����TM�U�����ģ��j��?8<�J�&����P4��h��T>�v%:�X�\�q�+�>:��t ǩ���ѣG���󥢜�"�@�9$�v�n��M��1�	�f��<��Ν9����X��Q�[�)��0��{.���jK@�8zn�FU���b݈T�"U�f��.�h~�ַ�3m4kM��<vz��O�/�q�d=[7��I`���z��d�7��z�,7��0�m�'�5"H5l$:�hI�=@�Ժm�ṣ��L��-Tx)r��C���4?x��ኒ8�zQ΋�������'-O�pD�;(���td�����:����DI���Vغ ��ƙڐd�B�"U��B������X���r���)΢��逤�K��� �7�}I��0���J�����ݧF�ˠ��?�I\}�2�5<�AirJ��Qa�����>��=�(�Ԏ�Ƕ+�	��Y1D�I��`��(�4���>��h0��(��DkcmV(&�Lʵ�&����{��c��:Gj�Ӡ��dڤX��EeUeY�ZW�
h�yp���T�  �����R��e�@�O�Yƍ��]�'X	�5O�(igO�XYF$B�����C1cj.%�I�x�#�U�#�$��wg�U����-�]RP}*����k���O=)ߗלSv���H�ύ7�,U�cG�J|$����yҙ$Z���;N�sj�U�J�^E�������ɭ��* ƪ�ԲĜ;���Y��,�V�!�@�Hm�:�����������6 �Da�t�`e��0W,�h���$�FP�e���0��dG,f�RX�J�%d{[�bi�1��iʹ�A(�A˯�Jt�����	HU�f�!3F~�c�瞓5���_��_���Ӑ��$-�8���וs^[��i �c�>�aP��1�w��S��h ��3�z����X���Ճ.:~�;�w<��	���J_��W�m��ip�}r@�0� �/���Ŀ�Z�A������������o쒎A�X�ѭ���1>E̝b��q#�>�4�Q��-�\L�A1�@I]�Syb�f*8�!O�E ��*��̊�Bbf(���1(+E�Ucm�/eZ��
�#�☮������*j��z�F�J�/�ŕ�/o�x2�r�&U��U�A��b��m8~���}�XX���,�[�˸xx3���<��[��.��/���S��ɸ ��Z��+�@*��P"��C*��[������2܈j-�8wFl�J�b=�h�nD�1,VV�B��!��,�ʬ����S���]�]�#�
41`f��
����UǄ�"�`�Q2ꠣ�D�T@:ѱ��r>ur����w�:��x�{�����EU��7���׳����+d����m�j�k�(T��X����{;P�K���G��t����0>?��D��6X#^ �5�A瘟H�:p �QL.���E�l�U�`��(��!��6x��T[�"E�8��3w�t#8�7��4ã�j>K���--4��td�N�4� ������|^IC�s8�����\\�����-�c?��&�.��ߘ"c F����(�c��W�o�SQt{+�:)���0�xXtp�^?�i[���J^�}RE��4��(/,&'���F2p�~����W\x1��8�{{�yWj�� [Fo�k>y~��#�W���u�o�j�Yr��pV8�J`��O�#u?T9����f������M�bd��T`M_w>���x�<w�	�xL1^6Y��yޚ"� �@R��b7�+VȳР�U����L�M�񢗑,�%y?�>M�̦�ɸbTLH�ԬjF=����!��)x��A����B��G��@&[�7�&EI�|��Eґç@��*� cW$3)/�LOO�l�0�/�o�σ�p�t۶nK�C�����5p����ѧ�@,�жi������dR,#��?�NͪF�55F�F^�A����jvOQ~�Z�ݑf�8�[}�d.4��5Cz�rQ�6[՛��tʿY�lXXHʦ���4KJv�f���O�%�,Jb�����kU�4�'��Q��/ݺG�>�z9�R3�r|�:�dE�Y��xe>��כ(V������|FZ�,i�x\�g��8p� zz���#�-[�7���>a�L�%�4�ћ3]��{�����n���SA��G:��㌎A�@�צ����3�
p*��~O릓�����P�5ifPb�Ei>�S�� U��{tu�"�S@��sV��V�����L��@X��0n���n��C_wG�n�.�H��"
�i,[��9�m���/Bv� �|.���C�JU.ev�{Qy�;+ F����}�j"�"�ף��4mi�{������T/��]���=���7��d���)�LGr�dȖ��::��{K�!��;��b:�t:O8(���}6�oHR~�9�b��W��ƭu����X��c�-2��62�(�F�q���'�\j^v���Ɓ�G��0[�
[�ynҕ<�5�Y�
i��yD��e�Т�Rnh80�D�#�w�+A*����#���eS8>5{؋�׆L�$`����ǟ���� �B�B��X�m��j�(U���
,sdşMy	5,����C��eR��J2Qeggn7t)��򻤻�E��(���^����R\��hH��	p�UYt��PAKG)�J��_ZF� ���R�1�-�8Zӓ� Lο�ij_�V��@�LL��/V}֟�0�Nx����U�5��&�������*���N�!�_�C:�ܻ�q��h����G��
0ǳ���.�gxvf[���d��n�,�t$��A��$Aݥ�z��I����%̣n�M@�s&���lص�� �$&E?�ǤҎB� �#&�J1sA1qR�,iQ/4p$s�/��sl�|6^S(�R����Ӌ��ǆ�I-����ZÖ��p�Y/����?���N������8x���:b�2������3�°.d3��%��d��������ދe�K�������Q*���T�w������'W����w�K�,�SO���<�_�{�-l?�l<x#�G̔'��V������96�����J��ŮOj��)L��!2�=D3<z~�Y,�l>�v*�l�m�M&�H�Srш��"�w8<�V�wP� X���J��ZY≌c�!Vh���زa��c:R1L\�T��L�*<��.գ�J��V�>ﵮd|����ݺu���ɀqL��O�׽�url�O��j��ʐ�t��(Sj����AR+���Zo�ZA�R�?G�0OW[�c3�@���9��Ws����{�X Ey�L��3��J6t���U}����ٰFØv�|ߴX��{�������[�{c��;��e�SX1�߻�Ӗy�7�����^�yp�Y��IY۬h���G��Y�8���.�d4X��=��pI��0 �bQ�����&
WM բ���{�f����礭^<xh?��N��!O&����fi�z���Ŭ���z\��1�hw9�|�Z`c�9i��&�4i��g�H����/Ҏ6o^��t+���G���>V��A�+e�Xn�"���Dg(�����<�g�>~�xRv��F�m���q8;#X�e�v�b�#W-J (׊����������Q�eAa6��H��Vgo؂6�ɹz:�0��cza��A�f g���`<5���!N�F��R�(���tN*A�l�
��~�aG���b��H�nk�`���XF �vB<?>͊�U[S�j�i�m�D���]�	Jr����r9����sq�8ء��6�N�E���c�'8D��D^��c�`�I�����Q�/�
�*8�@�@�A�b�NN��Y��	n�Չ����@���Z��ʐ�4�/z�+Ph2a�E�	�M&,�J(�Q�t����K6SS�L���P� �j_�'3�,�:�킿3��ukD7�*4P�䐍Ǜ�|����h�IM�Ne�\���ML����t�P���	�7n�(@����=|"6�*ƒ�D.�d�+H/�v��Tp,�O�oddD���80T��fbtL@�k�u�T
��P��D�M3f��c��J�$��f'ƐJ��뢵N�����-o����\��v���CC��س����:�b��E"���� e2	�0�kXlnT+���b�x/+U��u�����Uh�z�������
���t��\,!�%=]�8:t=�}\ևL�
����_(�����Sri�A/l;
������b�uf؍�"}ZU(6�d�[z�Rv��D;1s5�R�f�9I��9tRA3}iX�%���}&3,��v'�{�����n;P&+�t
�KfK���6
�$�Bnt�����؝@1�*�"2�kMX����	;fz�i�)_�MOk�n*9v�ʲ���?�l.��kժ5�4Y��)�ʦ�xz���������g�̖f�ylv��OK���uT�0���PQ[�����>6Ǭ�U�%~������3{��8��.��Z߭?S��V�X&\���,���0��
��b�����z���n	�n�c���z��8V��#�O`�R7>��ע01�`��ŐܵsWᲡT-�^� Gӕ\݄�4�ƚ��y�E�,���b/F�����@&��χK���]"���rV/:2�[w�G�@��{r�Օ������K�"mth�H�Za����*ҵ�Aib[�aad
�C����ۜ��~��b�����o}�Pm?7���%Ț�E���]�6�ߺ���J��r��B>�XAln�?�fr)MN��&���Q��s��!sW,��b�Trdc)�NL�%�7�6��?v6�����a,���C�f��ׅ��w�����R%���dT��:<�>9:��lȗ�j����J!/v�X�j1Pci9�u켿��}�+�ߣa��h5�}�ǅ a��r;e�Y*��IU��Q@K���Sūvitw�b멹�9���L��b�����sl�Ν�o�Xz V��Rr:H)���sj�Z�S��J*�-f%9U�7��,�q�OͯS@�CC��N�BY������6a�F�G`�;�r�Q�)͓���9<���J��t��@W���vzð�kp[�C|�ÇO��엚&���?WZ��8۷�E����}���/��@ͤ����{,� �ѯ�y��c�LW� �����g�ɦT35�8a�Lk�)-f��jQ%#[��QR)�8S��y^�T;�z����QdS��^+�p�9g���5�(���q$RY��̓p{7�-[�J�A7=䋦�l�(���X�w½����$�N�*����*�oXJ�����Y��r����J���Q�y+e�[H�����ϕ���p��Ã>�l6/��'��jF�˺aqZ$�Iְ^�KK�5�t��qT�Y�w�z���(���w^C��T]�>�����j �)H�jSc( ���a��`���D���n�҃9)�'paz������ �`���Ȥ����8�{8�50cV���z3%?�% 㳒��1?���C"G�-$0ZS�P���,0ӑ�(�%�a ��� �7�k5�[찰��ꐖd��J��\�b���f�q�)D'̶f�h��I�f�ZS9~�{�����C�OY�����ꭴ5��^�7?�����F:����]����y~2?P��`JUl@�ҋ�q�L8^�8�1W�{Ɣ��4`�����xۓ����a�m.���tGu#�p;Sj)XKc����	z#�:k�*���l[�`C<e�a&��.��F���K�7;���HR�Ʋnq1V�L頯�ܺE��`au��<얺`�������_>�ɲ�RC	`Y�l���f�V������h��	Ha��v�{{�c��bJf�P�"6:���hs�`�=�ʁx�[ފ��.�ݽ�w?ƇNH��|)���y8=^�\p5��{�X2Ї���"�Z���q�:��y�|u��8|}t/_���Ȧ�
D8�9Y�X�3z\��������@���{�|9V�,��e�D&V��7�<�u��h�Έh�\3��GF��e�Uj��:P\H�+Ԏ��-���ȳ�%�&��̲0'mq�]*Z�r�[wn��۬���@5Y��:��n��U�t���.�WL�p�|	�|^�V���.0�����
�a��N������W�qUŗ>W�pҺ�RKB�~��T���#���(Y!mi�,�[fJ���tuW,σ�o�LBҲ.7>���g�vltl+�hP8CG�V?>�G#�/!�F���\10(-pj�� �T*�R���5�Zdl� �)k2(d��Ʊ+�V��q�a?I�Gk.����d|��ɂ�ؒs_R?�����ɫX���<wǢ+?sɒ%�T'Q՗��4�6�<3��3�?K�On��G�WjL��R�D���᭑�7����j�7J�$��sOǥ��������ҁA�u����[*WD��C~�dJػ�����**�+Vaד��뾮������ֆ/\�9lݶ�л|��A{[H�|��L].��w���f���}]���
������~�;�������G�7�J"u�� �l#7�L�xR���P�\UڗF��,���Y�����>[5n�ԩ/�K�6ǔt91�?�)��519��H��>��������C�\G�T��B
3���@��H�Y�H
d�ZQ��VB�mE|v~�S�m�7�~�L��,
ϙ�����!``i	�g@oo� +���'��'=���zl,�P�C����|=�Yb^3�jx/�Z�<��\�Ĝ�B
�X�%L`��W��B)��h'b�y���p��Fq��Q/YjH-�_�T"-]���Ւ�o|rL������Iu.�#_ǝ*A���ϙ����5�̍?y��?�2II�sͧ���G"����
s��D���O'����L��tu{����W��t�g�Ꭿ����O5�}�^0a���|�����oּ��U6N6�D��a�Oa��6��U�/ Ϧ$x��6TsY��Z���G��ԩ]�JGrW�pyqq?(��ܩ�S(�/�
�j� ;M��4%`��f��ø���1Zta�d�砎����L<�Y}h���cw��1Џ|E5o�yyj�����ؤTJ��T��嬗�-������	��-���a,w%[���ԧ;�¶3� ����������W�Ы�É��v�/�sU
��L�RK��*�N�P*��F�P������R_�v7�|���30еDL9����˗![.��!��%�������WmT�J�X]X�хz�*���|�l�CX)���V��\|ޜL:��'ت)�%�8�ʴ����Z-e`V�
�'?e
o%��.��b��45`
imP�PRV&3��j����Pͱ[ǮfYD<�&�f��_a�#M��`L����u�MK%�������f��6K�~��;vT1aAAf�p�W�q�'��r�\(���GچY>r�R�
)Pa    IDATu�̘�$n$8=8��^����WUm�te#�(�0�=W<��l uw�����	��
��Yɸ ��N�vJf�:�����	*��@yqM���s~�jXI����>�+�]y<��daL��9M��:�N�S��=G�y�=W�ZA�`���l`~v�t�M�4Jx��o�_]�:\��/�e���W���;����Awo?�bI�3���E4�&}@������#����yU��}~����8{�V�ٹj'���+*�+�R���y!�C$�e�:HZ1��P̂�g�ݏ��D3x�w��G�( ��2�>���>��W�� ��% �Ҳ[�i䗾�|V�흨������n���d�K!�G͋�a
�x+W��.�}2vK�.Ömg`�3097���Ǳ�g��&fb�ĺ�D;�D;J϶F9�QG<6;dӲ���](s�PN��//uY�=2�n�$@�c��hՊ�D;�� �֘�
�T6%�P,y�i�ڵK��E���矏��q�;7$�"�^�gn#�0r9�]��c[UP����P��E�����V�.���	yY�u��	�=t��	nB�Z��s�!��i=7	�ue1�ϓ 3@̿��nZ���rN162n���O���3�*��u96S����KutP��V�=>�r�C�]7{^l�|ތo����ෳ��F����%�,E�k��^�@���5{iQ�a�}]�px܂��x����jz���fCQS��zPe�|0�N-DV����C��?t�&@�6�8u�ڵ0JE�CK*�N"���{7��M&�Ϙ�d/+6���e�9ȊX��ڄF�Nַj�jWD[�J�r�xB�Nfb
��K�5��R���q79||�D�R�h��5�0J@�+�p( f٫7��+h���4R�4�=�\�{�@���e]�e��u21�f�X@2�L#=Cblv��h8v�d�P/Cp�s���0F(��d�*�x&�d6#��z{��mX5Wƚe�(���:�Z�&�_)]P@�.�Q����*��f�Z�j�� ����?L5;�3S��c��a�� �4n6�6�N�j?}���A��ZK��*��N�/2a��x�:��SZL��d�0��xOx�r=�ɒQ�A�B|���"8�/��ꫯ��F&�i@z=��-��9zBGI@�֠��]��?����R��b�cQU�� �i:��G�&j�LƋ���EIWH�a%���P �?��S�ކ0R��0@���sQC(���3VpA���������u�<��f� ro�y�#NoZ���T����	Sv5T-e�Jf�5H�x��*�4��2>p囱��3p�n�>���vt"����g!�e
��.��6�Z�r��h$�x"��Wb����/}G�-T*�L�p������Qm40>>*�h/��o~˖"67���.qi_��B�!aF��Y�;ڢx�k.���Z�ځ�{D�B.ޯ}�q�9���_�gY�)QP�k�RI*`Ԭ�#+�Һ��TVZY�����E���Ǐɘ���g��R��7��R�	cOG�����6���ɏ-$p��q�����>�)\�W�?��;�0O��}��u���P��6�qZ�lT079
/;zs0�+3*8t�F� �M���p]Rڶm�6����YI�v�ja��:t����Ue/�w,o6�����|@���q�S�gReII	���kO0�p����i�7��-�>?���b|+~F���g�g�9A�X�C����lbB����s�H�,�[��s�{9gxn\S�;�A�i�-٠&.
H#���������l(��5tjs�u����K�۰������F��%�� ��w=���Ϳ�X3`+#�|y}+���t���!57�Z./���j�x%v�iUM�l)�7�ܕk�k��h���R��ү��s�R/I
�QŖ5+�޿��
�4i���\�v~��A�r�o1Vrc���U���4�6جB��0�ހ��	����D�'Ss\8��{V�x2�����_��p�����-�f��N�"3�@y:-�2���M+�����6>�³����JY���@�@|m���(�����-�]�+��,T�r�ҳq��y�2z::����O (�81��Ĕx��9��c�6�L�ٹ/��J.���=��,�Ʀv�a�(er�xCM���S4�|�&�IC<��h�('�f´MK�	��X�&#ƴS/�Nj�L��b� ���gS#h��o1�߷�d9��[l_�N�/�#��i�G��f�;�*�7��Na¸eW�&VyV%95=.��Z]Y|���4���(����fU6���9|tH�!�<^�֮�nx<>�=~��ϗ2\eK��u�'eP�z��
J�[S��Zs7�v�c�����l
@1���sq�b�k���;���2u{y9&&���-�j�x.qv\���p�Q�q�����d���4 k�.��|��x�J|q�_aO���
��j>{oy�%x]��ݎ�~�s������`v7{D��;�DFD��
C��0&.�3��㟾(#U�*3j�ǫ.=O��}WHؕm[�`lt��NA�X^�332Zd�v?�4�c��m\�7��uD�~є%�i����{�n��^����R��g�R�
�0ۯǫ���5�f��D�xTu3����Ϝϒ�4�+��M��b�U�>�Lb!���Uk����{�U�HA�a����M<��Y����"�-���a��բ�̤s�����ܒ.��N�%� ;�(3v��Ǧ�&n<y��Q�ܱ�&77[�����>�_�@XR������Ās����F�� ���� gϞ=�CȖT)��L�q�����k��� �s��m����|6�=���5|�jC�W]�στ�����y�|֏=���Y��|�Z���t��F%��<�n���r���Z8�x�ody<Ͳuu�ȵI�v($ �ϓ�����������n��嫮7#�?��;����#)�����f��P��a+�#�le��F``w��h�a�E4?7czu�P��K��e�nNv��icM�(k!�Z�+@�Z�	K�f��R�-��Y�*L[� g���A|��(��(���k���,N���A��/��MhP�+�\� ��M��ᴱ$�	^'7��ތt}玗�O�|��\�����W6j�8(�V��g
���]�Í�-��d#���'�êͫ�nwa6>��l��9�5���(�z�tQuX�p�YpZ\�9���|<unܭs�x(�,� �˕P�N�L_"����.)����8r�x
�lǇ%������f�K��f��Ax.����z�	̎N��A�T�4��t���Q�E�M�ݠ�[da��#���i̲�6M3�[�d��������������K*�J�� 
�)M �M�%��'1`�q��U��j�L_��&��ӑ� L�T��R6{H� ���R�&;u����3���6���������a��i&)���U�ٷCǇ����Y�tׯ� �V���͓������XmG!Z-(P&���EL
_$���S����LKZT��s�`@f`�e���La��fz����&L�$Ɏ�*Ѩ�G����A�L><m����i���1���.������a5C1aԖ��f�Р�B)��ǂ׾��l�����?|��X��_�~�h�jw�����;�!���B;�D")�HM���'�O}	535N���k����t�0X���'Dϵe�6���/ �?�_�䳠� �S�4��lN�V\�Ob�@��F"۹{�[�C�
ֳ�:��ܵx��]��7��I�G
�E�n6얢1ff�J]��Q�J��9�(X��s숰���![�9L�̊6ꪫ�/����n�|�{��BǇGн��*p��F���D���06>7�Nٿ��b����Z1�F��D|N
}X���K���N~�¼�����FwO��յ��`��A�G����hU+
��Ar�q��~q<�M��$��P+�q�9�1JM�-3����z���vy�}�\����V��E;�-��9��dnN�&sͨ�	�8F8/������&�JYL�9�i��c�M�,�Ȧ��3A�4;F�~|��}���P@�, -Y�{��s.�r_������������F�a��O��w���`���
iXYd*SX��5o[^ZA�I������-�}Á\� ;i����%b{���z����gz�p�18Hr%�2��~�] �����>�����E���ˮچPX�zp���L�u��H&�&}��,�RdB��*aS�N���"�&ub�h������b��q�a���:����)�V	�Uj����!?��'��t�3����p��1��!���h~D�m��?�C��C�f`>��a���3������XJUTrt�B��X�֋J�O�'V,wMB����.L�ĉ�B%�E��PG�nƖ�[��v���c�K�c��g��M����\>�SlM ���te��@�s���X�Ԡ���n���GfS��b�t�L�n�CR�Z���A�A�#���\�*�[A�E�q1�R0��ϙ0�z݀�\8y�S|.MX+�ө2�;I��ޑ�~7��}��1�͋Ɔ1���=�E��jM�=;	�d�-<��.=1
��-j����N۴E�m�]!���	|ս��C�."0�����;]�Mt�炰u��SSr����<�"Q;v���FQ;�L\�@��r1!��5��������	�vT����ul��x�Q"�%,�Yh�65�-a�?(�N,$�a>�Z��^�����X=8����g��U������>؜>��A8=~�
e��y�<~��81,������5k�g�a|�S_/,j\	
hwpݗ� ǧ��u��w��\|�Œ�{��������z9�.Y��x�Y�	��?���p�����g����؂;~���y�w�޾����ص�I�sDQ|��@��2���ݢ�-hI<�����Y2�yO>���Y�0m!��:n&�v��!��C�P��o�����'auz`w{Q7x��qXl�D.��
��/^�z�zl`G�%ZT
I�4s�_5�]���<�������
�����O�$,�2��u�P�!�����-��?A�7�I��{���:Yݭ7{����ѭb��VL���g�_X(@y����s��F;�͙���vc~~V2�^�A�MY_������#x&(�q٠�ϳ�w�X�P���)�:�aUr�hǎ����x����d�Tt��M}�~���A$��48�:��7o����k���c�m?z��[����\��%v�.��F
��$Vm�Eŕ��Q��n���T	2wk�zAZD������K�� ��|�,�� '{$m#��$t�ܺ���JD�
��"�h8�q�om�UNcY�_���a-,�(��ٱP^u�p��G�Q��*�f1��^;�n�JU��)�|nt�����>�dV
&SUH�z����y���1`�><�S�G�;��r8��tG��x1�y%���%cH/�qp��u¾��t"��\.%l����X@��U���c녻�-��Y��Gfz��>�.���NVa,6��K��Jٰ��f�'��W'H��f��G�PJ���V��e���l��u`�uH-�)��� ´p��ӁJ-�u	�M�J�d&0 x�b#�>���١~�]�Q**�ǘf0�b��Ŗ+'���A�~v
x-�К�DfŰΊ��Q�Ȕ����ŠUt�^���ο~�h	���,��y����������Q$N�/���7�~��ˁ���!�Ҥ��s%����LA�Ī2����u��bjzӓʗJ���0eL��g�UF. P�D2��Y C���`��@wr�3���D�r>\�0_���c��K��	´1���RG��~�u��uY �<R�j�P��-��۶l�#�K����>H����Ui*=I]����б�
P���-���ŗn�QґdD�5V�eq�?_�W��e8p�Y�u����>�O�D|��m�݁cG�Ij��{�p� �\����%�]���?�[��&\���pιg��?�����.��Mشq>���b�3����p�݀6��M�Ԉ�QVi0�7�N���QE,�&s�m��1K"�Q����6}�Qd����_ ���O$�]v�e8xt'���ʔkC�P��{���X�#�އ\��b./�|��c�H[�n�d|�vQ����ڼ�_,WlN\x��b��L.����زe36n�  �`����
��5�d}�ܴ f6�9K�bV�*cZa�L�jVK�>�5��AO�L�t�j�A.�f���숐ʈ���N�w������6
�=��p���t9���2X�jɸ�Qkk�!_�I��W�5����Aj�a���8JŲ��˗�Z�ϥ��켴��qx?���|�u��_��Xԅ:���*�ل-�z��xfW�{_�����|� L��p��Ç}����u�/_W*�`)d�F��8V�ދ�+�����F��b����lz�bJ������ M.����ܕ�>�*�e�71K�
�KS��p�����'>�nX
1Xk�ʕ�_�QC��ǎ��AXE�Xj��06��ܷ�;E��귂�`W���,QK��Hk���7`-�Htq�N��[�A5���P�K������5��TC;��;ځ@W+6��-�Ĕ�S8����"�0z�t ����,
l ni�gI��(��_w�l����J�(��!��'�0sh�JC�]�O⼳�p�0?�w���pxݘ��ap�ji�44rB(�@0���Kaa[�j�D�dF��zۻa��´��Yl3��
3�����c�4�L�Ӏ�	����7�Q;�.
lnSI�6��I�hXX�&��-I�'�f�:̴o��M��z���@��C&L���u3+u1�Jߛ�5������;Z�#Gabb\<�V�Z�h$��/V�a��tWWn�N�8���iq"�����B^�I�g����)qݚ��л�;�-b�ϛW��3VBZ�$�����>��Fa��&�ˢoI��_�A���z�(�a3Y6|��l���T�ͧ#X�f~���czfR�6?��5q��bڄ�6Ss�"���@b����v�zR�J�t�=j������f�ת�?��Lʅ
fg&��r!�K^vV� Z�%P�S�F��պvS�^t� ������P*��-�Ic�����=�­?�Cܞ�֐�)�W�v�h����K.�����rC�{H�qrr
�����K02<�;��k�.qx�X���zgo)^��Kq�]��=����o~+������g�뙧����VRβ�1�Wi�*掦������:*��e��`\6�C<����B��A3Je�R]y�R�w睷����կ~5���f�b�W*�u i�#;�����ű�c��๳ۋ����ހ�A?�lV��:%�
On��ib�j�
iO<+�&�UU����M*��X�/ L�n��aqÐ�<e���X�z���%
Sh�0���Y	�$-(�`�:a�kF]WGr�q���H��z������ۺ(���ܴp=֖0��sJ�{�l?�_�M�x������	D5��ߣ�v4#�Yg~�f�fj���cq��@[�[yl^����s��׹\��È� �K�e/��	��'�����~�u#ܿ�� �O�QK�X���-ݨ��9J�9������hԩ-`�<
��f����rPP0-�$���Y�J���q��]6}��qk��������r�k��,g�ii>�W���G>5�XhO��*���;���8���\���5�����b�W���AVfu�0�z�45A�B�$?� ϛ�}�8���,rٌ<:G���P���g�i�-�{��?1��}��;пf��,�+��A�\
��G�ن�7���%p�����2)l<m��-JՐ�I��1:t\��ڻ������a�.���4��>���KP-��[��n�.��869��g�=K���~)���"�f�2k�L����?��H��"�!r��yS��4�i'}��    IDAT"ϕ����	c0�~[H��J!Y�iDh.~����k�P���M��Ё�LWj`�C���4v5w�L(�
���T�hEL�ݪO���{`T�[a�X8QUl�b��ԙl�N�0_:��k�1x>M�Ƽ����i��d����czz��6����W��el۶�x\�St�/�;7m����w�U�����D���/����N�"LXr6f^h��4��HF�d���Y�⢢��6�*� 5��⃯!��s��38oظY���]P{S-��Ϟ�4�WMUFƚͷU4*c�s���¢��;<k�/��L;��V��� L^k�s�VU�	D'F�0?;�J9�����mY�}��/���)Tj� ���	a��-���#�/�-�)c��^~����'��>�X�4­��}�_����?b!N1�=��`/��YDW�Z%����׳d�?s�����Oᓟ���k{{��9�å?�W��b�������հ9m��{1��H�!�)�7��1��.���=��Q���N+ӫuE�s�1�4���� ��Uc	��moƦM�p�]w!���=s&ggp�;0;��+���?8�щy��ٰ��%�~2a�K:�Lw����З��T>��aI�/�f25Z콚N'�N��Kʖ_�@e�L]�i�,�֕73$��3���y��l޼kV��4�fxy�O�;=F�Ѱ��� V�_0�r��}*�Ym4�{��s�������z�Yz�����������%��d���$A�����S�QOǲ��	5��ρu�a5��5��0�s/z�@5a�v���߽�7߬��6V�~^L�Z��T�����+�-+U���<4�s�Q�dQ�fa�(�Vq!�-*�9���>8b��ԠL])̓�i���jX����*\�.x]N��
��ƪ�0>�����RB��
�k�Y8C���;�_=q�S@�BLmlY�A�(zDH�g1k����k\�]9�uF�)�EOe���ۘ�H���0O@�gy3+��9�҈n�P�y�O����ܴP�m���1�M�>#�߉ޕ�p�XX�Ev>��{� �lGg���KQ�60:;��Q�'���ݝ���t�/����~�&�(�r�����֗���Ԉ���,��d,&,[{l~F�'������d �5QO�p�cw�3�%-�x\�I]�x)�/q�rQ*#[�ޟ�'L��O���-B����hL�%[R��r5h�g������0�B��&�%�Y���YԊ�]�H�㨴�"���M f�fy���� ���
�tP��� �VEa����]��Q&��S�����=�s����2~��y|��Ǿ��D���'dW�q�zy��d�	��u�^��a�ZX���m(05wl<��*	��G��RԌ�=�Fa7�h;ɕ�K�9��$�vVl$m�A��p��© [UR�d Tz3';l��4P8ul�4�d����J1���a��B1�\M�M"�I�Q'kQ��z3^v���G#�_��Kр����T���wjU�	;Q*���D�Z����Ń�����	p�m����q��>����|j'I�QDq���1yn;z�\��1��}W���f����E$�!3�����go?���lټV�QbCQ���w��G�d&!w@k���@-����̦����֤�]Z԰�c]m��(�IC蚌�q% �쨢{���<�igZ�HS��q�&���L�t�w1�Ƕ���>�?�b��ݍD�]5�����j�`/��S��uަXp��6M�ucz^�4r^�&�(�ρרƒҗ���ju�:L�_�e��A�^��K��� ;��(3D�o�=
t� I3I���|��|�$�j�﵂:���,@`�j�Jo4�n�ha��UA�b�U���YU�Wv@Z{�s�W߹���i�7_/�ٔ���a����%��[���/Ff|��t���Upvl&���hT(c+ք��f�@{�r~"����,R�קʒ��
JE�-`�
�s�d-�$���t������ۨ����y�K4��pP�O��l/Y�o��Rxl��v*���E��H~p��q���q$m��U��҇���%��%��A�0��-�06��y �/؟�Z� '�������6�E!���3�K�|:6'���ŏ�d�c���Ï�����)=ñ��p���ً��#�׉��b�6]���3�k����a��*iU�� CF6��o�=�6̎O⇷�*)�c�������H{�D� wЏ��R�t^�ζ8�6x�^L��R���*��rKM��&&'�Ye�@`͒�@nZ��fU��zԻr.@�G'�F�ˈ�"e���A���|�
|J�N]��^�8Z�8ٛN�t��fAR�&�Y�5��z��� L�3����0�eb�	�( �Z����w����׈0�0g�'���EŔ����OL�����(SV�ϋU,�'� �*�Z]��h�T�h��1]�q�k'�6L��/}�+�?�#'�������KХ���	��k�E�c����P@[�X�9%G)�E �S L���N��ܤ ����ry�l����ʄ�q���);��Ud��d�N������$:{ڤ�a2�AO�RX�.x=a5�x�a��ۺ�ϕ��W[�sր8�S���ދH0�����}�����[�%�j���O�G?�2�4^��W�Yr����Çp��a��ud��u���\��o��P��{��O}�6�E:���'�(�袋$�{`�!��=�Ǉ���M�U��S4��ں&�5�ik5�t��VI9n7���.J�zf��bQ����7�CΏ��T��-�p��a�#!8�^ܿ�!x|��%KgỤۇB>T��]�	�1�M&�,"Dy�|q�n(&�	�أ֡�De#lW,ײ&3���a~9��V�5��oz�_���W���g+k�H��l����r�R�u�TJ�N�>j��ޙK����+ԺU7���O�X���������(�O�M�)�� qs�� V6�&�"��"��\k�4�졾o���f�lX�������0������������%�tﾳn�����§Uh�Z�I:�aİ|��3	�5�ngg�Ī�.�� ǂ�N��$Մ��U���K�L=��zgu�-�&�jq��9���q�c*���t6��ύMkW�V���^�U������;w��OƱ�q�@l�x�E1aNqy�	&=��td�=�4a���j�ܨ�Ĕd�$�K�6ŀ���b\�V/_��B\��gц�q�vG����~�jX�̌�`vxcC�p~��:�5Џ��z���Gِ�]1{�N�ry���T5?;�����辸��uD{���lZ�V@�C��P6[�e�G�Ш��\|�'~bR]���Za_P�=iM1|�¾�TT��y3tj𥟝�L�m3Ķ0R��U�:�uQ��R�Y�2ZK���sqt� �fU��@��Tn֪
O�_*�~V� �0���5������S��L�SS`��.��[]���!bqj�k��@�0�~��s�#i��s��&�S$&���_�7]�W�J��� ��Bx�|�S���3�5<U�^�_2  �M�*��� L=�S�C�	���3�묪@�Z�*������s3��M��JI�8
k.iJ�sYڿL�+b��i.$\��77xiԘ���*��d���d��3���突{�3:�	c�"� �tY#�M$٣cGNy�p� � ���7�r�c�*@��|��T��l��r|�V�` "@��O��)�Ҋ�֬���8>���������س�)�zj�����/�%�\�{��P��pJ���u�a�y00����;�I��&�b�_n�"�x�:�c��B|^2O<��<*P�9d�	�����9c��Ts#̿�>����0����ϟ����1Ѡԩ�j�H���J�rRm���@�+����)�?x�(.y��aX����=��ΈU~�J]�*h�	x�����ц��"��K�cA���u�PqLU+��R)>ѻ���Z���"��K5w��F�Z3���WHK�Ç�L��Ӈ�Y�㑌��x�8��|��J�Ō�K�3&�,�і����u�f��_�4t�^�r��(P�1Qf��2_+?7�_ZXk<?	���;A�-��/J��{vo���~��n"�k)�j
0������Up�k/�ڮ¬� �(�p4P�����;10s�z��I���(X?LVRZ�p���N���%�%6��?��ݨg�2q��Sa0`��P�}����C8��
��
��S�0�#5kՄu-_" �.e���шV\��d���'��&��~4��Τ�0�U��@u>���<���J��j��@��Cvn��s���ڜhx���}���ɉ�)xmD<AI=��
��J�r���|���}��6;��8��M�=���
5:gS����0>;�x�*D��72�H���
K�W��z��b�H��\�͸��������d@��N=�[uTz��h̪�/v ��b�T:Q*MWt���bA4�&��&�BG���EC1K�\��;R�O3S��k�:� �^j<6����P�b�������W�j���ڞ�����c+2a�O��j�i㬗����ł��y�\̦f�q��1�/,�Ď|�V�TkQ����#�<��Ү��
����2�M�h��~�s�"X�0��Cǎ�~~V���0s�<�lFYM�cE��Զ���7�0�t������xLY1E�ԥ�M*��uRz���_���
X���,���1�0AK�8XjR�]��Լ2ɭ���|U�
�ݲ3��YifC0�������+F�Ĵ$�� ���۩k�P�����{����x����>�T2�?>�;l�~�l݌_�{/�ch(��?�mo�>�{$�Y�\���1�r�M8���0KJ�+e�i�o�1F��ᢋ.�}����2��y\�N�,T����r�t(��"@w�]*]R�&�C20�;���Z*�@i0�uI�H	
��̶H���%K��R�wi?��s��կ�f�F���{~q�}p��8��ӱc�ܷ��#ظn%���Yo+[���N
yd�Q������g�eV����� ����#sd�[dLӮ���t�ޜq���y�#����#�d�4AA@�:&Y�5^
d��=�^����;l���+��W��F��"�i��kk݄��YoP�|ЩQ�^��\���V]�|�Y(u*�%L���ST\T �j5�k�9��0�W��F�a�׻�8�w=|c�ݾ��ޕ���z#�U+|�O�%�¸���Ó_@XY9Xϱ�=,.H3o���LUI�j�-����-�OP�",w��Y(ڕM�I��� �f�rT��څ�!�Ķv|���q���8��!I&G�ӊ	�ҡ-*�w�Ʉq|0juY�38�b]/�A�JY�h�Ij���dUL���
1K���E��@5�Cn4��B;�>t"�����N�P@�fA9���|�1L'sH4(�E�C�|A��L�L]�2�榦�zp�g��gnG:���󼙒a�y��ǥ���4LGnZ��1T�<�o/v<�k<��I	`�bn����8��\�ms�FA��-�XDȍ�;��5��:良ӆ�W�0�7�qsҋ��T��?�U�f�ZE�4����+�:STk�0]�ô�I�I)���3��qY�� ȿI��)�o��cCF��?�c��~�kP;�E6���0_1a|+e	�h.��}���R�ɦ�܎��]�Fwo/
��ɔ4��ؔ����2i�e��	�4�A�~^��Ϛѻg~�٪�J*�SdVo���3�S��� �lw��<�0]AF�%���]&)Ϛ ��S����9�9&�:^7A�T/�����)fF��O�z����4�=�	� �]2��c�S�hR���l�F��6�6���'U�Ǐ�I�qؽp�=�!"����X���h6���wZ���w��0�>'����'��`�+i���=юvic�/���ڞ�����WJV�O#�+��	��㢋.��}�j
Y��C�V�9����c�(�J\�/^-���-1��V���RW��~S�OY�%U�"��A6�U���ڴ�S<�T���� L��2tL��#4�����g�#�G�#�[�W�m��z�d�+t��`|:������������?�#��oz�bQ���$H�g�iC��;s���_�O*���`�U�'��b��dM@M�"e�,J�䆢�����0n��2���!1�i���+?�S�V��uA���t��OR�G[��Z;�*��s����j��%�ikP�5�j憅���Gon�	S_��t���_#�n�j5n���7c�����_� �H�����]��_>�oUǚ��l�]͠V�����mƥ����=�����ѷ�&M�]v�P"Z1�4[�P0-�,�o��R��$�K5a)'p�)��3��$=&�pR�<p�:�.��֍���.ܿ�N���T#d�h�^�x'�� �Kӑڢ��4AS��RQ@X�a66�=���T�$e�A��*͑���ȍ�"7<_�)팸Xv,mömk1�²N���)����͓{�4쨰I4�É�BJ|�6Ү4�������B^?�����z./��w�$ ��6���g�Y)��b��f��03;��}�xl�Ni���z�.ħ��p�es�������n�I�N:�Km����^�$�6���s"�T�]OB=�[u'r_�j��*p	{D��Ls�I�@���C��R�jǩc��"�haO:�<�~��� ���켜w�b�j(���a>����I竟U�W���d�9�sg�mvvFZoq�?��)=B{z��a�:�[�Fz�r��%��!���yn!�L.�]YN�G1,�2b}L3����E�S��E.`���t�xX�OR��z0>>�eJնFW,�	�$5QL!�]�=t{U�̈́�y���W�\�&#��l��xzzVޫu`��|e��NNI�+���������D1ar�O��`1������Ѱ�{B��:\A�dRe_�#s���ç@X��!�$�Ɇ��Tk�
�=�L��i=�u�ۑ�$�w�3ؼy��֙��E0��}�3�&g��g�/�r���+�����-�k?��>?v=��\s��.��b��Ȥ�\�m.?vX��GdD�
c�S�/�D[4��+ϗ��cMo�'��zCL>���L�.к��h�X8�|~�̃���r��?}��3l�,�K�����pbd\�I�pP�]
(`�!�Ó�=�{~~7�>*��9d�X�Jk	2ad���^���P��PX8��&�`Cr�γ�^Y��j�I#s�yy�7�j�[��&�(�̓5�����x��s�)�7t<��PU�z0���c��Ѡ�����5�I�~j`|h2_�����a�sJ2W��x���tu�)�9i��n�U`ީ�C���>�a{gf�w�8x�Ow��+�`�*���l�[N�T�ř[zQKć�v	V��貕�,fP�daq5P��P�T�p�1��f(v�?����/L�[(�Oi�A�K]*�ű�����%v�r$o.��1ei��ދ���n<��(F�u����#G�(�W�J{��Q��&F�2��V,Y�/�92aY�^)夿"igi�f:=3��#�	��Ϊ�J	n��lsϞ@y,��H7�v���4p��[q��gbYg!�Sڊ��l���㷿G��B��B^R\Vx�.�x�|�7o�_�Z={{w?��윤��~ו�̓�Kc�e}l��N��``9ۧԐ�d���+���b��(v���>.i���^� �ގم�%e�
�����H��e�6Hu<PK�	xOM��@�C�;5��V�)oM�����QmR$1"U��ހW�Pl�]?'��Y��9K�i��א^�<z���p�;h��p!`��bfG�|Nb'��Ea�~��:�
�t'�?��,)ߢXl�GNHi<+���9txHRd���ַ��5��T�rQ����ɋ���H�n�)�`���E�i�	D��5��h"ŋ�dƿIj��v9��d�:bs��F��~.�^S���8�Y׷�W�.|�/���=l$    IDAT~�f���O��z>>���.i<�ry�)J~�n���f!�s�'ap�-�>���	F�)zU�q9�B�Nˈ(���M�{��U]٢��*U)�,���Mp �`0�1n�h��t���19���LN&	���B���ʹN����k���2����w�p�O_���9���k�5�c�	�3�|1���dea�(ȷT��x{�VT��i	�;eP����D0����+�pL*?��S��S��{��-|��ֆup����~��r/�DT��/�"�J������u��D0T���.�w���X��V$�e��ߎ�����N=Y6��<�����Bqz$Fh@�����8x�u�r/�>�q0;�:�;�xdd��&SIx�x�X��:&�����"���2�1�����>�q�7�U*��.ߟL�O�'�]t4�L����b���v�������}��{}��� ���1�׺R����AaT�D�猥L�<2_Q0�Cz=ѣ��R�]���F(�א��1m.��|Y�l���y�5*a1�q&�Ы����͌S0'�~���5��9��y����A�a�� �̆����l��͠K__-�ׂ}-�����n��K�X,ޞ��18�c�[�}��w�p $@ۿT��,V�(gr���@efx)u᫧�y¶�4��(�ҹ��:[ɅlZ�h�Cj�v5O�kT�+�1E���2���2�5�,I#� x�s٦/�D�C�
��85'm������o}��bV����gW��V�hgA�bE�*",�����F��f)G�+%�
9$q�'���L
��E�_��)���Eab�$��jaˡ�w1��޲~�G�\��Y�#�/�{o��#���M���?M>��Ӄx�)�RQ>���C��=Q�ٟ�>}�	p�]Bo���G�p�E���_C��tU��i��Υ�<�A�*`������n�z�|�m�I�bμ�2�e9����@0��? :f�sS�!ฬ��޺� ��Ԭ�:$'M��1�92��jЮ�8�!�)-��b����qR��<��tW�Yw�����{��U�B	V���A�����_�w�Zs �ݓ�)uBo4���́F>�<m���#m<�;;�{10ԯt-�����8�K�b���رcN8����{������F��i�������F�M�~w,7Ϛ:]lx�E��_�L\8D,�ϡ���]4@,E���FG�"�����=�3j�ds(A4?vt����F���y���XtDޟL�b�Ug(���9<�:���K�3$�^�t��Q���y0�8z3Q��*�,�Z(��x�Ir��~�t>sNa<1�H��-�3>}>u�q���v8�^lڸٴK���[���g=�
�st�f��� �|��l72;�����p�c_��<�{�x򩇱~�kȤ9�ٍP*-k���`%�Rym}^}�M���1O�։ ���.�g�~/���h	�FDjq��w`��7$�r�%`��b	�<�M��뮻�h�<i�ؽ�S��2��ڻ����cڴ�U5�<Ͻ�ر�9��y[�m����je��U�uZݨ���_��,�s�)�4<�R���%a�|n+��\cL2�9T
y<�裘9�/��<^}�e��2���4�g5�� �����d�Хm�_&�2��}�x��^]ۀ@(,�a21�����7���:��r��օQr���`�ɐ�ds|�3���򟊍*f)Vlb��d����gצ������eQ���/?���Nf��q}<V��R�߄������*RFC�A%�	F��ۍN����]9��Rq�q��z��M�/���+NT�$_�k� O���ԉ?w$�D\�TRpXҰY�p�K�q�6�8<pX����Q5{�E��XT]~Ѿaz1���2%�i���>\�&Ŋp�0[��VJ���;�ĕ�=�=#q�i3a�+٭�;9`��́�Q�[E�����pܨ�R��Y�~\* S̢(�'�.V`鑓W%Σd��,Lf�� ��F��Ʈ�!\r��.�� N:��|�aȏ���7��V�\n�<�0|�?�c���=��E��F�/�K�mNTY<8���p�c@',���f��q�>����MTW�����Í��CV�E�ޤ<W���
��M��#��y���!�*���wK`�͑ ��r	���k�$� �0,�i�K���;'3H�(6~c���Fw��aC��A�n��{լC�SkEw�̺ E���8̺U���j�#��3��R������V�R�� 6���������k�����sp.�r��Պ�N:	˖,��K-���g��GAO_/��Q�P��m�x{�&i �5��3�i�T�)F۾$FF�����fF��IX�l�u���IY�nP9;���Z�쓎.�==}��&:�S6}]�"��M�4K^|(f�!�u������K˔ir_,h'��t���&�'�ߔQ(�(6"I^L�u�ۉ�x]}�H�ch�����_/>^��b
+;��ta��}H%-x��wa������ǎ1�es�B�p�Yu�4)T����I�H����	'#V��r#l�"��d�Rx�G��5�,���Yc�T�}c#������y�=[0g��#��v�k����/�]���[���d�4��O}�D<��3�Scٚ��\Z��o��F.4ԇ0<�����vn�!,��eC��Css=��������ކ_~Ut���Jp��q5C�Z���N����T�M����m�p4�9碷�.����g��҅����8��Oc��E��B&�L�]�%��n֯_��6�Wɗ�T�ឮ�D�ھ�m<�Ru�+2����D�`�k��s��9�'S�ǒ���Zq����H�,%"NBPMFL�ɾ��$����NK���B|3�1�0��&�dMN����:��c�ʈ����A��99���W�|}���g�E��e+A��Ga��5o��7�/{���+N�Sl�K��!,"V<���z7��(Da)�`��P�j�]���h�����ë�M�%��w9��F�f�RwV��fj,ʂ2F���X����>�K9q�;���K�aC�z�9d)��4�revֹTG��/�d�@3[�ᳫ������b�rQ[�3rc��>LbmP�ȦA�D���k&�jоy0�����{�8r�B�~�'��$��Ɔ�p{�8����/�~��������>?\n��o6���bG�/�#���I�Vc����z@��=8��ӱ���X%�	���c9�SN��+��_�ʤ	�`,Ǎ7܌'�~J@����/���˗/��yP46�x.�]�ф)1�5DV���w윍�� ����1Żfvb"����V3������]ds��:�耥��W�5�t�%�A�8�e9�;����c|&�0sw��@��A���?aeY�� m�_L>th����M�v-S[��l�2l߹��-e%6�xA)�p ��b�X��K���*$�LZY�j�e��6mQa���>΄�ҕ�<�������Y+�}�t{=Xs�K�P��.K��92�j�F`�/:㓽�z2&�8t9�����͟�HJ�ez#��Q_;Y;Fl1oP�Ɇ���٫
���V���@}�O�[\���@>�@��-Sgb���@W?���E��@]C38��z����rHeh��F X�Jَ��=}#��0�I�	���P�����,ƞv`��S�e6oOg�0�C�����x�;�Vaמv�}L�9�W���G	�ۉy����Md��)-¤m�����w��yKf��߿￷���8���ظq#�l}�V����z������>��w5
Y��Wl�(^/�&���ܹsq�'�ͷ6�����ern�L��(\n+BA?,e�4}X+6�8扣�����I3;W9+�MA�WJ��͍2E`JCN����\���a�ܾ}+~d�����˕�J7������f�5��I��/)�r���ҙ�j�142*VLfL��/|�4�'�J�ei�D�Vv'kGz�#��:1�~u�2�G���Mk2�Ҿ~���y:��Nf�b�{M5 ��ŝ`�~G�̺��a 전�#���9�)�fv���}�#-�yxñ�m�MoxA��@9] J,��`�L���O=S�%�y�*�9d�I�<���x��װ��VOH���N'���ōY/ �0Ԣ�E_$�N��ƍաj�0\[ś��v��K���x:������G���H� m�p��f�/��-Y�� b��d(��	w��HC5��0a4l-Љ�2T)�%Qf�ܰd5Z̙Ս&��Pɗ��Yѷ���!�D�q:0��_=��۬X��߰��w%�~��K�e�k���t
�>�W@Ul8
K���;��@a��D� ���ÄP�146"�x{taۖ-R�#v�a����8������h��a��\/><��T*V|��ӱh�"���K��M=K�P�X\E
j(Ҍ��Z+�cKo|�L�~fΚ(�Տ�Y2��#��t�v��k)�U����d�^�K��	3V>G3j��$�J�E��5�:
p��Q���5>،�?�f��� a�e>?
�]�`#9&AX����a@����N5\�|����4����w�_��Ԅ�%��s����>�eV�֩2��̏ي=���&�0�4aG>��r$�`{{�8��<+<n��x��� B��$,�lc������%?��>/zm�ɲ"�=?�8�3�ʰYfb܎�D�&usiJ��`YL����4q%ńY!,�'�G_� �P�w�QL�.���ϯ{��?:������sy��o�5�f*�EӘ�2�=���O�K�M�'z�M�ڌ�H{��ġ+#��e���]���j����b��|�
Q］AX�t��-�w����g��%���Y�r1��7��ߞ}�w �.]�ݻ���.�tzoi��T���<=�)w���]�r�)���2f�ضm.��b��%Ѽ��E��q{,6�pPMH`�c���;����~2S���W}r��0�v7J��*[asx�(���^x+��7w.:�c�;�"%����CV��n���3i�����_����������3G��Y>�N5�ɑ^/f��eK?קt���.�LI���I����f�q�D��sb��Uf�J�4���80��4�1'�����M3�"����:���ֱ�\�ʁ��H����f \&�<q6�����Dg�{����z����cɄ]��[���ٵ�݁Ŋ�TAd�:�%�<��G���*G�r��H�bkG~y�m�X���)L�L	�(�<�E7�	����B��"�DL����r:�k�d(�v��(�H'3��Fa-�d�bC�ZF��JQf��,6��9��Z#v����`��@}�LB@X��MkY���0�l�/ᰨ:��$O��
	���H��0���|u^f�ա�*�S�Y�cW/;���0�_}/mz�6��N`G��G.����m�8
��dE��k��b����5�_�\::d3d�`G&�J�*$���G��W��Q�o~�;<�����9w�
CC�G"��|��r���r!�PY���&�,(&�'3����w������JW��,m�F7,7ڇH3a" 6�3��7g_��]��ٚz�����7Z`���,��u¯`dz�:)��Z�0�3��(� L5�g3����e>)�@��K�\K2�6+>سG��t8���M��G4EӴ�2����[�n��ب<� 67=�\jx�͎"AX��iSZ�6^�����aIb$��ϸ���8���fPWW+�o_�)%>9��&�\(��ze�Z��k�T�1���"f�7�����r]�:*�W����"���,��F��ڒnfSW����*r����(���]ntu� AC�/svq�w�K��;�Õ����ll�(���`��yr�E��u#� e�6B�:t���O~~�x_q=RVW[�֩������c�f���Ѷo��s�oE��<���i���硾�6����s��կ��T*/��g�~B: 	dO8�8��X�l���j��b�&�jnn�������8>4<���;�^��E���X�~#�;�|�ܳL�����}(�����^3m�K���N���6in������B�D�oR9&�vI��	a��kHаt�b��+gP,В�@̇�/>�l����aY�k~�>���0��16�0np�h&L1h4��?�}Kv\�i>�1�8���;]�)���w�*g����Q�c��k����r$��a �̈�9v��F�Ƅ��3�\�f?j�_�er'�0s��;P�!#��I�9�����Y�,�����ч�����+�}�
e;J鲀0�}Kf�)���-�]��$�l�-����Ï��ņ��S�D�<�j<�pܢM�¢9�o$.�
F�)�U�C.:��zK'd��DS%o��g�j�R9�uY�g	�����%E�CN�H��
\^���9�	x�"�N
�z\ldR�XQ�P�K0��7ˑ�0�NX�+%x9�(�G���X��=�[mh�U��|B>�2�<^{�M������Q�ර`-Y�v�������j)�-ې������|�ż�$;ƀ���1������D��B^L:	®��o�ؓOH9�7[KK+�n�%���@P<z�`���g��5�-��5�?ڦ� &b��7�.I���z�����`*�-����S]z"�6hx^/u��<��k�`�&��zLɄNB�;ա��_��lC6@3aZ'���@O&�����Y��3��L���9)}��/�.�"\�ؿ8�n�-I^��¨�D���%�1~gٞ�r�Q�X1n~%6��1��E�U�?o�q����Ym�KR5&�<��.�P�YEzNM�ڊv���2q(L����`,�'S�C
�ݲ��鍍^c�;�g�V���5uD[e��d3x��:���Gz�Ӭ?�a��W{r��1�HUՕG�� o��Z��Ջt2�j��� n��x������[�?�����d-y���G�d�P<���W���;�X��K��]��I��e3)aP��6"��a�t��^�1�Y-��?�+�_�g��n˃��:�w�� N8��q��X��&$�Y|�SQU����(�߼	��{14�/����.N>�d<������V��/���A �J�x�eS���>�[n�CC�i���ƓO>)��l
"�[>G*�ix=a�-����������X���V}�lK�.F0���#~�����aK6d88��&�pM-F�b���q�Ēej�tvu`$֋T:[�����w�|4�Ԧxo�x�ǤL�u�狺�wFLq|����jΑ�6T�)���?CuM�Gd_bY�q�1�/}u���R�y�l��M$�4˦A��(��������T��g��s4� Mʜ�x�A7U`2�����*�����LWc�&'��l6h\���x��a���^=��7޻.g��-��(�(����.u��SW	�.�����^U���1�����s�S-Τc� ��7:甸P�O,���cttXuy�RE{�Y��K+Ƽ+�d��C4���-E�-�
�ec! q[l�Ė����z3>���W��dȼA?�>'�R	a��,N���|!�6s�qN�2�d��r#�.� Kh�����!���, 9<&3��$j�8�%D|>r	�Is�����X�N$��lq�ku��Q�
'��li/Z�.Yগ[��H(���rX]j��'�����A��Q(es�f�l��._��L��0�d�PD�mAf�Cp���w�����&�`�`�1ˆ�9r��|��~/���6*+U�����tW��%eVg��\��da���<��A�Q0��=��p�i�� �:�h��f}����\��t�S�wAʤ��|
	Ĳ���0��0�Bf��QrYa�8�X�����na����^^@�f��e��V�Hi}jC�h%v�8��݀��Sf��1�u�&�!��q��*"%5�;��5�, ���Ki�|L���    IDAT��<�ր?�/K�[�lQ�� ���Z� �eb9��z��VќN�V��0l������r0|YbF�T ;غ{�����o-�8n���xꩧ����~�r5'��9��f�ᦼ{�>T,.T�Q,X��"�,�[�^�x2+k��O#
`���cg�߅O~��}�����؏-[6#E0\�������a�{���ƹ瞋��w���k_��VQ�;�M�I��w�� �?�'�9N�1���&�І�&�sc�1�z�gq��7�P?��=Ř������X��ɸ8Г�9��/�����-���㶋y�N�,b�(^{��@���SØ�`���8������w�dq�����lu��Î��y��cO"�ȢT���3�A*ǚ��CMm3Z[q�m��Ef;1�ݎ�o��;�C4aLD�ό�>3��$�	�|b^,�u��'�
YC�O�ml�?)G�����ۙg�)�0t���U�m��)��Tv�zz�ĬH���5��� �\��06Y��c�8����'���	��h����5�\N҄Mm���CFM��O���U����ǽ���k�V��bņb�74��*MXi?�r�*L��ew$�(f3���(۽�������E�;�M���3R�0����W�R4�W�nC3C=�����QP�M����Aއ�N�%A��brX�CVL���ԣ��_S���(6@�[�����"v[y�0����
�Ơaa\cUr��ġ�����PS�ζH�S��dKR��ǒ���D6Ŕ�:��Y���:�H�(�P�����j�oB]U/��eB58e�	ػe;��g	����'�(�2��8h�b]�h=��.7`:�Ϟ;Gu�+R�"���.	 ġ@S�O���(����ƈ�i���+͖����j�,����$���on�}́a�!3ʑ��L[�c	�4��K[)���t�Pj~�Ձޜ5XS��C{9�A�r�A����L�a:KT�hXSe����j}Oh���YZ��? a|=[�)h��L�Q[_'�J�/Kv�n�[�Q
ahp］I>�O�a.�Otd{R��E��ͭ�|L�\##��c�� � �N�,����L�c�%#4X��#�[i֪6�!�	�9f�#��T\{���z��KpF&������a$����:��3���G�0��d��S��`���/�@��]�Ȧ�*�V���3��o�{4������567ap@��ė��c�<Ѕ`��l.g@���"�������i����Tc���BKk=F���`�\lݲ	��^�iC��%D͛7_�u���71{�<iؽ�c�,Vv�t�N�ъё�޳�}�k�pڬHg�"$W�d^�����`��U��n��f466�y�]2aW^y��ξ� ��_#c�ز�]̟;���X�p>ֿ�":�w��ct��T\4�Y�n��4YfB�-��A�PNO�nى�x�TV:O{�q�mw���o�c�=%��V�8?�������b�Ƶ���/�߾�5�u���*���'���²�~�C�c�"c�ħRuCr�k�"�0��ye��߫8a����֭C�XFm}�Heƫ?v���Ξ3�RN���L�7��EFA-�̟�3�a��$Y�p^�/F��aZįU�f���c�@��A��x�$I$.��c�#�D�iT&�� ��1|�s�^0�$iv�6��ݑw~�4a]]]����z���6��Vΐ	K��~,��7�������p�����a���A	.���?�����]�#�EP[6�7 z��#�G�9l�d��"2W"ڟ���fKfG�e��C!�Ȓ:�SD�bAY�y;�U����$�D�|
�6�M��j�n(;�~/jZ0�0��#f�d�Ȅ�Ό�6;(��gp{�)���Ν�t")��v�ltY�b~Ktbh�X,=2����.��H ��-3Ze����(����J�i�'�8��,G����7n�민��}�l{��-���7/nx�\�����Ɏ�������ߟ���#�����
W���Iu�u�J�1g�0^+�a4�x���W2ï������0-��b����H�R�8���v4McP T;RO�g�0
^[NL�{t�t7�*�M4�ҝ���Z:�e��]%�=��Cf��
�,��2F}���f��mR�����n�9f�-��Q��t�����M��E��G�R��=�M���M����,`��YԆE�:O�:���,$� M�#�����5"��j�!b�AU�����77n���}cѸ}�p・�s�;>� K5(O>����i�e^?Γ$���!3{n*ZGH+
�,�g�
j���U ��F�Q1G�[U�_�c�PAo_?��J�(��2~t�`��]x��-���~)`�%=Z�#��z�b-���с�&�N�Iklh��h
���
�T��BF�VM�u��cx������R�{��'$�aR���OG:�ŏ���7J)��m;�/�#0"@��s���}D�CX0g:��`���\L �����-l��E�Z5n��x≧��Hrd҅^����Ghk? ���7o�*��ؿ���2��'�����v�!������%K9����q�W��^72`�����K�w�	���݅s�clv/>�����DU��c��p���_z�{.���K�ٰ�������L�d���bӿq����a^,r������5��JB��$�M�6I���Q��\���K_���6+��8�e�������+?�F�@֬.Cj��&֭�=�'tf:n�K�&�3�t��Q����s�C��UMt(�ur9��i�{���q���\.�;���v��;�wo�u����̺��=�Eve���P��bAXf/.��Ta�rn�6��Kf��������y��>�k��0;��>z�p��r;���E\o�`�Z)`&��@�d9����M��$��OǱЩ�L���%BvyY�	�/�h��ٙ�Z�p���l���G��PC5F1a6���҇qX+�k�������g��C�gϜ��X\�����Q��S��]�"��ʠ���!�ٳG~V:�[�6TM�B�f�I�R��}�eKh�V�ģ��I+>�b9�l:��o�ǻon��.�m;w!���N�)>�aQ_�G{�9�t��/7,-(v�����D�t�̚�)-�8��C���G=���A��lt��MY�0��r��v�<�w �O��U�F���� R�o�VA�V:�jFUgx�V�ӫ��1F7$�`#0����gbh��@՚�۾j�����h6>��́�wtC���	��e�����hG��E%�w2�w9���ŀ���N�A~�s��ǂ��'W54<,A�k� ���5m��O��?��i.G�sqޠf�~�ۥ��q2ʦ�Z +�WƆ'F���Y���j&�m\����5��yʹ[���N�}��a�ǇX��b㛖�.���)к� �/�^�tx'�#���H'a�Ѱ��b��L��Ӊ��.dq�=����\"���>�SX�h\N����0�
��6GF��8E��Ⱥ��8���z�i��-EKt�'W���g��֭}_���l���U�5RU+Z'��#�1ع�C�6h�AV]���9�;v�&B�H	G���	ry����2��ߕٍ/<�*�~�Yi�PF�^�x�'q��.G_�$y
/���LI�5kvm߁��f�>�0��`����"!l�(�*�*4��"��Y�/���t����V�No5��!����se�U8�̳�̳/�pc�i��&����3O#���O�݋t<��\�Klߺ=�]"� 1�u@ �A����G�}��,T��>dff�,LZC}� Y���sS�l$\{�}Z�6I�
�̈́ac��1�C%��;��V���ɦf�%6^gI�A�~���hm�����ԩ����k}�iT��2�xRnj���!��&� �����~_ t����b��Í���/�)c�^�T�<���<��&���*6Tr�9�(�K������/��+I8�c8�@>+��?A��.����_*vS�=[[�):�>6j8�t~�R�����3e����Œc�a����,C�W�C��e ͱFԻ[���L�\�f�h���/� �����_M����t\uJV�l0ї��2�7�0f٢/�vy7F��K�������Y \%�ks#1EtdTn�`  硶�
�������N�m��1R�B4�f_-.<�K�Q�,�h�F���;�������.�pg79G͢��$���`	#I��E���,���W^�}�>�-۷��e��vN��I�9k�t[���k��{�U)+��$��&��P��M����m�� �|��L̊TԻ����;�gy��W)j�d��oh�j&��0�:X�jތUg��O�5�?a�h)�E����㥱�_|ބ[�D�����h\�'����h�J)ro{��y2a|>A����܅s�e?�c��G����J�iR��#���10��Cvs�����jٴB��<��'>���.�%�=Y2/e ��9����ɀh�;%�p긆9�/#��ev����۷o7���gIR�&��'PP%H5k��&��fQ���9S�Y��R�2��e�Nr�<���mV�i? �� ʩQ��?�+����H��<U�)�6��j����J��n@ ��I~V~�p$�M／_����x��9���n����^wֿ����K1k�Y�&h��]�����j�5
��A���j�sOF�c�����Nl��>Z��U:4ꮮ����G_�0vl�-�0����?���2���ڌ��.I(y=i�}�6,_�g�y:�A�߳C�QW�Ӗ6�Vɳ;d��d|f�\���K�����4L�C>�[��#q�Ϯ8�p�[�&V�<�t[6��Ay�̪C������S�=�g�z	�����r���vD��r�Hw��[Yfˬc53rt���ϭ1�&�d�X\�W�Oˎc�[�����%�s�>K4a�N�M�v62�iӲ՜f��ۺQH�$�P�2�dvK���xd��q�-�����������df�4X��x��:}�fL��ɱN'��׌L���j�s��-�e��"���o�Oa�J���?�y��O�t�#Ҹ�ĒR��r�T|/��ه�/>������a���C�P��@�X��s��N��3�@��Ef\�ҡE�T�%�eH�B������mTݫ@i8��sJ2d��.n����L��E�C��H�}�Z\�<�Ti�^m�*�P�P�	#��!�T��TL@\�%�b�J=�!��l��� L9G�1]ݽ��g�)��b	�b��n�/r�ѽ����[����� D;�p@@`�`�P��t�lU�<9��4bɬ����bth�d�r���71��-#h���O�����I��'�y(&�Y/�'/��wѶ���d�rf0�Ll�'��9�K�d��N;��H���a �|c~��u ��m�J��������byE�+0@&L�M L�]BPHͫ�Y���.O�uz�	�R���(�g�q����Ʀ;��y�_��r��!��L�>���UGF��L� 6c�1CY�|	�Κ���v⢋.�}��+���o������͊T&+��n��[��H�woB���c�0��@kv�V��Wt�,CRH��8n�,��}^V\c|P�C�U]UcL*`Gj	˖/m��ݻ��yo��p)o*P�͞��12�|�>xMX�ך>}��|5r¬U�[����� Ly�H6�%�ي:׉|Vtu�:{D�p[����)P�#S� �+���.�O<�/<�g�U�aU�hlhAWO�$=}���G�1�}c=���:I��N�����p�-7"��������0Z[[P]Qe�lA���%ص��Cc�d2%�w�"��q�z~�^���s��W^xooz%��Q�Z�?K�3��F:�٘����)Z?�OZ�\vٿ��U+�c�,Y�>�����f��%�]�_>�,�qtv|���6�V�d
�0+S睱��_�<3�
F�,X~*����Ӹ���op-S����� E&��<H%X�tK_�j.�؃���ګ�[o�	�����������Z�9�W�"u��87ӥ�%�6�2^J�I��؀����rm�ɉ�[|p� 5a�S��f�\�Y���0���
�Q�Lm�֞��蘢��G��`��F韏c�.mjL��J�(��o��?'��'��{�O�W�n8��b���},ZF��L�H �wy=�9�ޛ,���Ox�S@?�U�u��p���uˑef��(��N,��'�?��L�T���p[J�����_t;��m?<5S�**Gz�C_���&���Fn���B���yT��Z�鈪�ޠ�5�A�Tٜ��I;w�� ���M�'gE�Yg!/���_�*&�}����A]�=A�Z�AX�iV�0.@o�S�0a\Xd�da�UɃKD�@����:��(��0�݇��.ģ1Ѹ�>a��~]WQ n`@�Q>�Gۮ���ҘR��
�ߍ%�Ȑ�\*��ǋy3�⧗_���>�\n�#h�Z jo�ϟ/bc�)�-�[������6z��h��Ī�ܬ�	#p�f-����I���>ځ�L���'-�����Jώ�Ե�"&��ƈ!n�b�í��A�)m�;�%�̘g��D�A���k?9-F�;Ә"�2	�
�
���H��*٘�-�s�@�Nì�M'�x@F|6Mx�c&a^�9�x��Y���p�=���/�L�.ت*�\��8�3�66Kǯ%Gf�К�k�1r�������؀�d��9��ߋ�0R�-hjl0�䀿�y%#{"e�	��4
�Ff���u�u���Ϗ��[Z�+�E�E�G��ן��ߖ122ވ�o�2@���&�dLoԘ*�`~v��T(�͏�1�E�mp}�ư}�f�4 �8�}�X�|1�>�ۆ'�|S�f �.� �h�s1��ԡX��M�\^J�<�D:%�=���m�.-��o��ױt�B�؋7ֽ&��~ޯVU�%��hTٕ �n�n�����=>@XE
��Ξ��>
�{�I�����_¼ys���O�_�ut�߳�CtGGH&��,�Z}�[��W����qtuw�s�M7�g`|Y}��ػg/X��]�,;͓�����
���e�9���_�J��d+�+!�)c鑟D<e������{#cjL��Lj�����y�<�6�	�B��<�}�R\����٧&1���X2���6ʐ�;2�L���}4�:"�R�Py�V*����2������g�}���3	���1�M���c��,-�dV�az��:�C�3j4c��7��R�&"��Sω��U�Nd���l2�4�vKW.���c�tR+�#.�kNv���?��$�r�9��8����{o�X���>�i��k^��i^�/[QɧQ���l���9^xR���g���C�������4�zd��	��p�l�!WR�Z_l�� L�ᚄf ���rS�����,w���G@:���&3Y����mޅ-)��M���*��8��[DMAo�r����yű�c��4`4Mˑ�TL�6�A�KG&L@�[����1�J$����!!	BNJci��!=�������:m�C	�s*�W뾞>��� �Zߌ|"G�{�*�w*����Y3��\Z�i�Z��e�қo��ؙ����54c�<����_����t��
<�,ղC��Z����l3�SL��	81��r�������?a���!�Kw��n���K5~М��#�V�`:(j�%Cx�ńy��:�٠tI��n���	]߃�������M{���"����� �lY��?�A��`�&&D��A�zS�0� ,����B�*"@F��C!|�3����#��/��2����
�Dp�$q`4:&]�d�fN����>Dh�a���4f(�S�RP�I�k��n�Ɠ46�#�{�X�c��E@�I+@J
�=>�i/!�Ԡ��Nm�Ip
�Z���'��0�If_a�*�    IDAT��׋Xa�U�K�]��������:ka�|B�����D�^ضH���	n�H�����c1$3	�DpVr9K����Q�D�O�U�b=14���w�Rq#D�S��ˇ5bv���x�USS-&�ܨ����� L��[�{�MG�L��<ҕ�,�JT\�2~���uع�
�CU�~N��:a5����'���p���`����Y�{�.�{����%�B۾N<����"�<�+�"�jn��&̜9�Tm�q͵�W1-���!��,]!@(:2�dl}]{�v�w�Α*95��q������?�D*��h���G����4�y�M�x����0k�L��bs㤓>�{��3�������I,\1�]����㇗]�����.��rd�C��넇מI�W&��2B���ސ��Y��%U��:���W�Iza����;����W	��x��j6�|��a$�a-5����v`Oi���U�ks�0'��ߛA�9�h�K�!s���L<��G�k�y&=��Z
b~.�K37�	����@�N��,�F�>�]N�窏'[��{�fK�qe�dE9G7�1�փ��p�]x&j�xY���RL�_X����]enPe��)�ˋ#-��6~}%�2�3�LC 6@ɿHe�M�
��YA��-n7|������{?�{i:SD���(��|vG��l����(a��8;r8>zPwd���d5���8�[�M�%(K9�R("5<"��`i��ƠӃ�P�����bw��u
B��B�Ǣ�(
(f�H�f1�=��X>��S��ؠ2|N7�jho�G>G)�Ă�3��CCh��A������&�s��ϭ����3�L�t����ž�va�X���b$:&�/ļyDKDp��[�2��"��"�����QJF9��#�Y0ޘ���8r�7ngg��q������9	�Ę�c�u��j�3��[`)��ܸ٧f:X�!Z�Q�����G)��(\���<n����:^:�Aq23�%�ɜ�	���*d2�;2��R$���<���\��}�3X�p�t>���xw�f�L�a�C����TAU(��3f`���ۍF�� �L�����S^I9��@�|��%E2i0��<�sHwd�(�/7'r�+�lȿ�9�ڷJʘ��0��6�JƌCS=��)��u����:��k�P�)g��8�V���2�Qe#Q�,�*2p�tR�?'V�1D�b��MEQ�!� ��!���|m��׀��1EytD T�\�L��D�`������ǁ�dM�"Ǹ��h�l�ذa=j�Cx](�"��<M��),����.[�/��
������B�Ĺ�^Ccd�O~�8��%�����{�6|��p��w��u
�9�)�����ǟ��/��a���sϽ�Y�f��n_/	�#g͚���W 2A�qǭ��ob�̹8j��H`���=�PW�Fھ�Q��2G�!fDm�/5a�%��G��XΎ'��:n��n��v��ɓq衇a͚5h۷�h�4ˑ^��%�̨C"9�K��5|��/�����[o�A@X(D�<5
K���A��cr��XiI�T��˽�t2�P�54WenՍ�&$�Ճ�Eh��E���1s�?����ThU��1�]zT��9��5�a	��Md���Z�J�$�6�x�~�]�ړ�ϟ�E��9�i�4�SRW$Ȋ���a�>^�O�]�ПS�G6����?� ��Y��O�~K�]�2[�����j�p�!,��'��}�LT��������@��<8���s�$��ʌUke(Eo8��>B#e�=��#�,MJ����e!�D�25�6+�*��r�?�(=�ʤ���zB��M`_<���1�H�'��B�eD�s�R.�A%�g�H�8��qvd���s��H������L����wJK�c6���$�@䅹��`ϕ0�ً���èi�G�V�"!d2)U����s��c��� �p[��1X{��9=b����_���~tuc�s?�n7.��|tv���ys�o�C�����6C���("�OJ7�* ����]���.)��.#�`���WE��7 Z;�A�S4m7488HSe���� �L�f+x�y\dFv��.A��A�������N��+1�]�, �ZZ��gᆮ����|�M
�y���%��&A!� 7|��=߇ݑ<N]���dRe��r��lvrw�d���Lm쎤S��#�|"��M�s8p�Eː�˖cÆ�8��O�Aݔ)��,�,���9��d���,��fs�	Xэ
 �-_M]_bYb�����E3Ա�Mu>�lhjjQ�;�`dOx���gdeɰ����x�$�@O6eJ�\7��EF�N��`�������[���L�����c��d3��R	�R%��Ӧދf�Y�3���Ȅ�@��TT�Sj�H�Fac\��Iv#�4Max�6~8�~d�x�A�����Q.іr/��}��+X!E��6��T� �}Y�<O>/�]T$Y�6u���1��翊66�0M���v�q����'���x��5Xuءr��޲̴r�Jtwu�`sf�G<��ٍ,K�����bѢyr���1�6����>u���� ���0�=�HT
y��J�u[�N�n+�/W��(ǹ�6)�ĊX�b5��F<����Ϗ����W�m AY���1X-.T�8\V����:�	_��8|�!x���q�UW�($����<�k��5�1�bP2CW{�G\Ϭ�Ý���������3���[�|9��bhk۫: ��4@�Ӄ�O?] �t� LO �gP �)l�صPO��a����m�l����CM��JF���{�^�����x�|A�".��D\�r/�$SR�)�e�ۚhTCȯ"��&(6���X��4J/��jj�աHz���o|�q�{Ƒ��!��y����k�ɪR����.������?��Oӄ�����Z|-+
+r�Q��i�؇j�.:���v"3Љj��t+�N��/uv�h�����!�ר�����*�L����8�\"cBh��.1�)F�Zg-%0C�(����Aj�
�j���-]���}(�y=Ɓ�t4�O.>]A��v�Y�;��a�����>a,K���hvx����Y�\pR�.�A�;|��l`��͍T���4�T��أQt�E�U)P��a��Ձz�Syil�������5��=�p��?G>�����y'����#�7�a��9bM���T�@W�2�X8����Ó�bQ1d���?Ⱨ�Ď];1m�L	2�.ļ9�1m�t�_����={�m-���y��b9�hi��{ܻF�f��EÇ���m� o-��W�g�N�4���.S��0��f����2��z#�*�_�s�M�Zs9�����r:�����5� ��X�����(s��D������d��N������>cr���dVQ[8�����u�	1�jٕv�o�.E>�������7_$gȏ��)ZG�;ѩ����|A�x��a�u�k��8�Hg�<�`������1c\n'�ly�(?(o%q�=��pTYX^�Y����5�yb1� M]�`�	���P�^mbи��<.�������ߋ��!��5T%h�l�@�j�`*�N<��%��/��ٴk7�G�ʏ�*/J��L.˜�PDuM�H$|��Jp�ع����U��V�(�x�j�<�`<nz�U�bdJ�/~�}�B����فb!�l:�T͙�~�e���fpp�\�?�0���h���SjS�.��"N��j\���_��}g��Ni�:�Ӎ�o�=��SO����Ck��P#cI��6������E_��� 뇋ɫ��1)C�Յ��E�N��1���F�����P��U�<��c����e��h#��:����r7��*�f�����p�i���I��؈��)j����կ��C]�%�ȵ���kq���{��%{;�{�4��ż�7&��.lN��/���ب�Kv<�L�J	���:��d����O�<�Ē|^��
#��-&�F�7c�rδe��f2�Ҩ�0��9�wx^��##"9�5A��JN'�kj�y���M�����a�9���m���g�01��x0��/w�Y�����������Q�?�\^l�H0p���e�h�2gjK�$��A=}�p9\�TWaldTz��	U����l�p�[�idp{=��i3�=g�?� 슿�q����|k�ۼ4/���c��b�7-oq�Y�':��^lE$ǆ`�זף\�9G�ėDU� #��d�f0� �E %��̏�\�sF	����(������2�L<����m�b_x�k �C(h���y-��\��e���8�,U�yn����
��s[��)~ޤ�������ő��T��Cf�(I�LILZ�+|e?�u$�B:�)��a�YHXKHes�?00��h�L�Ձ��R��i�t�6V-X�}�d���\u|6'Z���ֆ�����1�9��ї(/z._�C�sę�ã#r�����x��װs��Z�x�hs8��:��Us�Q� 3|��5�ͨu[;�A3�b6ο*c��]��I�D�lݞ����(=�Y�2�Yk�7Xa�
����e3�7=��#?��̈́i!7AϗD����|_U�,��8��N�q�w�E��.�kЩ�CͰ���)�C_g貴&L9�^��s?b�\^��Zh=¬���ǯ~�+Dc�b�ʌ����?ގko��r��:T聗S>S,%Ξ2�RN2��c��������i���VV���*	��K���iǶm[���F�H�0��U�D�2���uu5�)���M�睬�h��~�	�ɹՌ��^�w���5��i�#�6A׌ү18ȫ�9�-���y[��$e,\�\̜_X���0�^��r��rZ��&��
�N/rE���Q)�a�xņ�nq�Hz�(Y
9��;el�_��x���R���m��ޮN񻪮ᨣ����\s�5�y9��I��{	/�}�W���^՘���U+1��
�^�U�v�ux�٧p��7��o��e�p�y����_Ă����O�'���_��X
^_X���s���G����f��,�)�TȠ����}H�ȥ��b�>�m6�TQ,������1�^d��X�B����Vtt����X<�?$6:�:�+V,öm�PSW�c�>^4UUU!p����Q�R�M7\�5��x��RP^U��}cv0u�ҽ���²e�Dx���9sg���K�.���V�d��tRʀL*��5�Ub���Z*��]$�H�J��T�9�R�}Ƶ��͝=W*�fz������_x�y=�.��1J7�0����s&.�u�|.(�#�/�\r���cU���Q@��	Yk&A|������_RMm�L[*��%ag,P3(����&11�BV�9 ������\�l��=��~�����Oc�~��G?��������BN{�� "�<f4{�L/Ϭ�e��2�8l���Q�gd!SS�L�\T:�&�����u���NM0t�W�)R�+$K�"�w����e�,��+�p$�\�����]F[x�{P@A�i��W�t��a6�{��#T�#�&���	�d�,E���f�jmnm��C.��;w��?�V���Kʊm�l�m4��ˍ��M�nm@�����d��u ����F��C}M-"�*�~7oz�x
�� �͚�ۯ����t�͵k��'q�1��{�|���`�F:���^nn1>�����{�(ɪ2[|ߘ���y�ʬy�b.e�[[��}���q�v�6�FA�D}j;<�F@���������ʚ+�1"2c�{c���w�Ɍ�W������U+�Ȉ7�=�;��o����چ�~~��Fbf�]8��%�	��wX�eC�A �\Q���](
�Oq�Yd�4�РD���5�~%��M���#A��K��'0��CkȖ�5�ȽЬ���^Y��:^Q����8�ݪT��J���5����?�^���k�Sa6�"i=���n|�Ϭg����&[s L��g��%=�y<|)V|<� �����dIM'0ĠY�`QO/v�܅�mn��!��ҚK�tV���U�J+��L��_�Aܾ�L��~�hƉ��i4�T*!�s�X������y��Uk"�6>6e�|���o*�Zd�#ã�qqḤ��8ǒ�^�g��g�����:����\8������G�|�X��"�j���V1�����J�%{�A�0�x��5�����-iK{�d�>4�v�����u{C
�9����������U)���hnj���+�o@)�C��#Ȧg0����cT.�l�MS��/�o~�(���]���-�1����된���m�{�z�{��x�7J%$��t&���V���/��b�L� ~$SY�]s:�����+�7�Aa�Z�uG� �2����fQ
�
�"?R�	��1��gӸ������g�:��E
�* �W���x7֞�k�o��F��It�'N����ĸ0��\��!�!��(UL8��u���G�H6|�d�8B�	{���"V���,��5kd74F�a�za�؀�㷧�G�"�EnPs(�0Z0��Ky'b�����%��s9����c�oZ�p3�k��8^5��c��ս*�T���j>U8���:��w���U�=��%�Z�l��eft�^�$��xԈi�9�����$�d�T�!�2S�Q����;uݪ=Seɲ����7���YT|�gO^���^��h[��u�QD՚B�_ª�q��Ch�԰q�R,�nƒ��p;���i9�vJy�6��z���L���5�zVƐ�g0yHz��h�h�ʼwM4\�Z��(��ȥ'��ٕN'��
�0�|�q�``�Ȕ�0rornLnJ�� ,��~lj&��I2a�����1y�̩�ܰX��LI�nl����n&SIA�4�%�88���p���T��{if��T*�&3��>��iol=5r�\v�Gq:�oK;�3�$^{�e���Z�q���Ǳ}}��lmk��öI2A�NY�;�TR�66�%K���6㦯~EL>.���4mj��= gK{� �`th�Ph6M�A��f����c���R/�:T�	<�,?�x���f�89���=mЪAU��KMɄ)!�W}���]���N�U�d�r�؋ E�v/J����k���лJ�'Q��,[���j�WF瀫K���(�
�Y�l���q�{Ⱥ���#�026��% �����lF��X<&�`��o����A��FcW;��\$:����]%��g���t�|&�@�mYp�ƅ��8�;g.Z�nmk�Ν;���'�;�/ٰ��qIE�!g�;S��Bn�J�m�tړ�q� ���;��+d�t�����k_9��~�I��r\�Ō��\Zu�����.�~oP4�cS	D�Q�<�K��b.�ޮ����-g��|����x��gѳx%j���xm�^ٴ�r�j�E�� �1���t�$���fi�����ރ�I<�ģR���IE#��n��z�Z�M͍p������l�Qsz0�Ja��5�
��/\��υ��[7o����/��?��8v��j	�o"��) ��7���bP��_��}�X弜+�@�H���9Ew�Mj��R1�t����O�S<�����)�B���z;[e��>x�_���cM�������+�K&��t���qd3JSy{4��C	���mx�G��e�!jZe���^fij�g��MC� ���a�d�-[*��m�>Z�����舀.v���nj���Ĕ�K��Hc����'A�?献�`��iL�-��*�,�z�S�?������t�y��v|^oNԦ\	�E�
��4�}t��k�N�ylW��\��]��8��1UW�0e�~���<W^�H$���Z;�"��M��&�~_9o�����ο5C��Mx�)LX�Vs��Ϟ����_��䎯ʲj̜����I�}��2��y�����z�B=3�+��43�Z�!�>�c���K���6B��^���\]]Q    IDATbC�ži�ǋ���:�U�1*������ ��|6J-�dт"��3��q��p������,� e:R2+v:��w>?�5/�����8��	�XW�i
5
�Đ�T"৷� >pVD]A~e7�D��8��Q,]�)����H�%118W (@���U�?�tj�G�QH� Ps"��"�	�*�%�p����n@!�������[��JH�:��n"c�rx�σ�7o�7�u��"�~��k�2�p��}΁���ꙹ�, \<�����@7B�	eW�͟7�iK�T��K���+Ɲ�Wk_,�>���Ս_�U��5�C��&���`��ǅ�;I�W�!)��I48T�e���AT/��4W=�����\���4��x�B-n�y�-j9�G�p��{GU��n�JUȓM�w�J%�l����cC�,a��g���FDkE�yO[7��*���z*M��$�i����|h�g�f���}^P7�$��<��fS�����S
XQn@Q3ӑ�/z��m�x�x)��`��E��^�n�n6��R5#�7w|i�!�	�� ��a|j\,u|A�(PL�q��DZD����$���".xa���m���f������`Ǯ���w�gQ2�a`�	��+]((��w�قg ,N4j��,_�w�yF����Q<���ذ~��m~���Va��hl����>�U��6o{.oP�<�z�q�7�.�v�<�8n���L ��O�t~�a�v0+���D$��Ȥ���]����(�9��e|�P���;R��"Bf]�	�>@��Tf�X(���&~�㟠�^�	L�](��r�pb��5���D��#�dW+X���RM뒩f�Tȉ�t��9��Js�|�����*}u9gs�b;m`$TT��P���oVd�����]��&ӊ�H�17<�����gҜ��l,�D���&��,���8$8��8��� �c����0��n�6b�m�Y[�S�))l��i�}��x&3�<�w�sV��C4f�QU������\�~��t�>�:�c`�{0��T����D�W�~�/[�#G���R�����z�F�x�W^�I�*ߛ�x�@��?��_<��=���+3�"J�)Ă@&y�n\�|vNg���4�Ŭ��Tk�#��U�$�L�ҍ��*Cf�i7}���o�Ik!2Meq=wx��_@w�*��w^p&�X��#��߃R�D����5?n���7+{�0lq.A� �7 a,.�&���GGa��"c��=���l
�%���K-��8t��먑�e�i9u�qx�T3h�֫���.G��`|l�DCǇ�pyD,���7�Ы$IL��!�����D9���p�=MIs�]�����4�/�E9[@�*sy�S��B��ѣ2Q{/��َ#'��O?��6m���������,���Ěޥ��-8H��i����?���$ VdNf����&+U��3٩&ّ��4@ҋ����w�&'+�\+�ָ��0���N>M��]�>�fXd4��SZ\�������U�A��V��_O�<�Ne����e�̙t��B?�	� �#c�����js@��ě�������vV�REA~ӂN�.���q��x���M�U���U"�ć�ɠ÷7��`5�$.����XeG�kM�vm�+2����eB>�I+�q
�y��M��t\|}Z>Sy')�S_ǀ_�����tW�.P�/�����ŃsA����Zq���L��DbB
l��ݱ��+��[�8�����S����b��v¡ �'�x�9V�o����۞\�|¨���V�\�ˣ�}�����&��3������[���G�����K�:>���ؿ�O���\�f��kz&�H4��/����~���?��;w������������Cx��-����.��bi"�uc,&i�/<���v��{Pl hUA��7|���_��s��rc�F�4��	��T
��ѡ�Gg[�h�
�&��D����s�.���̴*���ʧ�!${n,�zz��_>����9�݋�#X�l�lK�<���{imRF ���d�?�2��|��w���E#j*���H>֮^�L��J���Tb���X�t���^rх����}� ��<�4��MU2ን�!+* �����^�����d�� �\��$3��Ci���P-�T���I-2gd��G���x��\��Km���)�G�E ��EO��Hp�3z�zr�Eƌ�� �b�)���$d#	�0�V34��t������w�>_�𛀿��&|r�Vs~��/���6�j[�"[,�Z�Fs̍��8��e�GQEpQ(�P�(D4�Kg��j�
����Sa�>!�&;`�N��;�u����%c���
����PEE\��w�ӗ�(%ᨙ�e�0,!��Kw~O@���0aa�pԁ0j��3a��/���Ըl�RŜj�D��y��N~/�E(̧���=.͢�EΪβa�G^ۋZ2��p��&a�bN�B9��ȱ!)k_�x�z�Q��Z�"U��|e)��^�\E�XBblB��LP�@g����l����ֺ;�p�-Eȴ�2i4�6��v`xr\�y~�Q���(���P0t��������=�[U;&á�G�TH�G�Բ��N= �)��td�p'c�a[.�\�5�uVZ�ϱ����9�����,uf@�ϋ(��V���N�����uѧh�p���:�)-"+��D?����9�ﯟ�O]&�Y!��;�`F������I�\F"9%� p*L6�ぞ_Q��Y0�EaL� �Si�#!T�.@��/A(B�������-*��j�����퇔�
��k��0�@�>Vq)����Cp�q��M��LNh�LeU �kCtd<�,�6��)��lǆ�!a/�'�C|�?��,H�0(�7K]���$������{�����	�:$�g�)�) ��6p��AlCV����g�ލW^~�<�2������e���Q5��8P*V�DU;62���x��cJ�B$րg�{	7��E��*"/�/Z�;�y+J�4���)1��3�,�ƌx+�J���֮Y��N?�>��z�%Rm�ʎ�d�G�������}�<��r�F��da������ؿ��I�.ѳu�/�����>��O�O|N�oLY���>DZ�wh �dF��ǆQ+[�}�f��\Q�^*J �oL�Q>�k��ҟ� �����H��4o.�GO�df��e�p�x�*��!�b��K�v	���q��碫�n���W���o���c���Y��Q8�z��4ӛ�<��n�U��s~[ظq#&�&�'7Kz	7�XʦB�8������������_ujJZqsL�h�{j&�u���&p����ƪ�<�r�"[#�T#�
��q�l���8gl�zͼivXO�ߞ���r���g7F|�Y���4S�������t��+e���P���7�ɶ,�h8��/[�{�a���x�j5��x��}�{i[�+��;,�7�19t��/@��@i$2c���EERE�L���T(Ѿ��h���M#�+��Vө4\n��LQt�}7��pr���'�`�<{0.�k5�2B�>��w�KQ͍!覠�&��w�Q�F��o���a��� ,�M�a�=�O�`���ʥ���L�4o�����Sr\8�� �
f�ܖ���v�c���H��V���B��#0'2�3��e��p�B��&���B�HM��Ɏ/��� ��I� ��K:izx�L��qD�Ƣ�^���tؿ_EN��Ǐ�kQ�b��%�EB812�pS�0~�XE�5�*N�j.&����6�
u5�:+�_V7BV0$Ȕ���e�-{�B;��T@�o���ɉ�EU���S�%�,&�JL����wiA�_��ږi�DR��Q�0��:(i�Ŝ�B�0�G�v����v��z`RϬՃ0����J�bul�uJVm�Q�Ie��RZ6��V���C�w�L�g�b�_�=Ѿ��m~�jE[+E�=͝�Au�P���.�,zL��z�R9
�2��~\Ȩc����� ��ܹsV�B��YO�����������������u<���� ,�Q��Y=�EKkyOy��p��#SJ�B��n�D�#���B�bn(X�hUU;2ѭ���s�����C��
������w7��N�;2�{��!^ٱ�KW�Ou^�pLD.L��2f�<�pu��3���]��-߂����;(�1�ǽwݎ���F�ȡ>ajhGp��!1	Mgs�76�ΝƆ&�XA��a`lL�
�ۚ%x^{!�[�{����ȝ]�^5�XTlP�6=�n��߂� |�Yg�ڿ� ���b̤E�ؽg7����x˹ê�Ef��܄L:����d ���".�^2/LK��+�T�q4ߴ��n�GĚ���008*���\A�������RZ5�ްg�}���?���=�Νw�{��.�v*�L��G[<^6K��.�u��thko�j˖M2�9&y������jQh�9�X±(��u�W���������}����,W�TT�����Fβ;�06��N�c%�'��iN-��Y]̢�Gx�x�L�&�5��jzVW���gq�h�����1�A+�IK>���t�Pl�!���s�Ź�����<����1<b�6ӕJŬ��h(��0��o��1a�k5���_��{<~W-ܾ�BϤ�$�Fd�~���$��$��
����&\]35Dl��8���'�*x������U��Ơb�&�R�w��fK"�Ρ	�n3����'>x%�8w���R������m7��+��[@؞���#�� &UI�P����	��"�o�nECG�0`�C=�����d�LVk��2!.�BjGTq���a�<U7B��^ٍJ*�x4_<��g��X&!��w��chin�����pl��H@��Q0ͅ����C�S��`�H�).;��B{Vafp+�,�o=WXŇzH�:?����ǿ�)�4��{�������?+Q��rJu'@��,��)��5�*q�^��B7Uh!7Rn�m�)6�H�kG��f�t�O�M�`Mj�y����S���&����g!��1$8���f���^�Ō�V��;2�t�лR��y0���|o=�Y8~F}jL�U%�,3�є���Te}������rufA�x�iZ�����>��:=�ړ	#�J��/�\:(طO�?���i��l�DU�+�<n�6u�K�J
P�j�T�å��|Ĳþ�j�l>��k�N�j�nţ�+�eJ '#@�K���^7�������+#�����y��b�?�n\�y��8&t���~ժUr�}}}"��,���F������Ʉ�DR�*�<v���5m'����tb�JK:#��+_ĭ_�g�C1|��?��Ds�/*pI��;f2��(��H��6&�?<�	w��W��h�K���4p���3.���1��l
l�#�=L�ʵ�;N���~Y($@�I��C�\��%K�w{���Ɖ>Qwө&�&ѱ`!�|b3����`ͪ3���ڮk�}?�~��*tM��G~�����?��E+1<D{��=�����f6�'3���Ї���p�]�ٛ#/�.f2Yt�,B�4a�}X�r����<���"��kH����	�_��ؓ����w���ށ��{l}~��m�9��f�cU�I,�R�U]�n^;�<��a��ԩn�Zp̹γ(�׊�q�+�8��WH�2f�<'�NLo
u���>�����A �s��:�_���S��1���?�����T2^���T���������w�5�X����Y�{ܘ5�<շ��{�Mф��<�<�����Гw:�ΔL���4��Ww�gX�8	x,X�J� }�HQ ,����t����R�{��l�t��s"ׯ�_1zeK.,�g�U�J�|�CW�ҳV�������E��ad��p�=��ґ�Ց�	�;����m�w�
����#�`,�#۬�l��h�LO�4>�&A���@X�+�PKѨN��g��h:Ii	�����8ڛ;m��cq'F�c���]&�F�lZX/2�".����Ra��4���<s�i���hX����o1S�aǁݨ����'ư`Q/�Z��B��p+.�KU8�-��ea��U��=�T��Ձ0^�7�21��J��R��뙰9`��}�O� �4��k�(�c �}�Te%��)4��)D=�5��A\��Y"���|/�[�V� xd�.`��9�L��(=�u����$�����ܺVEu@Nk���헴�˫0z������뮓���]����O~�Ǟ}
��V�XEb�1 Ë��8�(K�7a�o�50�s��΅P��Y6{�,"(�V�
�FD����KY�8e�O�ۢ�:3ME���e�vKҝͲ��o�%���䘘��(������1-����?�{Gv���y�ф�}i��6jD;\dy��^?
��F�D��b^දބ���5t����7|^�6�u�OX����
�fR�ق��/��M��F�����w~���#�f�tU3��|�������}��ɱ�69�q�+ ��Kcf!�v&or�蔔pY�˨U,�8~�d�;%>7�e#�1Hf�iB^�@$�����m�v��Y���0�o?�aIG�:r||T��.����]Hg��+���AT��餺N�����u���KW��λ@��Ͽ�/(=]� r%��f�La:_��U��w����	p��c���J�eI�I��K�q	��݁�����ϯ~>���q��!�t�y,��J��j��H���F����\�^��i��׼>&�u��Y_�ns���KZ�����c!?G3�^�_��,����|^tm�����Uy<~k5���|�S|=u̚��c�0�c�1���5��|ԃ���_\�{�Բ�z2��~�14���S��a��z�O~��Ng�����UɢfN#�/a�F�i���F�E��`Eo0�j���0�YM�,b������E��,�@��/G𜲼��*���U���p��^ ?g����
#p?r����n��'1a������J%�΅툴6b"3-�����NЄ��C{2xL��) 0�nH�i�����d���𔝈���Wwkd���0���#3	����	t�tI�{ײn=��Q��{��?�ż�?'�Lp��SoS*�.-jx��)�h+;b��܍7��Ge�~���Ń��8б�m�e!f���A�	�0ߨ�,;(���)�[��[v�a=�Nas�!���QA��{kWǼSiêb�����¦���w�:��Ì�w��0�*�	��-
�Ӂ�]�����m�&�|���[uoB�dj���Ȅ����i�t��N������#B}*٤���& ���׀i���=_��%m�qyP��b���~�#����a*�E�QE��4�4q!빢�AV�Uh1�3Nk��"D�C�"V���L���ж�N�\oF�Gj8U)��������b�@v��#�4.:��+MJ�0���?2���.L����C���	KWG��`�4�0֪���/�J�:�^�V^@X!�B�UFSЅ;o�7|��E���?'a-��dq��'�	n��Y�)[���Z�:�|�Zlٶ7��m�U2�ܨ���ុ���/;[ ����Ii�F� �+UUe�Z�+hjh��N>�˰TU��`P�S&�ƞ����tho��2�8!��֬Y��{�a�i����
�\����k�?+r��_�§Q,e0��@�s�^х��Ϸᩧ������V)��<����3�)�nI{3*U��)K������8`�܈�-@�4���Q��c/��ObÆ�16J/�Q>L�/'���ݳ�=����k�� >|��[�*Z:Z�rY��A��VTe�քrC��J]Qm���zT=�D/fi������D���	���^��K�'�w�J���lQ	��?����n��@I��Gn��Tk��O�0}�zV���Fl�ɱ`���    IDAT��c��5�N��tV��5���:���]�;�g~��m6'�������y �[.���|�l[E!i�j���zY+��9�Q��`����35�]�_���UUv[�s��%�:8�Iy����Ԍ�2]���SU J� 
�a����v5�$|n����t��߾'l&L�#5�OG�m0C�|�i�V����@cg��0j��'F�J��:�b9��^�����U�&�����*"}�D�0م0A���0R9q�İ��U����5��8Cb)Ao���V�妐u��s[�1�\���Su`@!UHW�b
3�+U�<�o���X3��;��>���.9v��w^z�58�~a��b-M"ȟɤeѦ���0 +T��T�ؾ�K��Z���J5�Ac�W���$v�DR a[@�Oz�_�f�	��0G�����iA�&i������6c������N!�
Gm����g�(Q^{ש�}�NP�`89�fSq�HG�3�z�z�]�
x��&�h͝^x,�g���w�#U�H�;�v�T�5��8=���V��w~p{:eM����UC��`yK�4�����Zt���t��l�nj��"����(���XbH7%J�=7)��bG��*�7}~�/��ל����]�Tj �E��մL5�u�&�~T�\y-�S�� /@п��6�(T�<�fU* �cc/�b��c���%��� �y�Wp�m�"�������hn[���~�j�M ?��*��t��ak� ��{���q��?C����n��-��ƿ|���AӋ ���,	2A.D�1�0&�,l���@=����O��Ã���N�~�<��R����3O=-�1�`��5x��mx��X�d���*:;�1><�����q㍟D�Ɩ5�����~<���� �gq�����%�x걇��Ccԇj)��	��Ma![�!)j�)a�؇8�@�����w��^91 �c:�E�J�U:�-�B(Z%,[Յ��A\v�Ÿ�C�����x��mR��j�xC�MU�֟���T�����,���c�s��K�"]�������
�ۻ�\r��SnT�"3��Ԝ���ڦ�� FN=�X�G|^�"�wP���@N��H�(�7���K���88?~�\���ta�r��l���y�j�Z��p?�?x�6��o�������Y	�����YL�f&�s�����0����,�ZB�\��K���F�Jx��r�ªr�aLq��jEE��Ya+��Ц�e���G�L'e�{�ế�MQ?�BR���M!	�<ȹ����<'̧c~=��Y�0?kF&�����ӥ<<��0VG�����Na��&� L�>��>`
��+���# �0��F[#������Gjh��65"�AEd<�*L��J%G.:PJ�е�P����
��7_�3SD�%Ų���e+�Eq��Q�ܵK*�m(9j5ƄI�J�Ra>�?J\������ӑ�,�N�~b�j�� �_'���ҩ�c2��t�����2q���k-���M�LtvUp8fw�Z���]�yk(�������jN�Ŕ�t�%�f���L���Źt��M���� T��c�c���6��A�Ç��$�Je�j�3�)aNo��X{�<��pbx�^z�p ͋�a�k��Ǭ����T�%���A6�OI�x>�w422�҅^�Tu�U���B�/MWu�P�]��4?�&X���1ڷH[M������d�-���R�b��ԩb��!㘡w����'3������EM�) ��Q�Q:�S@�v�$UD?��\
ǆ��UB�[E�߁��3ؾ�yl�������5E{�b� �� ���n��a���a�(������g�r��� n���p��c,���x���A��v�_���F�L}9zXb#�[��[A4�A�Gx���r�R|d�Y�)cZvǫ۱t�b<��fD���A@�Ykο���}^|�5��t"�.b||�bA�����_#_��?�t�+�wbϞ����m~d��x��X�����)�jo��e� F�L�2�nX�K��
�0��� z���	|㶻p|pP�k&G������([~����B$�EbrW^q^|a��o��$�[[��ەq�(:&[��J5��;�A���5�>�FBֲ��Rd?GgA��-����d�q����\��?YYDHRh�ǰ����F��Oo6����V
��#V�N��������/R�A�AX�1�Xi6��=
�)Z����0
�y��~��3ߩ�����M�Q�AțÆ�m�NFs���]~.4�������S�*�j������ �^������ieApfWH��qD�U�}ӝ��deB����b1��Q�jى�3���_�a�{G�	�qCіY�`Qj>��#�1цM$UJ��Ie� �Z?
��A� ��=Sȫ�⤭�a1�'I��MXt�J�'������!5� �!�;�v"���*���V�%�d�"�ɷ|v<&�]O�B�&�eHK�X0���NՃ��^��G����L
��4b]�|��B�ۏt6���[�t�̄YT�V����1�Z?�/��TC���z�S���#��:i���^a4�E����&�L�=f�o\���jk� �ƊF��z����C]Y�cr���x�.���宓�}o�=��֛i�& ����AU��A�>0��nX�{ճ�݂��˪=~�C����	���=&����7n�\z�۱��<�e~�ȃ���Z��XCc(er(N���Z�a�(֯
 я��yS�'�@�*��7���-[���1Y(t�C�B��D�V+����z)����t$��y8��&M���p��l���x�9�x��P���\��ȳ��lVi����#��J%)�������%��r���`��^d�i>
%���1���t��)l��^͉��A�2`V\X�j-��r�*��3RuI�V�3Zq#��c���ع�n��;px���q�Շ�"��B�&ڵ�4\�����.�<��9x�E�z,�E�g�y&vt�<���2S��?�[�n�µ�~H,����X�r�[��w�~�9�L��0�>:��Չ��Vছ��i�+(��^�# ���!\t�p5\v�[����͏�U+���A4n�jQ�Y�e%r��)S�FVר"_ȁ��hĪ���1|馛q��q�n�4r�&M�''ɬ5!��d".kB ��������~�����>�H�"�\>�d�[쉴�,͜_��l&R����5��D�,��;�ްi�?S��s��j�i����Ɍ��e��5����Z�A�ތ��ÿ���Mp=h�g����|&l>��F m>`���T�0��c�F�U AX� �aJ��_�xS@}������~����.8�Y�JLÅ��jX�0#;�3���o;��4��4j�����j�nc�"��z���̛�r�t�W�|���p�l���0�jp`Z�g��b�L+�VA���Qu#���� ��[,*���g��f�a<�0VG�~���b�kj�'��YM� 	�a�0źPB�*Щ�h�OF��@� ,������l�!�ٌE�W�Dj�%���W4ހe�W6T�A�倗��e��Z���Q�+�xO�c��	�Y�����(:�[�N�P�La���>q�FO����L�^�J�1����Q�H:2X�I:�[��SR}3Y�$3�5��`����)����M�0^?����3�L��4�*E��h&� ��X,��P�.�����S��	��7]-��]�����ےiaZ�`��D�GWb*Р�Aa�w���f��AX}�O����EkR�O��^�������� ����n��&�R3�W����;���Mx~��p��Xz�j�
`�_rܤO���.bi�.S���f���z.ۍ��3)�'MMa�T$Ҋ��*����	2,0��&`������4)]A�C�bl�T�)�������O�o���{^{��x|�S�?>Oo'���5���yl�Ф)��g#��4k����t��҃���<�n���1e��
81zV%������ ��V����ҙ<9����t#W4�	k���5�c�j��B4܂B	Xе�?�_��w�X6��gu��%����)ƺl/������R`��!���L�������UW\�+/�L,n����)�}~�{���矗v<��br|B����;�z�j<�m+z/���vc�s����C��K_�W]u	�ā5SX�CG�����3y���l�#y�47ߵc+ʅDÔ��p�k�7�.�p�_���j#��5G�W��=�q�W�.��gd��\��,l���� <�F�e����Db �|F�`/mۂ��#fR	��g���2� h해�Sij�Ԍ�mJ���f�)�
�5������&�7|�.6n<[~�g�zMH(&n.����k�.h�I���R	�u_��xh������S�`���Ǟ��Mg��W�2���1�~�7�U``�����A�0����K�7�Cٶ�Gwn�ѯ����4m`:�R�A1?�x��q��S�՗��s�������Z@�QEU���5E��?��B��SB\E����ޕ�©��'s������b{Hq����@١���t�g��e��%P����k�ܞ�IU3��GY8�$�I`XX��%�����D��+֯��Ԅ��"�u�%��	c� ~G�c�F�cp<��y-��"F�_ݍ�t��(�Zл~��r��!14���D��Y�yg�x�4�(M�]�Ņ�7�)1kC{��SY�����ϙ�	�h�Qe�6Kt0�` �ی�/��|��tcb|g�� �HGG�E|ﷀ@ɀ7[��X��ȚIf�����I�A�B�7�~7�'����ɩ�q�s"F���q�'Zwp���E��� 	s´_�`Ο���H0�L'���z�a��g�q�֚/��"�¿���tlSE�yhRH ��2|�Aͭ��:I���k���>��
���:�S�W��?ٳ���`8�
T3a�����?��pŻ���.KV��d:��;^B�&��M�5��45kbM5
�,\�~��0�����gOD�#��I)_𕜙�j9�T:�'�n�Xp�����
�rO@S��Z!��9�k�Tb[[�g�[��U#h|sV$�E��
�a�ڵr�t@������	6���S �ׯL����e��=#�Q ��G�`H����I�d�+��s�����jÎ���eˋ���T}ǚp�[Ηc�Db,j0�L���d"I�x#~��_c����i��������p�|&+��Y4��"~��E�V� �+���}�_z����&L̯��6P�B�` {�챽��F�Q�Ν���#]����w�'7c��]��H>�W]�����)~,�Jw��-͙ޠ��JO'�k���8�܉ư-MX�T�%���}�eD�f��D�,��6Q��G-�b)�������_�����yn�y��x���G7�,rL6�d�XqzL�շi��G������L'��eՆ�G��1Յ�k�!f�{��H�]��W �c�s^�U���l�����TbBR��h���2��r����+:}(���Lv������2��C�i6\�e�u}��c�
DiF��b�o����N��*9����Z�V1A���p����0��cg�r��~�����2
�$`�;��F����+����8��,��*܎
,3�����^V��)�J��l;��wٹ�C#N��e�H�m��FG'�Ob]�4dц&iY��"3TM��e����9�}a�ɶBb*�D�d�(�us�X�"�Ŭ��Y�@�p�Xy���0�dDX�N� ���7����T�;w�z{�`l|~6�6-AxL"� ���:j�<.�;䞭�Le����X�q4�u� ������HM�@�=�B���n$F>��o��n�J�J��G��1-X7k�G��D�2�e���+%�U�X�fF�����4ad�q1�8�(e� [&���`*�J"i=#?�,�Z�c�T;#������`�5��J�v"g�2��#�W1Lm�Y	��8aY�M�L�s6�-��1*�i.�t�惬
����ES
�Ҭϙl
�2.d�t+eTjJ�� @�B��A�.X8������%�u��J�;����B�sy�{���j�"�M������`��5��=��[�����+c�'&�}�N���5Lͤ��֎���{��_<�j*�YSi2��K��1E ,���# � ��h�޽r^L5��U�d��>��\��T�;�Qb��pAc_S^;e=aJ�b�F�&����H���|���¹��x|-��K(!=E�7<O�C>8dS��Ƚ%��S�b#`�ŴJ#hz��O���/(n��J�Lc`|�b�q��� �a���&Ǐ݋a��B���dG�5�]Cb��d��ҿ������g�'�.'ʆ���0����ȶB���9�ۅ�t]��s�p����?~��Y��0�F[�$�9`l*)ը'L�2���æ�%���]�LL㢋.F6��믿.L%��V/C�J�_E:<����^�hT�����sxוoG[s�ozA/�y��L!��j�Sf!,�Uу��8�AL&���]���p�����[���!�J#���M�9�Ŷ�Ʉ1��ֱ�]�����{���L��w�~j��g�نƈ\�\fν��V�)CQ�͍͊[󦦒b���DP�MS���7 ?�|�^���~���e�-WT7�yJå����5a�1Q���?y���,|/Ƕ� >i������1l���كS�8=��f�>�!�z}�����j�e����W�=mS�M����C��?)&�xd��Y_��'߫�N˗-J	�90�޸���>�!��Ѭ՚��7�q^	�0p"Pw(ڮ(�7T�+i#H�*̀��z}����J1G������2slo�xV2Uwhl7������7�_$"�8����"FIA��C�D$D�V�^|��2��I��5�vTZ�r�=�h�\N
y������n�v���Uq�U2�����0-tuu���	іf�E�ǎ��ԑA��.�TI��Eȡ�l͂�
"۳���Ւ�b6/�U���(��xpYU�ۙJN�P�cj�����ejG�����5nr�m@E>��'�
�=���a�~��9fc(]���LO�L&˻Oᗥ'�f��'+ϳ>�yb��b��Qc���]�c��8�%�e����yH~W�:�T�~�N{F	��I%r��Ur������ ��g�o�H�PUm�A�\����0�nJ�1zch�������;��lF�5���FbT�֬[�֎v8�':?j����*�w�bIs�;|m�-�x��ؾ��\>x*���U��m]��"^6����}Q�Z��8�k������W`�͖_��4ȢA`�Y/�dWU�vCd� ��F�/=��	�8ι��I3���j�UZd��P�
J��y4O�B�t҂!��Hv�x��t+��4�� �b	9�&M%UJ���$EB,4�}Hgg�G�v��4B�Θ�3�0� 1n�s�V��F��¸�l������{ ��!9��/d�-W�������h���֭Z)��d�I�E��љ����;i���YF����)F�4�̐2+%ÓM3��Ex�^�O���W_��������G���t�&�m}
M1���\zNGn7Oe8~��<�l��Ma��(�xy�X���ع�����`��cH�rh������� ���na�H1������W��9\z����?��c"��4��YҀ��t>wX���|U�w�Q�.(]+���dJ�U�%㒠�׍�q<�\�W^�ND�a��
C��GU��$7�������_}z��7�z]�sz�X/��t�o����阬__��ة��ͱ���t��p��
��*���)�\x��Ɂ��^:�w�⾊���[C���p� .aQ�]�⦿�s8��#B�H�-A�b�P�Ta9�8��c�I9�s��s���?�    IDATK
�vџ�Kg;��d���go� 0
�k�c7+c
ES@�����ڥo�S����_؅���#�B��)N�{NJυ<���a�jY@���D2�ƌU����@����j��۳�;X�5��8A��9Lu:�7���*������ڌxG��䨇�T0xt�Ǉ�jE0���sV#a� Uʋ���ѩ0�p�a��D������*e�H�� !VF1e&lRUi��D�Ȕ<|ݵպ-jVc�]�Y�@[���0�#)�ݪix���u�]䈶��j���9o]0�;(���gGNTI�̫�%�¿q��E���vJS(O�F�h�w\d�XW��Ѭ����ߙ�de �0���x���1����s�^Cdr�(�QЪ�A���3aev.��l�[�9�*Y&���/�Ub8��y�q9�d��)RWD�� ��+	���K���f�,�8����0��Y�<~�ϫ6(S�6[��O`L��ׇM��@���/7$�-q=��cGO��Cg2�N�h��Kj�x�����=﷈�3ax����7ۮ�cBZ�ؽ�x�x���Q����I�����j������fhY5���b!o�Ӳ�!}aim�]%LKWL:���a4�� ���*�X�F�e�="�/�j�y��7t!�̣��"�&��bT@X�sQ�0�yQ��"70�8��wt �؈�0�@)�Gs�A�����0�� ��!�bâ8���j��\,uf��9W�pRj�^����ȗ�J� [("��BӪ��H+<��%�sA%@6��M#ͩw�ޅ�Ǐ!�J���/ߵW_܆+��6�[���������~�=Δ�VS�e���l�ǧG��aZtշ��w�`�	|�K��I�o��]�g��,���xB�;��t��]���n���c���([y��3HM�����G���Ç��N�|����&Eu��b0p��X��8�y}	��`�+���6ԤX�]�J���-Ob��tjR��y�I[��5��̓��h��7b���N��u����&����ӀQ�ou=s�?�Ճ02aR�|ǯ^:��⾲/.�H��;�4�L,m�)|����#�O5����3�9=�ǚT���G�pHI6��Jv�~}U�_�]��`k^RSS'���N1�2D�c�q`�dj`��UHN�𵻿���"f�LL!����2й��{U���a�&,fJ0�Df��*�q�I*�2B.z����;�����L>����3���tN�&ޯn{�4��������u��Ibj*��q��A���m-Xv�rLYie�0݆8�P3�3t��[��x�pQ�̇|66'pd�6i5Ķ�k�0C]���b�\g.VU���M�(Z�1����>Y $�\�ؘwv�&�VS���h�I^�n�@�fF5@�B�����cAW�Q�Z=IG҆#�l���/��@���f�4����E���@��C�M�szC���Z}U�;�V>A�q*
���a�+
��JTI�ZvjRګZ��w@�{����-��F( �k�v�zL%��P�E[��wȋ%+�#��[��Tn��E�6̌'h뾑rm����1�NP#-^�6{H�JnLx�x����#
<󘜇d?�:1�E�-�����Ӎ���Ai�B2�N�s���L	���ػw/�.Y��}�ͦ���$��ƾ�ρPHz �i��!�̒�^6�p��2tF0��>��9��C�m`�,B~�=�E*7��&V,��N��'&�s�Ĝ�Y�yBO9�Do<�6�L �4��&l&���H}������>d^X�=:9��9�_	���OX���K�� ������o���.�{�y��/�������r�j�'{w�9��Ҋ��V+֜=�L��_��wU���y��߈��c&���s�B��Arr˖t�*���F6�BE�.�(�����\�@��7�c�8����ڶ�=�	�|�p{����F[{'����|����>4kDcS�F���Kq�����#�f�j!���Xy������}�x�.��K�=��$j�֙��m�t�2_2���qQ��)�܋/�{���ê?$�n���H������ �ڌ���L�bz3��0�N���5���Z|��������/8�9�tV}�����=N��Q����&�O.��ٶ#������[�7n(TȄ%�4�hl���Ӌ�Z
��Ȼ�Ɏ�Q�D�YAt1O��f�N�<x�z�.������7C��mc<���T�ݢ��0��hGk�U�&q�(��@1�桍��J���v���lٌM�w`��Ym6�%��c3�i������:k�"+TJ�^� �aLgӘ�gD˒n+W����Բ�T���(������t�Oj�������'l]��>��s/>_@#���������܈���F��M#��V�[k�Z�1*.�YL���X�l`��-��h��@r:!���Cu7�<
�-j��(��n�ށ�dJ�<�|p�i>2<(&2����ޠ4�$0�K�)�F��Dק@�N_�{8��t�A:�Hk���L��H��~�5<��+#ެ�Z.۶����I3X��(��c�v�V�t��S�mg��Ts��ݝ���VG:=�s,�T�������B2��ZSW��#c:��%Ÿ]�~q���5c���سw�B���J��Q��g��t9[@Wc3��v!�̈3�2'����v�©l�D�E��i:��mb\*� 畵A�JC*K�S�Z�7"0�0d1\�b)v��!כ ��՚;
�y�y_4I�	5:�nd�x|�r�'������p��4���ȑ#r�M�yVM�\�,6�
�P���0,�*㞕�#�C�<�����a���ho�à]�QC�i�
���0�и1>�Eb*3_Cc�C*���KM��av
�^�iK&�م85a����+�YTAbj
RH�*N;�,i[�6�p�&��//�[�)�㵝���14:*��dl����IA˖�6���ƻSb�@�l^���<_��ga���AK���b�p����[��_�]��8~�z{�Ϯ��l�w������e��Ie�����Z:�����%�~�j��흽����+{���]b��ѵP��i���k��߼�6lټY�~���l��-��nĆ��P*�`�r���Gg�ضmz�78t�%S
}.9nY��F�(>��e��jE�T��	�&;.��ߋE==������2��[�nZ�"y\'+�ŚB��ҙ�����엮�<ѿs��c�.ұ��ԃ�7b��k�k��o��u���p��$�GK��u���}v�� �>aR�0Ǐ6|��?����P��R��R!	���Vt��UM�s���~8�\>C-�*B�xv�|���q�RM%�I "V�^�mތY6��ŕ�gM9��w{Pr0`r'/ ހ��0���a`<1%)Qw,����7�|0YEBA�YU=&)Vc�H;ɪ�p0�����a��յ�S9Wu�=ӓ�FY�E�`2!��M�L���ls�� $!#���@�Q�(L���9TwWW�U��~��S3�^��������J��y��k��6<A��<:z;�oYK�,��2ʅ2��$&���D�~D�ALNLȆ�񹱔\����1x�ni���gM�-��JҀ�����&x�n���ʆ���152��|
!�/f�ѕ-�0SH!�o��MQ�H�Ii14<���Bb1��E��������L�!�L�z��lz���LlCU)��Ʉ�~����m��m�٪hnh
�W`)VQ-V�r��S�*�4\�-�Tv���uՋ��YO�ŠiFLI��u��Z�J ����ڤLA�r�̋Js)6T���y����C�N���b�gij]/ ���5� M���i��3;��;����K�giʿ��y\�pp��1auYʾ���k�n���,�oZ���=GX0�Nx�"�s������ÉJ&��ۇ�`J����2��4��ׇf�	㼦9Y)�=�摦�f�s���5AG��ԙ���m6aLer3���2��� ��V\�5H�)F����x��9�y_*��.�0"/ܼy����c�ˁ�Rj��a�j媀
2f�JǇ�a6>���QF��@{c"!iv��	T*6�\��9��{�D(;�sEP��cl
TO��ZVlv�4t��
#N���j���G�c>[C�9�l�CU
K��g�н?O�D2��_�~��_���oGCs3FF��W�� �o���]����+��!��瞋}�������r���"x����(R�2~�����'��[�y%xc?�ŹY��_^�ΎF���K��V�u��1�(!�e�<����Ǯ��hhl�%_���t+؉���;w�AWW&'ǅ����싋��z���W�U���B.�.�"Vėr"���Ǳ}�c�UZ�lv��3�#�`��tU��ö[�\r��P>t䰴Sr���V}+z��7��`@|�t��b��N�&�Voa���eZwZ����$8����u���0���̊����0�����t�������5T��z�_��!��Zl��'�e�,7����7����!к�5u�0aa��]h�����Fj����R5X)8���w?�[�{t���ȢƅTU�(͎���2���O30�ᴀ3�e�p�j�|^�P������Kq�#$�$2Y�i=P-��JL���r��o(�9�0�(�����%��*���ndKy$r4{,���4FC�怣 ����j��>�A6���.�O��='�8)�:����-`��^q���zSӘ�����B�)��QB��K�"RբXP��.&�06���2K�imcs�D�-��R�:=]'i����xb��s/Dz`��X%���*�����l	�X
��,gN���jL�0aJL��Mв��w�U9U�~22R��k����ӈ�:eō��qq���#_�4 s`�Ľ^�2t�����`�	��zVJ�g�d���'MWO_x��Ӂ�6/�ݲ��,|�gQl��_��ժ(�
�׍�[7axt�h�]x���G<f�V[��YZY-�	#[��.E'�zv�Q��Rk�L0����n���7�-F�:m��|��JT>�`��#&�ubp�q�0��b�%ϹN��sN�Lijo�7�2^K�%3���?�A��Y6���0o��s�<�1���X���el�����X�T*�=T�H?��0��%�6�����KX��X�`hx�}��x�ٽ����a�#�Q�nQ��>��h0��l���˟:&LX:-F�L�.�Q�/`Ŧhjj���l5g��p��~��G���{����W�@wOr����i�x�;�)ߛ�<�����T����`�k1��G?�A����	V���Oa>D���3��[_�6GG������E�tZ��^�7y�ݿ�Rbl�Ca��踴�)W,�e��]��ʢ�D[��܁��ٍM��"��bhdD*�y������:�08؏����돐����yJ-���Jhi��V�������L`r:�l&��h��A��i	���妾ל���يP2�x<!)a�
�2��<��T�2�֬Y����-bO��'�_�>(��2fb�M����[1j�[�g�Xŵ�ȯ�O}:�~=�g���(��z��R 쥘0���<i���}<'��U�0�ۓ^���x9ZT�x��Ko����,��u�#��Ѩ%�p
�����#;K)�
X�b�������y O�G��;$�fD@�Z�X��+�z��1��$�y1�k���"� �]��XY'x&��C�e.�y[تVi�CA����ی��Oz�x=�	�
h_ю@؇L!��DJ�;TS�F�#���I��-oÇ?�A��=9��x�	��]�_�{&c��/BLoa�*4�͎KϽ �F��W ���G���4���kU/f�It�_��׉{X����8�{��*b�H�ݽ=hlm+.v�@GF���BIQ1���E*�r�7[X�Q��rR/���f���D�7�b<'ͻ�U�dZ�f^3�Ubr��J}Ճ��b�ꅯ�R�f۪�J�j�7t=i5��d��d�h��udz���%#��$tP��׬O��7.p⁥���zSp�7qF�h�}j������5�%q���U�<^n�r3�T(��,��G�"��H��8?��%�reK�x�k_+�6��XU9>9�l1o( @�=H-�2:�M���M���0=i"i�0��\N�Wmm-�XQ��Ҍ�-tԮq��QZ��R��@��2P&SF�:j�y�x~53&�L�^�)L����z���ɞ��);b�|�rq	�r��1�X�8߃my�Õ�Z�ui<����KgPȕ���.���8���*�)lGwk�Ꝙ��Ù�^
�ӏ�~�;�Π���N�b��#(-��ا� �&Ֆ,6R�|��gυ2[�ŵX���O���������]�=n'�.'<^'c�,�p�?����Y	�Ãؽ�twv�8��&,�H�&��������YI��⎻�g������3�����g?�.�d@�Hd��3�b����?1��/�Acs+2��	�\Y�zV� E���W�uW�?����[��9J����82����_�c-����Yj떖Ҙ�����b|^���M�tdzj\R}W_�)\��w��8��!�r㹧w�y��ݵ_��� �"PC"UPU���$��:h��4�>9q�AǔJ��P��J�q�2�rz�p�쏌I���|;#Q�3"�im�$)����L[ ;��0�+���ט�?S�F�룞�z��ڳӃ@��N&E�ԃ,�J׃'�Ω���s��sRϷ����z�S�}|�`y��v�a'{ ������?���Zo�~���M�`�:Fb��a�,!�c}���8>��+��M�Z\�ը�\2�*<�&<��>��������m����|�j�
�/��h�*BI�U�@�F2U!V��KVa�~��Ve����B�=�}j�HSK2;X�.|f�m�z��>')AX��C��nx�.�MO�j�]��-49�D��3_�;��|���lI����W��;����`��l7D��9q��3�7��+ĆǱa�*bb|+׬�������o�;@�gG���p@�b���d��Ʀ1;9-aj&Z�Z��ى|� ���ԴJ��l�	Ff��"��p�Ծ@=�]����'�y&��-�(��E�T�9�y�7 �U�jM�/��Du�K�/�8�1�0V����i'�#~�!���]5 �s�]t��=Lk����/�丙�6+u��z�����<�BAS����/�:ť=֤�M��e&�ߡ�S����H�C�$��9mE`]_2��	����%���ufڅd�a��7��R�862*��{w��_|�2Y��V|��c�cO�."0>Y"Oݤ�܀BA����3�4�0V��ƪ�&dy�uT����!��g���	�c����薬��i����r���Јh������:�p8"L�����b 2�ɤ0a��Z��&���Ȉ��8�عs�ɤ5�q�����Y�L��R���+��8:9�X|6k=�!ثi|�����F ߹�G(W�pz�(U������5;X+CF�� ��8R���8:0�٥�Ч���w�gP����
"jU4�`�����k+�WJ�_�*��r)�����jk�������E[���@Gw�P�p@2�0:4��o������5�V윳���n���1�M��w���#i�>�,2�v�=�bq�Z:=J;�O�K�a1N�k�ebbz
�	47�!�T���UV��f�:47�`�D���p�x��	-z�esI��`ǆ�}�j��}o�����|������.@8��_�*�ܴ.a��4�CR�R\�5Ϫ�Z��|��Hj�,��gf�Ã��S��l��RAZ���x���*�\/صAO��L���UR��҆
�9��7�Է S��Q�.UXfNg�4x;�9��t頒���Cɢ�ߑ�P������\�O[�����s�Y�/���_p�\{,��F�/�����o���m��e��Z�e	A_�\��u)�t    IDAT>}�끥	�*K([��#�d�w+z�y��]�90�IK����mH�H@�d�H�3�}J!( W��d=�_Q�zp�r ���ZG�+5d�%�_qNUdPRਚH�� �J��[ʹ@�Js.%V�a~$�Ya���3��0���`�a<��C��!�|^y�6��Ո��Z�1���X?�M�����Q���s�U�cuW/<���gg�?>�����#o +7�W��Y1�$H�'�e7jY��M�Qp3�/O.�������� ����(�2B�03��L+'	�5���I��~�'k��-=kQXL+�YJ!������������Ց�s�O�0�=*�Ѧ�k177W�p�qs���I��Ao�:b����@&L�j:Z�E�9.���н#���)��i{��R�`.��`��9��a�Ӓ��|a��i7�� ��J��,(+ YAx�9�H�Ş}{ѽ��?����3��	�U�.������1E�L�,�fu�fkU�߳�1*F���h�N�֧<Ȃ����EU�ڤ=-�8��dK2����bU���G@���΂ך:&jgȘQT�먽��{{�:񹚁�q1p�{�y�ʲ��W�5H���UE-�5�<���\���<s�,f�0�8�QDcЁ����/���m�z_��k8��0=l.�f�bp������*�!�49=���4>� 2@Ϳ�����4U�8��ٷ
c���R�fw��
g��)�n�J3l�H5ؒsx�?�.�LǏ��<��Y<�����������E[ml��]{�{oٲ�R��� ��@8� �<���i�:���J��XZL�oxr�|� �ia��6,��I��sfD2him���n��,,�cv~sS��؅�/�\8@Sܴt3 �~f�s���bi� !�X��IA��Ɛ����G?��?�Qdʢ�ǉ#����EC��B.����(��Z ��n�v��P`@�:�ҁ�0�嚌/�[�Oq�9�^�l�1�����mm#ȧ۾a{a�}R�g�X6K�������ꥀ����N��>�h�MK>�uF����1��V�O}@y��u���?�*�������~�e�~���Kn���n��[6�2�RI�f]B�_��N�l	|����d�/�$�9��?��	ܷ�,x�� �R���Ku!����BV&w�]]���|�~��VY1]z�� L�i|�D*�(H�Ӵ������r�צ�[�]X��eY3�|�+k&�CMX��ξ.�Q�Tln_P���2�>Џ�a��V��E�_ �a<��I�����8<9g4����m�D�X3ҫ�=҈��)1Ϭ����j86:��TFȇ^y�4�>6؏��Yz�n���PCS�4���ؿw����Q��ni\� T`V�_3��Ϥ��t���\̨WK/.���!5���ᅑ�"`�"���ס*-�B��`V��4�Z�NZT�G �d$eVĚ��ZO�}��V���q�U9��,���&iѶTݙ&��|�}�f�����v��T0���<g���5�&A�7T��Z��ȱZ���[f�4��|�;���`���΄,%)�� �hX\�Y�̟�'�f�.�vX*/��(�M���[�G��H�|A��#�Oϛ �Q%�i%*f+)��y��kB4��Q�+�#�*��a��U�OY>���sJ�EA6�!A�b�BƁU�W���	X�FLU�'�����b��GRN�l\�-����s�2���	n�|A���L��aTȰK�"�S�j�A�B,1���\�2�n�u�����%|��kpb|	7��-hk�����n?��Y�4�c��V�۲�R^ie9�V�Z�B���ՋO�:�ϣ�2�L�F���[��阀0��/犋\�Z��R�4v{���,���8���E�у�e�d�*�n=�>��h��b��@�@a�������T�H#R���F9�֯�m�G��3�$��n�d�<�FG�����m�Ȟ��XJ�e�0�j�lřgmƗ��j����������z�LM����%���F�VHQ �#�w�"������y2�G��s���_��/�o�Z�a�;qϝw�1��V��m��ܴbtX�gQ-�$Pb��=o��J�@b��UL��5C����ϴ���݀����
Ȁ�5�y�T�r��t�3�M��Y^GX�
�}�r[%s�/��K��k�Ҟ���:�~�ڬ�I������N�kV��Tϯ���g�N�|���ˠ��'v�Y���I�~���f�����t�}�+;��S�D&Lӑ]t����{��'��+qᴠ�v9� �9<��N$�>��JT�F�%�S�Z���Y��Μ,��d�A�ME��~4����(�e�rS��S�N�V����FMK��V�t�g:�2%�ᄨ CFg�8�^a]���-e0�4�Hc�T4V�e�b)L8�VW��4��Xջ��3�DB��������<6^|����l��J���,���	�K ���� r`j�J6`:���ÎM��׍�'D7��bS�͍���{�S	Ѳ;tX�e��~/<-���"�E�7n<�ДE�mk�׼>�l�.����fQe��E����<�Ky��3h6�${)���hHO��b��A���	�vt_@j�H�3�����-�<I��x|Q|��S��,]A$cάv����ǖn�����|�b=�R��s�]�e\���r��t�����>����%�0���G��=	�0z��I�T+FJX���"\�Ӌ.������0��˸=x�-�X�ыJ6;51���� ��i�o���k-$�}��F�5[�NDmԒ�c�� +cU��+�\Rd"�{:DC��#ׇ3�<[�5?��A���g�)�E9�0\,4mU�fLY�%��i����E|��n�bA�ѵ+Q���^���Y�-MIk����Âsׯŗ���z���ӂ���5b����F�~�&�b®�����������׌/��M8>2'��"�H]�VchjŚnOP:�Tp����J�[��^�ɘ��H�!)ɡ�~���}b�0��q{�� S?��-(����=�ab2��|noH�i0���<���7~����h��T�C*��)Z�h��=�n����yD9�+^q)���w��5��P\�a�P��T��臷b��_,���36����\v�er��D:t����/����	8l�48ԏ�^R����Ł�`X��MO���n����Ŭh$X  ���QF�bUaJcHxV.�9`Z.)p�f�ޓ����y|��͛7⢋.B��b2i�Ɇ��j��׊M�׻̾�o�iV�t V�r\��ԙdk��R��Th�徔��f���g�[���L�d�Jʅ��|*�S����:3�z�ty����p�e�v�j����������q���2K×氡ˇN#�O����ό"���g�UC-�E&���'��x
��N�3�� �:
�f$ApU�:p��q�Q@JEL�p��V|�/����f� ��Iu$����@��@�jG٦�I���C@�U��srӪVd[��Jݫ{O/b~)���.��5S@f6������(l��?�a��ŗJ7�u��n<��v�86oKZz�miBOO��8w�F�ş]� �pZ$�id
y��g��_���"}���
܍aT]Ņ6E��se�
�45�i'7���i 	Jׂ���(�T6����lĬc�-�����3��		�e#���@�.
��v/\e+�s)XhTK��������k2_�h`
9��L7
V)q�����M�)M�s1d���2��\�hs��5'xW�{��_��i���^N%9'�qpt�)⦠@�J�8�iqb�.Ѱ�u��y�/�	3��:Xu�T�4[?G�*α���=bqiI�0�0�aL9Kz�Z�T��I��!�C+�-[����n���8A�URqk+��:�i���Pʼ��Lah)WT'S���+��� �K� Ͷ76��f�r��X VJ�Q� �
�V�ڵ�e�CSS�lf�&���-B�h��n�l�菞8.�������M6��D�.Tki�������\V�Z��V}OZIp�(#W�`fqK�9��i�Y�����|E;p�G��H#���,�ޠ��Rɜ���y*�6+ڽ@8 bn�+�k�����iC�R�?EG�*O͡d������2<��	���k:��{؞�\�bf|S���#�L D$Ҁ�٘t�/�����s�!Υ%X-��q����>��3��o�3���אL��<@[kbqDZ0>9��z�e��\�����?�����;(j����~�:�����o����=�.������_�e�^�L>�Î��Q�	�\&�Y\s�g1>1�Í�6ʼ�7�o|�۰�ŽH-���@�����$�ż�P$,�O�k��T�\ʁM�	6�	��� +�	,�P4}�<[qq�`��H$��.SGF���/^�/ҋ����lWQ�x<w�|o�RKWy��VW}�_{z����t`�u���}�5������y�)K���dv�9= ��H̀�dj�Tϧ��G�	����ŷ�.M������[�i� �|iK�����G���k�|�$<�
��<�؅��!��cpl�
[Y�A�*�g%�lT�P\kK�2��5]&(f
��ݾF��b(HYl��"5�I�L��`bfV�'�$,!d`�����/��ܵ��Y���XrO���bu������vv�-
�=�f�i����^lZ�N�%nެP���3���w��V[�1u����k����k7������;�R.�l� Uj�߿�&i��64�H@�d�%���W
��M�BV%�0<0���9���}=BuS ��y��U�.[$@T}�Y�y�.I]2���r���������腛�ȥ���t��B�D�"`��4W	���M�τ��ϥ#�h�h�:%2Z{�q��4�J7�'���MX/�zHq!#H�sܔ	���t�<^+/;������|�s�O0�4H����P�0o��֙�<o���a�`�S9���2����<a!�;��Ɉ0kSYCag�}�: ����$rKX�֍ٱ	>�h�皖1�銭\&+�HWB�������e�{� ����x�g����9,�rS�)�8��s�O����R�/SP�z�IK�CQy>F?0�"�S��d���\�y���q,�Eê�f.�]	@���5��^��R�`�j%L͍!���Zɡ�����.������.B�N|��$V�H<n~���wf�t|0u�JLz��}���翍��Y���b�@C�V�	+[�*���P==i9�2������rF6��n;PȖQ�$���1p�T�\d�9�"g cŴ���w�w�u�����21j�9p�e���]�K���� ��pff���1���Ǟ؁[~��2>�Q$q��u�§����9�}n�����{1=������s��`1�N��[o�ƍ�q;P�e-�����g�߄���NLN�5"�HbaA1�V���:ӳ�(e
�h���cGP)�D���e	�JMZ)ҧ�GvS�WvYS8w8NR�p�YgI0p���e#r�.1����,ߟ)I��y	�8~E�h:��^է	���Ic'k�U��7�u�c�ԧ!�Ǻ��5J���:K�����#������V�ڠz�ky�3���L}ީ �j8������|Y�0�O�<q��o��M6_�F��Jy�����=At9����oGeq{��"��8�r>����Oh|F�Tɢn��F!�ya�L�~%P�*̛���z���t�[	�5t���Vgf�����a$��BŦ���C\��4{F��� ��U�	M�tA��5+�/e129���vѳU
e����sX@X���u��UlY��'0?C)O��~��;��s�xr�<�=����nmÙk6�ڿ��@G�P#��뮻����T)��K�8XB^X"؂^4����&�GQNe1;1%ƫ�����m��-iY2z�|Vz�QD`G?�����sI�z�v8�J�p����{�Z���4�n������a�VD網�B*���N�i�|T��4azQQ�5�v��9�	�8.�i*(mKPoHH���E��i���"@��Ǎ����qS&��f�|S\4�!�
S3]Zv�������u:��H�N.����S��EJ�e� ��aqI�0����qQ���R��N�d��-����Jۢ/چ9/C��e�r��`ŝ�ƙZ̈́�E��4�O
�7�{�V��D���҈x|QLb�l�q��5�Wd�����8a1��6������ӏ�b>/U�Sdɚ�ZeP�����������M�+�8�yM	�G�G��&5�Ǳ�52r�_gU|�saڊ�VE�Z����Rq�P@�߁�=�x��^��}훈W��|�CҤ{�������vz��Zb��O�V,� ˗K�������c5>��o�D�4\~���PSZW��td�`��6?���E�QpNᴔ�)��_�!?��0�� i�٩q�}��8P����Ĳ� ��q��d�����o!��_���������o���Q��&�M#��G�!�Z�&}l�F'�k��x���x쉧�b��T$^r�6|��W�VcqUN
�f��������A,-�02<��?�l>�������.��/�z��
>��k1?��
�rŊbpI�,,��uo���#Ȥf�u��������A.��j^1���qGv��T��d�Z&�Y78.�eQ�J 08 ��s8�9�Ȍ	Ke��G�qΜ����5�sK�I��׳Wˠ�P��:�̔6�>Li�����[:�����LY��� L4��k]�Z8�z�ӑ|��\�b�΂�c8��|Ω �R���v���0����eeQa�ٓ'.���z�3ص���)�y��l\B���O_�Ndf��9Q̧P���_�!t�pB|f�e�es17����-�oV���D˃�N�e�Y�\(��YP�EdM0���W�2v�x�y�yX�b�l�R1�R�"�W4'�Џ�L,h�
B� |A�T���^������66��4%��4�v��Љ�z�覸��/[8?���W�Ўg�e�;���@sc�n��7��w���E�\D�Q)c׮]��_�lD���ǉ�[����d�e:���"��C��:=N4�6��(�*\���ȕ���sx��q�������@2`�Z^�l�t�LN��i�\p hq�+�#W��P���:�ѓ[[E���#)����f:�T�4A]]�xӓ������Z-.�\�d0EŅ@�q+��r+�`W�f��`���5������|^�
E�{�̹hr�!`���2)��s�M_�ɔ,{U�T�Gel��T���Ӧ�SS/�#���Zj�99~D��� ��?I�rr������r�A�P�����b˦ͨf����3p�2RJ��b�p����a�9�է�C�Ԣ�ttII)q�����	ٰxL�N�hH�<VI�7Ӌ|��ˉĒ����)F^��tZ�>�I��Ѵ�����k�cbU��Ĩ0�= k�M�cE�5���S۞�I�s��d�4�dҔ�s�B���oS�[J8w�*\���'�ݎ���oy;¡�w�"��!��AXFZ�P�984���"�mX���IXlڻ�����;8r|L*[�­-h_ه�������+�����z/��~��4\��˟ �^������@sS6�[-�Aj����Aw��-�٤{hx��<+UJb����,�d��X�C���뗴}����C��]���\#ɀX�(!>�"���#}l|���<��N$�r�FsKʕ<�}�����M`�(���d~l���11C(܊�i�B�Θ���
�G�8�0�A*1�-����t��E1fe��jP`f`�j�%�W[���_�LX0�mW�`^���ҀKg^�Sfd�]I��"im�ڳXp�b۶mr.�O�Q5���S��L�a���A:yX��#�{&6'~c�I?A��d7�>�!}_�W��x���|��D@��s�z޷�&�a��F���    IDAT,��3�kX�s��+��,3�|��C�-�����s�W&��$���<��;���-�5����ґƷ��q���w��k�O�Q�/�i$��m�-���f>�7 =5������\"��Ua�_I.��I�k6ӥ�4�T�aj
���[l1�p��*���NTX���?����f���J��|Ɋ�Ã�� �]�H���bZ�!��)f��|Q�5%(	=���=���B�jM*F�ӓ����H�%�����6`S�j���oK����Ex��U��,n��ϱc�>�>r5��HS:�:�K���K^����gQ)d�v�Ϩ(b�G�{
���OIZ��fΐ�p ����~4�4�vct`D�a^�6��kW�%Ao_/�f������|\5نM��( e�����%�ө� �\"�|*#�z�[��N㯯���q�ztZ#��ʤ`6�[1U�P�q"q��S7.4x�����z�K��I=1}B��EoϞ=�|"�%����>w��ƅ�&A4=��N����%+�M����o��8Q��4����-@5�o�tO6��e+([ma�J�iL�u�o�n(͔�II%��dZ�,Wc)}d��x�y����6$��tM`������[��D�FIQF:�Ͽ �׮���K�[��`��+.�Ç���s����T�&D/+Ӏ�s���J_?89����cI>Y�BQ1���<'������V<.nhZ{G�>��7n�(��ĉS�?/�#�.����i��e�ߏㄟM�G�J�����|�K�#��}�xbʛ-��)�B��]u�(�J*�k��g_���n��Z���p��ߌL.�{~
V���mB[{7ވ���&Z>�$�7>6���drIi}ı�J�����_�tZ�rg�����L�T��������U�pV8,U����G�O����?���Ʊ����ރh8 פ��/}�����q2��[�ē�cl<��9���"��z�F�s�-�e�H�c�.h�����i�F>���xw�y?<��k7��/�������� ��=�p�m�������(bs	�cQ�0����7��gelV��]xd�v��w��	��&�X*�����pJ����p��cbz��l���$�EL���e�K�:��4T,%4��8�֦F�#�k���U��tB:9P_(�ٱ�����m�b��p{D�Y�8dU2��p3�#���W�Z��=���Yh���On�G�{�#�Z@���xbI����}��#I���j���0��R`c���t6#������,��L}1�7D%�J7ZM1 �Ք��Uv_��}��k�dZD
�}�2~�3ҥ�k� g��˦��yd�i�
�aw�Y�v��^�H���B��b����Ǉ�j5���v^��_<|}�}�F�ˇ��	XJ1�D�X�tF�ؕ���쀳RFviN��Ak e0gs8hէ�4e*��ƄU^:',�i�h͑M9JC����LG݌Й�)H{[���͋����xl`
���J9�e��N8-6�XĤ�!��$�-��#��A�L-�H�S"����c��8�Z�l�;_�:Qw��9���$�}�����ǐ,�ii�B��p�<�|�D~1�Y1�h��}���o^'��5�+{�U�?�L�8xG���[�I�b�jL/�о��֯��il������_��W��75D��	��� }69��>x@��j�$&��guZ�����HW���(��@����4"��2D5#�����+�ŀF���h�dA��<�Z�U� o>���Ӳqp��̈��Y�q\��5܄�(jDk�tJ���U�C�^���8�5��Iv��#��RU@ S�ʳ�a��U:T��1��*0�E����S�6-�{3��l��-W3S��0��hSR���Q,U��)a�İ�O<ޭ[�b`h��3��bw�[vq�]�A6���ԝ,{����q�t��q��v�ycp!�T2�,��"e#a�p��`[�7U��UkW�q��O�������bA]?�1�s>��_�y�.���I���?]�A$A5�a2e�*J�̮kM~�@���Ӱafz
�\�v�]V��&���o�}�jǡ�C���I�P�I�O��V�.��#�� n���`���.g����cp|N6AF�pm����Tibw
�5���-�i��A�E9�B|�ZW��v�Yxz��͌c�;�M%Q���L`���:#;i����e��D�(��Y.8���Utw6���/���_<��w>��������԰�y��I��;$�J=\lvg��U@XK[���p�m8|�h���cx��¨�"���| [���j��bC�{~+>k?��o�gQM�=�/�t�w����E�K��lV�oC.����Q��.8$��}�s/0�\����1l=���یV,�=���Y�AWg��!�),Qc[N6�]�cf�~Sdq9�|�� �6�U�)A=W�3&�:Uݵ�c����] T �]�xԅLڬZ{�q��=\��8��0���ȹA�/�.����iQ>����DR`�v��%/qHl�]-�s����D��*h���uC��dP�ӻ����l=�k�����]:�G���w����H�f�B�͌��3{�� >�Fa_�̇`ϧ�f�)�E6� �����]��T��Bӣ"p!�jd��5��e���ǋ�Z3U�#1g	=Ū��J������e�����x�������C&�X9/e��]@+�$��j3��� �°��JE�n�rI�/%$�шpt���Xj���n|�k߀Q�¨YP�e��g��y��ȣ��=�.��u6���[��UlC%��ۮ��X������ZV�"���f�5,�/ _BljF�*1�t��	�v�4�4��`az
����LK�0�v��(�j������|?҅�169�l*�ǅ�׏��6x^>�������H�D)�����IG}Ō��)&L�#��_�/�0�\bD�IJ�G���2�0'>�a�L����y)�_\\� K�&sF��Z[S��.�\ 86��R)D�̅B|��'���{J�>�Z��=Ƿr�Vƹ'��ja�|/2������A�0Qf8F]�D�ZSa�
�p��a��Q���i%Fʌ^���^a}�	f8,l�b:	_8��ج�Л��l퀫XCz>�遶̄�����-4�㲲R.�����hX ���0���r.j*��E� ^��Yb����&�Ug�b�Y�'$�I��A�2i-/����5Тan�7��L_w]���n@bI�+�e�x�t���T���3=�*�X������#��:��q�Y���׼m��'�x��p�P��!ܼ�,��tH%0q�"p:�;�t:��E	�L3s|�_���T���_�A@���j��a
`������k3S(������u}�3H'���M���*��Z���zq�w��v�<X�g
w`q)K�?��~Y���5�|\�+[�%�p�yga||���َ��%<�سp�iEҀT�թ�����?ۆ�xt���Vvu����=�;(���s&֭_��~�ALLNcrb3�	�<z���\��t�d0;�{�eb��N̡V�F63AƬ�!���$#�`� �*�1jH..���4�%�~���M°��q<r�g���x���֘п�O=��HL�������h	�@Y?�t?���s����`IK,h��1͛r����c�s�s������D�*V��1��Y�-�|o,�P���a�4:/(�[~mq�c��y�A�+��/�֙�<i==� ��i���|��Uk�6?���^V �'�'����[?��K5�f_���Ch[�v�Aw~c��h.:c�L��2H�ϠZȈ6��4]�ij.���^YjЋ�[{�,WJ�e������z��hK���3��+_���dﵼX&X��v$lN�t���=�B*��r^D�n�X���4�AX�R�?��턥Z���+$�@��X|I�F�a��c���\!\��|�+_��XC9_�ֶ�fL�O�o~;v�3����<�Y����+�=z5���Uų�=��ȓ�K�5����mE�̪�E$��-%a�d�]6M������+����R�1x�D��ZI�/����lp�����,� ��� 2NRF,�W����C���QC�a�ؚ-#30'�(���p*�V��Lm	��}_�& �,߮OGj�s2+l�+Q"S,�R�5k��j!�����O:�Fg���X�Z��W�u��{��!?W��	�KJ?^^8�"E[]贚�aF���(�Ǣ���&�S���H��|I�Ś���Ƭ��=���T�1RKĶE��	C��H*����_��|���|��E~t����Ғ�+������&T����+�ul"T'�fjXD�cV?��mP��PP��aa�a�u�)F�Y�Je)m3����s��3��w!����:�PU�d�Vȴ�M+��k�k�t��o]��͞yܺʖcK����*ퟌ�BY6UUQ���*�d�T��S��H�ej����E�R@0���7�ǋƆv��a�����M#R\�0U>�er2xu18-��~L���ٌ���z�e��At�^���)IEZ����m:��9�l�]���g|A�aMaV����^������a��=��֭g`dlT$#�S3r=���/�3}Kc&�`��1:>�/$� ���/�[��F,�N�m�gw��s������X+ع{�rH�r���G2�Eg{�-�X��o|��ؾ�Ai��,���@�(jU�lI�g��ή���x�'�N�i���E|1�'��T��C�ٹ����9��ӨUsh��P�-ajlX���!��B	㙆e�ǱJF8���"�"��c��Ur<d�X�A�#�0�h��BH WVF�����/�K���6�Z.A�Ǥf�4�K��F�e+�q^��:�3�q^3J ���^�$ĕ����6!<�v�s�$�N3�5�Ǡ�6>�s���@�,�*�i�4��������lg��'χ�Ģӭ�~-.���/��T������ho�<���u;*�X,/�t$/�Ϟ�������Bmaw"�N�nKc��T�p`aw�oތu�=�ii�Ǡi`^�52���!�a�ݢ�/�&���m�h�,w���͜���b�YT�&{F�q��Q���T��\U',�i�7��wx�G�	̳��G�*L�������~v��Th�H�$jĺWv0�K-a!�T���əy,N������\����
 _FS��'��j��o����P�A��q�������ro��Up��4�U�rT������a��ͨ�������0�ͫJF����wl�4���b�%!�K�ȁ1p�0��4�X��K&�Y[�F<���wEl���d�Hꓞ6Ѧ(^��W�xs�� R��'�9N�]�x�5��yЮ����f�� �ד l�	���? az2jf�������ˁ\Nyz��LRb|�^�(a7�P.n��C~��2$p��u��fZ� h�L�VXf�4H�8�3���+�0)Pk�1Siӆ�5�˓�BU
��3��S4�K3a�̗�SU��K�b�S���Q���O�D���n��ĶmJľj�jˢ�������b��6���[�31q��7"3�̩��e�U��\�t$�S
!�-}��]�n������,|�+u5ܔvh����v���]=¨�1F�<'lbvJpk6��}�0΍�%?G/��n�>Cw�Ћ>?_ k�(��0�����[���Uٴ���>}�l7�9��v�-2{Y)��>O#�F�S���zHf�vJ+X�E.OP��?�vҥ"\� V��( �Hy���5�ղ�%b���\DzvZd"�?�ڛpޙ�'�uSC�5.���#b�+?s.P{�G07��t��������QY�3\�(�dp��ލ��_@&�Bc$,�DW�씞����ţ۟�,S�¨t��.}Ņ�GG{��鲙2��>�d�s.(�c˖MG|��Tm�5�n���T�@(��ŎB�ͷ�-��Wdך52γ�E�mi��THczr>�M�襧@�a�m�VQ�+]%�	��3��" �\Q`���M:08�xR�XI�K[�DZ@�s�=��g������
&r�ƨ Mk	�}�_�S�z�#����s�+����L�k?H>�A�����<��ù¹��:th9��g���;v����3�@��}V�?M�g����@5`�Nz��Lg41#��j�ڵ��=K,�a���6������m�_Vf��Z�����.���n��-Ҿ1]�s����ڌZy�ۋ($�����RM��%x�.[R�2=3#��F��:K�|1}�\�	�d!_ֆ�ǩX`4n���ǆ�hV�J��jGG[�d�L�R	�2�s�Hٽ��O�ā�<���1W+�a�Q�{ٔc�T=�a6[���+�[ѵ�K��科-V$����R��E�#�s�lƧ>�4�(g�
x|������-?B�f�B&��\V��W�Z��χu�=��k��QT�B)���a<��y�|�-8��s�o�`j��)$�I����f��b����[��5��8�����CX�������t��փ3��%fO?�*�>?FFEG�z�Z���t�\u�U��������¤V]�Vtaa¬e�CF�@�ա� L7�V�䟾�΄Ճ0�Ʉ�����A�D.�d�$�-�$}&��4�鞯� 2a��Gc��15F�uZ�����BQ|��1*��b���q�f-Ǡ-U�T��ᲊ�D1o�
��D�&�ǍF�NMG����d}l��\N���gg���>����e=V���Cr엽�X�~=��wf(�g�nѰ"�т�[����fc�Y�h�$ɠ��A3��F[��ﯯ�n���s���$�~gr$�P:'��"
^>���K���Q!a8	���t�ò�(@JW�D�<�����d떏�b���3%�c��q�P�����6lb?�������`�"�[E	b��)����ҿ��͜:ֲ���P+&��D�nؼ(	HC����j�B���'iX	�屘�U���ѻv=�&�A�e�U`��uM4®Q�$�E{Sn�E��G�㶋6�}�R ���7�|�_@�P��\՚�x�_��LLM���+�:q��.\s����~N4�Ԙ��W���F*�(curr7��1��~4B�^�M(������}}+d����V�~��E��v�d�[�F ����m;�}ݫqL�}{��/q"�6i�NFQ�-m��4�*S�jVK	�^��Ec9�,d�����,�o��lJҧdtV��z�h�8�)uX�v��P�-�:�J,)�7'3�f�?����c�c��H� �w]�����Wix<re���N�� A"�I+��g�}V|̴�Bi�U�9AǺN�s��kt�^W�30|�ނ\|?��%�<~�]����{s��%�	p���5Ov������]^�>�3ֽ� �n��/��v���@��W/L���o��lݸDʿZ@���a�6���l�xJ�N'��Vԃ)ϟ�L ��2h
E�A���]��(�`��"��0��׸�bA ^C$�Z1k6��6�ŧ?�a$&`)��fN?o���G��7n������"b�f��V�)fH;۲y����inD����n���S��f�R��*�͍r"���":<Q�����/a}�jу�������G�~��P���c�Ζ6��a3��җ��hkj��\<�]���׿�+V�!�\���(9m`iS��B4����Mv/n���x�G059)�۟��MX�f%v�ٍZ9���@&��7��D�T'k�Å�O=��|�h�:W�����)����ځ��a�N�x�n��[�p���tOf�nMK�M��H=ş�i �ǘ0.�d�T�R�.����R�F�!��b!�*��VF��!ǟ��ͱ��lߋ�ץ�R~nU"Sbv+�h*`�B��T�i�hy.[R��6FvLC��L�����C3}��Ε�J�Z*.Ԍ���!�'7�0��ȱ'NAv    IDATê�NM���5/y��	��f���C�#"�'�2�8G8���N�ۺ�t
��2�E4���������>�$ȔE���Rh���#����Bf�O�s��=s3 �@0ě6���4����	���F�Țz���?G��Q,A'o����#*��A�b6r�Ap3���bͲR"�b�����	�*�~Q�;Ƨ�D7Y�`����T���:"�q�|���u�n�\v	Cf�9P��p���7bf��,5�]NUq��V�+W�bR4aLG�y��Q%��LXF���������.{o~�kp������O�5��.I���ǰf�Z|�����#�yb!�ɩEl�|>&&cXJ���׍ޞ6�ݳ�~�[1p�������o���x��ߌ��A446��� ��/�T���aqȹnl�Vp߻�x�����l�w����ݛ�J���k����8��~|��_����>�ox=~���p�������a�]���sU�&g値�(���,Y�� c�6��2`�Fa,�J�(^e	�J��&��ιr�U�������=���Cţ���������{��� 2!�B���V��ʮ��_�U���%��EU%llM���$*:�J�x�E���$��Lj6���iiNa�	(�B<��_U�R�8�Ľ�����6!�V{��9J_0%��W�2���z��Z�.�Ka|O�9��t�k .@ѿ�s���j�����{~]��"�/Lnʥ��S!�;g������gt�deX����W�j�B�2�e�Z�|_�����%�WI�(�e�D�k:��̍?����ao��H��:v­���;��z��C��E�J�o0��v��(��.$"���	�f8�g�`%�d4���d+Q�3���E�T̞���j�|��8�E�oGI۪�cX��h��,"`Vq�[N�W_�bjaO��t�+3ւ/~�>l�a�Ls���mZ�S���*�*Ua����Z�X."��	s�}H2Һ����z�{��e͝�T�8a�:!4�!�ٹ��(�y�i�L�a�nb�R@��A�DK;ښXݿ�ЇaR�2aR��k�;߿����+����3:���n�;�p��S��
�6�ek���ţ?��,���λ���y�޷G�DZ��6��2,�-� N>m#2��y����.���1JsXum�����F��ݎx��|ᜅ`ن�/K�U5�e/��9�@�¦���(�����F[_�t�$!�;k�PSp2���-��U뉇�KT���\t >���c�b0ҥv}�3�P\��A��rM�ϡ��e]�>�j��9A���j�G������ �T��&-<������0�������:9=!m���Z.�R�c���BQ<�����G�&D8U.�C����\6 v�DrtMD�
�tE�`���芟L�9�0E�Uc�b��!����M��Y��y)��)AA3�˼'�[�F�0��#����6�p���@�w�ὕH�+�2A�,מ�c[�Y��s(�U����'��������s�1�~��T��B��pa�}R	�D���[�E�nA���:4!mT�/&��j�%��j�:v5������}J��^��P�}}80>5����$."G�0/�����c�����W¬�g�|�s���]��g$%0�7�fgq�I'��_�fg�0,O�0�t���+d
��q�%��k��m���pt?���G�@���)�y�f���?G6�*#4����04tP@ص�^�ɉ	������E���A�����!�ڇ·�����2��ͣ���x��ٟ�[�3暥(<�	����J�A�Z���n��192�x4ҫV����?V�T���ō��NY<��
�y������^������L�`P
C�����#���'m���'<��D`�?�ͧ�N\tʯ�aZ~������ӭM]��^ԕ4� V�I�g�����	�%ܛz��?�{C�m���)��[���7��g��1@s��k%>�mM$i���S_��
�V������l��r<O�ϧ�����Q$*�۶�ч�o��O5g�ה-y۬����A���/���
%U"�|�/d�1X��yP��sE:h��T�~�M�ʯU둜0��3�~	�A�[������L�+%\z�F��ꋑ�A����N �B �/|�~<��ҁ�mSl?�%a�9D
���:���q
�U�t9G������E�\A!�G�/_�B3|�	5#;1����7����Dq~bd��8&�"��ߍ��	�BA45����#�,��߶�N���C"����)�d����H����޶�LI҅�m�p�����	�+Q�Majd��ø�m"�O��Ɓ�;���lw��B���[�؄L>��}w��G����;�I�
ư
�Fz[нl >^�L��9x
U��T�f��v�=t�@Q�F�	���}ۇU�Ň.�-��3���^�@kp%_��)�4�������ԀC8�diw^�m.�ɱ��?klG��M��əiߊW�)*5�Ç�!U�կ�ϭ��V�J�d�� ^n��$g�P߬�M��7Ǣx��W#/��٩i|�[wbێWh���{�2,?vF)�aA$*2#�r�N�]��y!�$����e��T 9�ʠ�۾:x�-���uu��/L>Ee`�֓`ښ� ��p1�s�xx�{Ԛ� L�y9����r�
�tZ����"!9�*墬_�Di_��
]��lrN�4}ݝJ��\ҍ�0��1��!kC0��;�g���Ʈ�L�����E����(�gE,z~�vPqT�T��Dك�����ڰwd-��ț�k�b>+�u�	r�:�3(e��77�H ��<��}��v��M����+�׭�l�6'�b�&L��cv:�X�%���:��P*��[���tv��*��$n��flذ�̼��B��?��p��f(!�k�v�j�����W��N8�rY\�����'?�H$!�d�G��Sa�c�[�r��(�+r�}�I��-���.�2�ϡ��\�����\:�X$�V�B������R����&zu~%����Pk��a<���M���x��[r��(�h��p�A �A���Me\�{E����Ndb���8�ר��1al�i��HMQk ���+n��r��Ɗ�j�*��~}�X���x���(�����1�w�E���!ܫ:Icȕ����>������P(���������{���ჿ��Rͷ���B�b�I�.#�R�IT�)��������kJ%�2-5�'��z�JgЊ�%Ƴ�B�,F��5is3Q!�� :f]mM�uD��<�,����Cnv�zA�N��?�b(�[�{?��9�)ۃW9��5�vPBb��ũ#�G6z�9�����0�b�d�a��v�{	;�5�":�Q\yօ���V��_���N��:�wҳ��ݸu� ^=��lF���@��,Cw�	���cV�Ʈ�_��2�Ju�\��X3��axf�kW��G^7������߂+ϼ ���C{�I;��k��\f3�ڋ����i�M F��Yg�/#�O<�k|�k_���n��oUE��ӠY���/�(�I2QIqɱ,e>1�fJ��r���!�|&T��n΅C����5���Ց �A#
�,<����*�(y�'�x��XGڍ�t���_��#5��ʢm��&��^�E���*�-
M��v$���
��Vn�geQ�X��]�b�S���ɖ��ފW���+.����G�I*���Ǽ�K_�/~U�97пn�lX���Q�����0O�B��J�� L'U�5K�q�;ν��} �{�,��?ݮ���z� Y�ZE��y�)®�jr��rV��>t�?�d��"��g�uП������w8��܄v�d*ˁI;4^�����L��ZgvfR��Z#~k����11;�������)*庨�v;_?��I���l�,�(�{�n�<i�����,�f����b|��������F�7Iu�F��rt=${!Ė��ƁW��g���̧��C9��}�� �>�K\�'נp<� {�qY����!�����m��be(�d&�ZH4S�����y��>�X���nαXHZ��^&'��!j�E�E�v2�3�K����va����i�almm���{Eg���գ�0�bK�uxh^?�{9��/�N�E ����ܬТ��X�UF*9l�A����5�X  ��n"���'*�"��3D~�㑵�yQ\_|=&��U����O�}.t���k�=V�ͫ�I��y�5�SF`-vY�ɗn�2��\1�4`��L'�����a���+�m���%�*��W'V�5���������*���hהF�G:	�s�j�����U �7�b��?�?���/�]ѕa4R��,����`x�IC_.H�n�JXZ�?���N�f�	+qU�
�z����f��I�2e�,N�Q3���"�da��K�:�_~!��q����z���Y9����+���(����*�^�OJ�lY�)pHi/�q���̓�1>3�m���M����L��
ք �/Y��>}�=���œ�>��/o��O���۰u��
yQp��CK<��W�����׶n��Ԅ�S�k��U�f���V̕r��vb�	Ă�X-I��!��	��^�+κ����}0�;b���_�h,���a�L�#g%�����̴+8}�YBh�=�'?�)9��Nd�a��%p<�䷱��S0SH!�L#@�=Y��d!`��Z�.�H�~�����ͫ����5V��-����e�����4����AG�������b Z���?�Si⹬چj���$�����K��D\E�%'�PA�������I���Q�X�0���?����U�ScB��q���o�}�����#�� �s3*�����/}=�(ܱҰ��uX���c��.��~�g�Ƀ�7�#�J�c�D���:��+�o��u0�P���J�.�?���u�W(K�y��9������ziK=u��䵋��V�lc�0��1��mM<B(@��~g̽c�i���e5�0O��R!��CG$�ӏ_���
�.��&����g?����;;�`b|�bf��{7�5���c5�E2��l�X�p4I�7I��{�h�@���LGrj�)��{�|,�)AX��V�÷��e�|�R�VL�M��W_������O��[�\Nb��ߎ�+�K5����ػ���T�U��UQ��V���}�~7��v�����i��b��vU�x��YY�X\�`��I1Z'Ǐk������L���
m��G�"PE���)�L~��	U8EZ���K/7�W^ۅL��T:+S��uXU��3hk���S���"��C�I���Y2l�}˟s ���+W-�u�s�N�ZH%ͭ ��B����I� +8f�\��r��%gEY_&��d����±��v���|�Z�����u��2��:��O��� L����?� ��A#����k�����Ñ�z�8���-��E@�_o����A��IZ��/�����n��b�o*�"��|���?~�/Ժ�\�._	]}� �����FNiݬ�N�Y.�b`RK�VA� �ΰ�����(XsZ�lW������"���e�X��m�b���Ӧ�K�:�^~!����|�Z�*$h&����܏W��x}6���@�˅�|�8eh��#>uU�8��D1?�;��+��dUP0��Xш���:<����	ة����A�6�g�v*�{�w\���w�C�܂Cc#���^$
�ˋ\2�+/�_��atb�����ߋ/��뮻N��_��vT�^[��;n-̺��ڷ{�4�D������'��nl۲c#���p캵��������r4�\��NQ�|�x�Q�_�:��;����K$s���0<1���A֜u2f�i�e��c��k5�⸩8a����)Gӊ���Ig�:8頡۔o���4Ҝ���]lq��
	םnG6����t�K��a�)�X�bZGKs�t��&N��#a5yD&�1ǘ���>��Zi��Ƥ��$) ��I��?����qx�0b�����D#��/���_�f�$v&|�h �{| �޼Y�+A��]��U+09;#.lC��)��T�(B��>p��a����y8�G�%�I�c�p���;-F�f�����X�'�y�|c��k�C�|�����}��K��5X֟U�0��:�׭I}@���
��\�������.jVQ�%���ჰ->�h�ڸpө������������ϻ�//KV	?�V������c���~)��L��}���lizL�K�fE�]K1�LKL2����6,�)�0��o)����;�'`U��K��m��y�xӻ��}O�o��"�E#���߂�ͮ�Y�4ô�P8�\>���ۈ�n�����hD�s�GI���B�=�:q��*���I�r��B� �&�{*�A�bQy�R US���U�En�[�`�T/m��e011��ν ��~���H�(U���b���C!����;����Q�$��lD�����hk�UU�C�9�߯��|�s��g>�<��j�é�kuz�,G����Z^�x���GF��O����I+tP���N��F"?+�l�2����J����)��t�+e���V_����YM�`K�a�3�/=Q�����_�tN�uA����'ɥS������x���~���?��a�o������\��Q���S@{���f.�9�2�S������*u���R��q͢��EYtUmH�g/�lGe��R	��v�S�9x������.\H�����M��܍���X�NrU]ȑ�Ԥ@؞���M!p	# $h `�)9Z����	�/�2%W) �K	���A<��G��9<�&�f2���n�x�	��⋅��R~��Ů]{05:)Ʈ�|�a��iv>���K��o=1��Z�k7����_�*^~q����Z�w�j�%ɰ�Ȏ����Kڻq��c����$��`���!$�q(V2��t��B\�k@8�r9	ۑP�YAO_/�9�x��3x�G���iŒ��#[-��+a��$<9A7m�aښJu����:�՛r!��Pߡ�p@:�ȅ��� #U�V�<����qJ��Qo,�7�!;��mAzC�/�"�A�a\��<�s������H�0��c�/���k���� E�X��e�ADC�.Y�@����qq<�aaU����@�X�e_��.{���).��?��{~��_���noF��Uh]2�d6/��O��p�����5�?���d�N	�AB>�>D�4���!��[|V.4 ��٪���V�^�?�e(H�fk�0�V��
��v�n�� ����X1h�X8@��eIؼ^�X��k�,���phh��$��.�p��x�9g
��W�l�G>�i.]�l��D��P�D�xJ%�t՚�j��|%E����ڎ�ַ�|�*���m!�֊��>��UbXa�0F%Qa#H!gWVz��~t6Q���{�~��W���7'��Y���dۜ��m�@(&���[v.���j��3N?����pß^�b6���I��RzVt� `��-_���e��%�u��Yte��.��QU��j�Pu{����Ƥ�l����) �ˣ�o]t	^߳�_zY��m�WP�:�E���hU�n[���I�����|�)�^����i�~������a��O����I�N@�*oG(W���~�{�-듃T���SmD]�R�h�6P��e~���%ū]^���%�4�\W�5�s�P����"�k�9�4��H�p���������1���J%PW�uE�i�5&�:���hz��|�W</+a��t �����?y�K�x��i�s�nT+s��c�ۃ�9�BjM~?�1�����i�[Q�,3�p�^hCj��a���@,�i�@�?Ï�N8��v�*�Ex��c��*�Poo����#�H��(r��IϽ�20[�p¨J�BZ��    IDATNDeC�\�JH���Y	x�`�����IdFg�h�Pũ��V��:�Ŗ�/��/����j�ٜ���D�!X��0�2�$λ�\sܱ�����!9=k3��qa�-W
8�{/2SSh
E�����+:a_z����z�qQ�n�Ą�J_HNؐ�a7�q��X��p����$KͶd���X�ϣ�<b�>�m�\�RM*aiGzU����0`0�r�A�5k�<y�0�U��d��b#@z#,�a�e���)��T5�p2�����Ѽ��2���жA�kY=�(��o�.�A���ENn�`�lͬ��
�Li�r�xu������*��@�>�.`&�D*����Y����x�l��]8���Q.�Кh��%т��#����Q��jkB��H�v#GQ\�+���j��n�E59����7V�+MGW,���l�,9�y��o>gA�\N�:Y��l�'cUU+V�g�|3pNf�(�荧<�p���mܲ.Lȏh+7�k�-R��ɹ�:6k���ڴ�	166,&�.J �������/�;�yο�l8�4����\��F�	W]H��@��"�&�`6�1��W���/�ƿ��]��T�(�7u�#�ف�B&\�r=h��,��၀��˂��ý߿���o�m���ӏ��Q��Rԛ�g�.��R��m�"I�SO?�ã���n4�v��+a������x���U��������#�`�_K��t���')��8¥��@�A]������(���I�f�����vX*�9�+qkZuX�*�;f���He�T�+ި3�ki�#7�+��T��c�e���ؿ���?��#G�e֞�CN�ց`Hilq�i�����.�w29�(۫�j&\
�)P&�qN�B�6�FP�����4��k\O+/ $G7Os�t�k����	������ L߻�ϰP�:"N�v�&�/����*d���N�D8W�77�痿���X>1�F,�Y�A��ζ��0;#xۦ3�Ӕ@�$hr�`��&���v���`��qY��QM̯��%��	¨���)��z�&"��ZF��Y��*Ԯ �rE�]��w���	�Ǧ��8T����C����LG�Y�b����4�j�	LAe:�EJMW�Eu����x�RC�dML"����c>���e��	s�U�vt`~r������!PM7?�xl7��8�mMX�
%�B���1�|:� O�_ݍ�+Vb�102:�C�F��� �N�j�L���<a�׬!@�(eERI9�Hȧ}�Lj���:ٰZ��
ª0&�jp��ʠ"9����HV���M��4I�Z`��}�y��t���|fʍ�$��Ɗ'�X9z#�����4[x��J�z�R��U���ć����x�.S"E��T	�e����V	�:l3]@�*a65'|�ׅ�|a�[��?����g����	D�a���u�����]w�y �+z��D:ۑ-Ď���#Ru!D�WV����q�,�������n+H����l󈹶�TOS\j���o$�hq}��!�p�`�=�db����?'�#��ʢp_�RIi�^.��E �x��� 0��U%�@�S�|]��z�ԯ�137-	O��F�[�Oş\z!�{�-����w@��Y����%Dm�Q�B��WQ([b�cx��h`A�����?j�O*aL�:�zH�1M.��KWq�JAX���e�8=�g{Ma7�r��<���c��%Ri��g�V���C4�&Jy-)��Lep���v���DgO?����q�g��.@s<�|�U(��I�:&_��ۓt^���(@�`]��R��ao��<��?K).�R�$��G� ��+B�uQ���b�`ú�����������k&���cr�����"Uv;|�����e|��������^�z�-r�=#ʸ��V�(��5�ʘZêmO~�\Gk�g�p�v^����B�w�;z�I_c�4�Q�M�9����pʿQ?_1�A�q�}�I�$F�TxcKT�Y��k��������0��?��2i۶�����m>��k��eÓ�hI��R��"�O#��u�l��v���^̡����]C8�I�#������Q�\h�!�:$u��ة��Q.�F*��#��}��.�՚l�?��aW-����w�Ů�
v��"p#k�2�"Si,�3��3��gD��&؎4�t�r��,f3�2��GK�sSp��hŐ��~3ʖ�v͊h0mݺ]�}jB�n�Z
�1`�S��8n�Z���*{8���\�W_�>������&x�q��Y�UG���R� -�Z��D$�X$.��f����8<2����8RS3B���=׻x�Qݞ�c�@h8������*����Aϒ>�EE[�\��,<��5>��v<�!����A�,��Y� c��r}���m�`|�C;+H#��J֊�Ց���R�'_T��_Q�v�w
"�ha*�.~n	&��4Tq���R]��Ƚ�ε芨H�3-v���g�G��`��u�-p�,N21������]Ll�h��e}Τ�U�152�~��˸��Kq�i��*��hoG&�y���g���-V�g`��� �тt.�j��j��'��:z���s��d|H�oP�C(����n��<�5�(}B�����"'�I�!TiU-�^�Cڐ>��������	��|z�RY�{M�S�=�Ŕn�;��u�ϯ\|�V纑�ť�+�f������x`Q� &�'0;=&��+�;q�E�ayw;>��۰qәx��>(�Vk(s���xQ��H��"0:����aݱ+�
�mُo�A�E�`��g߲��F#���	M�.�+�A�C��&�an����ho�������O=&v;m-m"�&g.�
���o&_�G?�iC.o�`������+/����]x��®U�+��ֶ �A�]�W>(M��`�Y#�K���v�A�PE���$�R��Y=V�%��'��!���75#9�D0S:�,y8W����n�I�R�<oN�*r;$���2������=���sv���xF����I����Uu�@(�$N%���]�l	.��B��}䢍��#a""N�Ӟ���nI:��%ɁS!S�w\:����;��)�Eָ749_��I�v� |��������}��u0��)������H����n����a���?�~���/{�o5��e?���<�[l��$NZՊ�>HM"�vUQ)fQ��E���Qr�RL׋�����h.�X��Y�t�	��܍���Ϭ��grZj����L��H��=x|a��P߂���8\a�T9�&�B
R��]-&�K
�Ʃ�P4$0+1[I�4j�2�E�079-􉬚&�{�P�Օ�7}e,�-�k&Ab�F�t#��yv��ɡ1�
<��}X�a��~�i��;�D�-=}�[�T*ri3�
`G��1�O���� �l]�yx�d��E�j�Rm����zM�qb��\�&ދ�F~L�3�B~d����`���h�C9S�Q�����,�J�て�F�Jqa�\��%)��:�����`�!p�Pd�.�i����${�w˖)<;
�F�##����CiV��$� (&:��Io�S|[�3Ԑֆ��/J�ti�8��u�jR��0���SIqH�.�������C^ly]����=$�E�GM`�t\8���:�K�5{�%��=��nn�U�E�\Tk�,�bN�����p���b|tM-�x�}|�_�g�=���<B}�Xs�q"<1=#��f�o�B����*�7�{��-_�=+��jV��"�M�\�<��ZZ�d]�0A`"�����Eتr�T E	ߪ��/ۅJI��F�����u(��"V�ydH������p��ѵ�W�F��Z�Z�ݑ	=r{,Uis�
��Lp�%�����;H۷����8">���.E�c���.N=�<\z�5"I�5��罏DB����dZ�Ӭ�p����b`p�yzn��; �R].i���۰l�Z���K5�:[f~�R�E�0�!������A{GTl��^���S�� R�����ǚu�17���ب|���Fp�]�""�!�W���N:�x|�k_ƻo�S�K9X��$�`8O`�x��&�'��h r˴�����@�⣿j ���:Q���8�ʩ
� /l��I-�t�Ol���f$6q?�>IW@e�H��/��1��T\08ްzR���|p�)K��Ylo�FO�2���'P\�l	���
���O�ߦǫx����Y�3�����I�:��^w��P�l��LG�.��J��v���9�]�E�td%\�-�|���+ZG���}�9	^#�֩�������o �ˆa��@ؿ��ԕ>���5#�L���yx��|�{2ظ�W���I4�i��A1;/=� �}��R�j5�)uŃRO�� hݔPVW �Sf|(�2��H�IP'��^�f�0�ʡ��G&��{~�����2e�*��+v�j�8�)}��D$��rap���g �K�J�R�V�}��^�{��` a&�R8�ۢ�ǆ�J%�����`�����&.y���Ξn���G�.�W�!7�D,q�%�U[4]ɣ�#Ϯ*�⪂`�d�E�ǫ紽�͉M/m<��LyU���QuK�u���k��,+!4�e�	�'��Ɩm/�*v�p����ݨ����B{��w����hqڭ��O�!}|/��i�!��?��/�{���.������l���ۇ��'���jYڣ�~�8wE��=A?
�
,��H�@�\^�Oy]�Zl���� ���tr�m@�/W܊%K1;6-�'�Jb����u�D@U�D3��=���q~��J�R����>`��)��y��n���X�=�@�/�d�E��BѨ�hXH�s�O�G'�oEe*�������'�����Vn&�ǟ|�q���� ��V"�ъ�tZ�ﬢ	#]�MUo0ٺG\a����\�f�M�[-��.���y�hUBy�LNxNԻ"��v/���s33�G���U��@�˭<:���Qe����dd}��I����%gS�;e�r���]O�Qn����1!�㵧81}TYqڀ�d����H��	#�xH��97=����^����f5���GW_��������l2%�0��LHX�?8<"m�kWc.��JJ,������_��g	�[�PK{��km�a
Vj�x��L�)C(���Л��41����m�4I!�RC��؆��^�߳��@ww���d����.s��8}��­��C�&��H��1��w���8�������7��V)�Q@�\">/�2e�ն�Z|تZ���ev���������]��K)��"��
��ȩ��9����
Je�&�q_y��p����SO?.UY^?vnD�K�g��lv9H�6i5�����f�Na~���&�ݱ�qD#MX2�ZT�&g5l�ڵ��+P��(3��T¼�ǩ�{�9�*kJM_�+��;�Ts�t[��w$q`���|�L�: L�6+܋;,,�.��osěu,;�J�PIs<u�,���}Q�U��Grpm��-��x^2�ذx�`���U	��˽O^��c[����2N�lsk�����⭧��Y',��Gw�W5�Z�by5^�~9���,����h�X���9c L:aMY�H��ĝ�m4�W���B�PF�w7��_���=��6 Q��y=��5S{��#Aa��e�<��zz�����Q�&�d�;�H�F:���D ��#���&�e.?ۭ�́1߿��B�0�z�1����Z�/��������D*�2W��Qn7+4l�Zl5x���$C7)�]�!Ƭ?_D�@s�	��9����03BHML��-�(WQ�U���a��+�ig�˨ar�0�Di>��Cc8v���A��J$I����P{Gff�ؽk��UNNq0�/]�B>�o_|A�1�+ll-pʓb۶m� ����D $��UV,�.!�s���I_�	��2L!������/(��Q�y��U�����+�Ė-[��󿕑���1��Cr�h)��]�)*1�&�uA��6��kn�TTؚ�*�>x]hc��)��'��fttwȐ���y	�<����2��2�(�5��j�07=��p�\�7���k�E���*g)���k�w���܁����Z�V���9�$�U�]�[�&�?�IKi��m��eب��0�%ªy�q'a��>��ڻw?�[[��E��X��XK#�"�*qg�b�A^��O�XL��8�/���[*�yVM!���br��#�0�V�:Z�_�>[�$D�=�qQ�A4yL.��:C�C�ḺX��]A>�*F{,�&�W_|>N\����]��*�?���,]]="���`:�AKG��;�@$����������?�c����?���'D���X��]���ئ�Vi�z�j�r�ݵ�p>�!��@%�;��6,[ֆB�D4����82�y:�������-Jpl:��۷����/�)�!�X@FS�fg��܄������{E(�,��2Ma_��g�����Δ�t����Sq��sgG�[Ƴζ;��Tv\jz/_4�����|��G��-�Q\uť��G�Ça�ޝ��/~�l6�R!'�+��n� e��.T��n�Iu���a\{]�=��OL���>oX@���`�������ᕩKJ�T���8$T����ͤKO��MsjU[q�?M���H�Oz�AO36�6���k��,5���4fC �S� ��6�#�qG̉ú3&���8(G�0 a7��o*6dہ���?~l��
F|	�n;�zeǬhF��睈SVv \� ��<�[�R>���
�K���V�h��*A��jc)&���#����".Hf�l#����x	tH`�aۢRC�Y>�bk6J5�P���;-�[�u7����(U̅VZ%�e�ג*��a�3X>����2I��ʘ4EK�<n|��F+����?g�)�PSH��(�J��n��O�aO��6�r����6<6��tR|.�*��j��i�a�}���S�9�HГ���)�31L��(��h�ı���cc�y"�`�^�"73���c�{BÇ'�l[���nDb!<��\��#�avd�hBl���	��S����DB��(eB@�w�p@�a4���GSK3֯_�����>��u�d�o���T�D���8{$�z�-T��S5�DOkN;�4��}p?~��YcQ����-��ݥ����΀�f�Zlܸ�s�8p`������Y�:a`��ސ��
\j��_�b� |�o�*��:$�*+
窀�j%+�o�M��҆d�'gg���f@P861&� �?4ڥJ;9B��2��]EmnRY��Z�v�i�����5@Q�bzb�d����׷���(���F�U��yݯ���w��=�$Ĕ���T�V�����Ҋ��a�߻_*`R-�f\�+�2�x�ч�ͲqxtD*2aX*���!
�\Jwg���=A15����$^��`K� ���G�lX�]��*���R�v��"��b1��`�Ф�:A���C��7�	��AKk+���I�F�]͂נ����|]�EzY�ݝH�Lc�kۑ�{��q�o?�>tP�}h/���m=��U�Q2}:VA�3y��m]]h��B(�͖�ۋ'{w�� �ވ�:8�Ű��s121)z~l_vv��g�F�?�`( �,�<����o���S�%4ǃ����ʗo���8�.]&+&3�!���ˤ�����;�FKs�p��e����/�3.��\w�U��X)R�۔�+��VU�g���Ρ���t��� l1iq*.7K�%Kxm���Q����(B�U��l�3�q0�{ԧ��E���M��g?-ٴ�{�'p��~���z�Z#��ms~6N�KUU󭜩[m�M�mF��%=k}^�NL���
�E���X�W�ĵ�^�x���9�j*�{^�#uҨ@5Դ�L����-HZ8P/�v�n��=Z���Ўt*\�1���@Ob�    IDAT�0�,1�[���.�6�0%4�~�Q*aa?��������]̓$�z(VkN��U��U��������Z�+�!H�dY��@,�*-�85���D�MyJjХʜ
q�aF�����i}$U�`+��I��
�w�ys�������V����ᑗ�a�lc�T�eU))�#��deQ�`h�� �xv�;r*=)�,��:s��J�2\Dl1(�>�\�"��|�\Q�
z���L��)�BToM�a����V4��v�t�R�jy�����`'�r2����I��Yz�pb��*_)�*d�X�U�b��ϦQ.�����3�S2�C [)�h�5��-b������Xٳ��+	���N�t&Ʀ�1<��#$���b(dMD�a���R�dRbl�hn��l
�㓢H��(<���R�=��Ԍ�.��|CCC�g٬�T)J�U�9=>��!�a��������썛䀛J&Q��sh��Y���DP�*�qVH�#��=r8��M8����H�U0�42��I�䷰�)EG��ؐ���6�9TC�[��5[�H��S��,�zq*SU��^�2[�cWWV�Z!������̟/�Bak��Jӥ���H��u���c]�R|}7b�:[[�Q�f��҆��<��_�g���C�9XA� [W�wă:'�8�P��S��e9<Aj`� ��WV�8�eM�m����\Œ���go�F�EK�4l'(���I���6E5ɹY�� (@׿q"�����r�)l�e,�Y��;�#��XU9f�3�C��5�/bݺu�2��c�Y���A<���x����{$9�d3[�?�ȁ���b��E��)��F"Ajz��q��h�]��3�܂K��O�\v����&�m7"�f�]>���q�bMR}ljnE�r1�(�S����
�����V݈&�r��g2�x�&�^<0<$�[�P�V<iQE�^V�sS�e����@&ǧ��ӁC`ߞ�xm�+X�fN>�d��޳O�kY͡����8��gؽ�T���{�D�_��q����ށR��.�z�T�ru�hȵt:U1��ؗ���)(4=�'�͘�JXP� �R?x6��**e��>(iĸ�`���%�ߨ�M��_�W<���x���b�ݘ��=O �$��V"qr�	ܠ�.->Gӎ�א ��J%, o�ӽ��Ue�]w��������aq7a��B�
�9"��T.�z�{�/�
z�Es��`��@{�ʰ���-V�[4��rڡ�8�AlU�y'�)Qꤶ�C�آ|#2����ߋ�l��m3���Fm;��>}�O��򙂫���ǨSuǮJ���{�:'.o��8��a�c[�(�e�ځ��9�ju͊x�X0����.⦞����|���1
��%�EOɖ�)�����Ŋ��<�y�����-�0�/b�v!os�{e���_���abB�3$�&i� }Ɋ%H�fE*�X��!��"��"�����
����L��(�yǰ�,��Ȳ�azL��9��T�E��#� ���oY/�1���mڨ�k8���<؅�rs����s��%i=3���ǥ�W��D�Sw�jU@L,F!�U�� ���U^n�yٟ��.C-_������m<�<�ԣxu�Kp{���ҋ��VʑG�W�(с��KB,G(D�����	�e�@�6%���XX�''�D;���=�kʠɀ���o	�=�/Aݍ��ZZ���6���,<���}>M� ֔�`f�l��`�����3X�g��(�<X�v.��mصw�h �'��I'��D�"��ԡ㽗�]x���rbQ'r�T�N|V��z/ٴ��p"W�����?���TjEtw*��5s���a��ۅ���	�-Y�!Oi�P�$��8����<��3r_N8��ś`T��hj���Q�:�T��g���|�1��"�~L_�z�as��SVC�I;O���r��i��r����E�Pۡ���.��m/o 6rX�I�<�5S 8�6�f�3#��3�gպj��s�-��mUQ3ͅ	9}4v8H�f��?ЋP8���^C�,�㏓)�CTN�0�t ��@�Z��c՝}"�ޫ#eC�X�}����Gy>�0��P�r*.�t� ͊Y�o6?/�K�}H%8��Ӱ|��]���r�	�Yc|����C�zw|���1����x�Q�1kH�4czj�����\r1~�󟋫�Y{S��1��g?F4��k�J-G�"I'�V��
F���I��|���/n���C�X"C,���\s�e���!��C��5Ð�۸��@�vDYt��o�f�� ,y�a�C���\?V��K��ii�SS���eFT�mY&������������8~�_wcxxXT���ZwZRC(�Z����1�PH*撔3����sֱ��"�F[H:A=�]����E"�N�xH��6���A~�9������I"+\��J�q&'��'�)�
u�5�A?Gl�"�`��$��O lA�bQ�`l�~��7��^yS��	�������ӧ��CM}T���ix�Y�2+s�z�_�
;3��m�mY���D0���kw~W̧��\��d���ʄ��� �N�x�ɦT�B�s{$Kd[��a¸�hu���R�?���L�����c*�C��EŭY	�c=�ƉE�.b;HMz�;NnAS����*$��Q.�-◪՝}"Q���h�"�
+�'�V�t*^���e�止X-�f/�f�f�����	=��H��b6=����E ��a`�,_�
��_�$M��Of�&g����Qs4.&�H�Y��2�ժ����<1Xo0�&��%Xy����߾�������UL(����c���Vb�������G.ˤ��E$S�BXP#�³�#�̫��b�ű|ʓ1 sp# �7 d��h�"���J�LX�! �٥��*������T��<��o ���L����.�u��x��e��m��F���c�-j��t��I'��뮿/���:����g�t��ƩK-5pB�U5p��SL,Tێ�0	�ҊW��Җ$�p������	�xK���t��a��e"r��Aѝ����FД�g��Gn��\�J��V���ذd��s�V�\!�ˊ����%8v=~��)�-kCSc�������4d��Ynx(ʪ+��l�8r"��#p"w�F�l����ZD��9�%o��dO?�z�����D��k�dy����m^Wːֿ$i,F��US�ͅj'|>�>��9��o�@{k��螾n���M�bjnZ����8�����*ԃ|� f<����1⹺h0�*$N0�̌M =9�& K[:�7w{�N&k	�Xr[S�����`���IJ�~ETݢ��=�)l��)����h�[��yr���e���E����wH��^����p2��w�qH���M�]w|U�ZE��R@�ͤ�.�n� y9�\��*%eʒ��=��䵦&�����-1N�s���?��}��!Ϗk���`��
��q����b���PG�~-@0G��	�Z4�g>�8u��( LIV�	²r�D"Ơʼ�ZЕ��w��7�+��%ڏ��v�?�Q��k1i�q���m*��]�-Hm�߬@�L�U3&�zS���	A����1�ߋ��;�K�J͂�c*a��DmG�}́ݶ� �`J(�J���i��AX�t��#M�V#7�R���O[ bGW�+��}�y����l�R����h	
�)k|ncU���`�w3�%c�����#	����������~�`'z�
]-L�eM��M�s�����6#7yq�!ܤRل'ǁ�	|���C���g����Ǒ�(��K�\�^�u-"�E���<�V�.�ټL�P� *R�h�Z%�h*��prŒLU�!)�.[j�S�G��xG�� �ш(>�IV��/�c�Q.V����-N�q�pb����ORm��2��9�!"f�@�Lc:9%���N�<Y@�DOO�����-�1=���ĴT���>nz�� F~��DWD�Z,c��\��5\X�l�|�Ww�@.����/��3ss�#\�Oc����]��G>�w]y��LD�n���+[�ò彘MN��&��{��/'E[��R;3S�|���hi�#�/brja�|>0�$ɗ�D�Pd��4�ja����<9>!�zj�����0|���xn�K�dM�v��{p	j�-=�8�����O��2F禥ZutA�Ζ5!��Šv'�.���163%����Tl<�K�0�c��&�A�J��VrD��� Xۢ��¶���.�ZU1o�ArgW�\�@(�=��addD�Cvub��5�W�Hr2������-`d�~tŚ�a�r���O>���U�kr�n~�	\|�0}��ͯ�eY�x'kE��E=%�]��V��\A�2�lT(�B">���F��k:P��ka;��7�O�d:�*VQ�K���O�Yg��R��{�>a��\��eKh�ݻW�y9lhI�(y	�>����G�a�g!:;U����R��T�z�
@`<=;�=�v��{�G@�trF@�$�.hV��5Iz��"�쐧]�^w ��$�F���p��a�sx�ʈ��(�L�]},����i��F8ԌH �'�X�	�\^�{)��j�l2�@���-_SyJ���DbC IE�� �oGg�V�N^�O��!t�5�,P�D���K�28�pR�؏�%�r��T��aDcM���EWG��g�Ie����p���۾�m�^�����Ȫ����]Z
���ab`-�FM�q7�{�D��cr��jL`��(�n��,�&�泎�6+a�����2٦�J�s��_�	/<��򡟡�ϊ;�c��RAr&c5��A��# d^�T�JJ<���"Tʊ�W�H�ӕ�W�-o9�}=�mCV���@U��Ry<pز���٩A��l�'��T��XF����bi�EB���rڟ�ĩǢ�}c��h��H�_�*��5��J�Sq��v���X�{# �^P�0�o*6e������w=�������}l	��Sȥ�a�I��n�j#NX�O)����+5�������/�H/���HuD/$=m�M��.�b�UU�j�X����HK����n��#�U�b�EM+�nHDf5�C��O��#σ��b	��4�=E��]��dHz�u�u ]�%��Z��k�w"��G��/���#za�p}=�Ԓs�B0onn@�qx�E�c ���R�y�YD�aD}Q9`����v��OՂd��^ۥ ,Myit���?\���_t!(]��+�������K�ijG{�V��%K��{bzR�*D�)9��l���_�������.�&�p�9�������UxY�)��7����O�-O��He���7��rI��v�3��K��d��R�_s.�A��̢�O�(g�z�%��@�}w��H�#�jJQ��������.�?��'x�͸�7b���163#��G�~�_|FЏC��21I �ɴ�}}r�ħ�0��@�#A H~��h��u�+ز}�V���&�u��S���5%�v��L�j�k&Br�W��Ctv�X�$㗀���ъ�e�2�Jk�L��{z�d�r��e�EXn
����B)����a��A��x��뤒vƹgb���h���SOcx|�H��������a��u��suW�&gf�AeT�$EEeDĀ�����b�u�uw�WY#(P2��<��<�s��]9���{�ٽ����?����{����y����wB����f�F&�A�4�$���[����V��k;Q0�P4��&�g�Ȣ���P�HY�Yk�될5K�Z7 Y��kp�EcfrZ~�xbY��\� R�v��G�_��0(�I�sYB�-W}�:!����*~����"��*����hfq��(��'��_�6�]bO����o��*�4EBO%s�ɳ�3,�1��(P��fqbvj�8,��Z�X2�p��VA�ՙ���׆��	d�%�}-��20[C1�N)�X�jE~Q 3xR,�U���?N�
���X������eGR��K�A'�\�u���Q���zY/��F����W�?��K�eȬq�5�Q1�"X�u���v���A&Gx��CQ������'��(���AN����U��fw�R�c)���R�Ź�p�T)�\@@��g���^{A�:���f�My8����8���&<IG*+��]Y�T.���&E����
K-lV��X<.��4�}dD!.���V���IQ�4�(�}��B�L[']6��A��`ԅ
�NI'��Q��z@�@�-�Cj-��x*����0���1�g)���f��V�pH��(ʟ��/E�u����<�̮;a
�E+P���4�-k=�d�p�gcS��J
�zI�"�0�ŉ�|�wC�a0YD��$Q��\�1(vm�āF���b.�%��bJ�{����Q�A ���#3崢�ie\"z��Z�4�����B�jl����n Af�����!� ��> ��3��8ٴ�4��E
DË���\е�T�������P7kQ���ce��:�1jk6�Eߺ^�F0:6�|��D<!�+�pyS-F�<�P��ُ`{+��	�9]����َ�p'�v��y*�Kx��GD�E���
�Z��Z��k6`bd�\��J|��kd�`ҙ�KD��?���Ż/>_��=�]�bv#]�Dn�:�_:V�ň�\��Y�����I�k#1%��]t
�5id�����BW��j3"W̋�<�L�O>���غ��˿ߍ�p�s�025-��ÃGqx�����2��PXN��J�億�zc�D?�*(�AO_� [��]N\��+�k�^I��Cd~��\�X��K׈���5�f^��+"5̒�LO�na��)$S:�j�҇��NX�ѨM����Cao��>,�3�5B�X�
��2Ƨ`���\EWG'BMM���m�m~ad
��4t0(�i���cȍX9��0h�Ф���G:A,_��G�wl�E��nh��p|Y�Y�����R�^�"f��a���:z��p��g��2;?���q8��
��&:'��e�Fȭ0)�Y#���H��T#?��3��R>���n��ט�bB*��`\�/��σJ�L��RN�?�[�etEEu1)h�U�,64{��YF���cnz��Ӱ��pLȧ2�S�4�$�֤�C���܎�B�ndR�m��RӢT�)����i�l'�Ĕ<2pį��x�r'�'�a�T������+���K�l(er�٭�U���/_N��*^�Sو��q�8E�FuZ����Gx���倔ɦ�r����E���*���`�q��}�0^��j|�	%�Z�v�d���t{�>��x(g.�$�s�PW��7�L�l�t�2��i3%oΠ���`���&��O�a3!�I��uUiD���{�����>� `'�y�z�`vR@y�:��$c_z�%�tr�P$�9��HM$���ک+9�4�jz��:��.���V��W� `|.�%�_����T�'�����Y��5�4����}0��a�����7o/i=-B��#��sX�a�67��\�0a��2�u�֙%6��1bt.�o���05���|�:�.�櫞��t��F������Div�	���H��J"�	�ŀK^h��n�N�>-�tBi��4����$E[�.7>Ybt5;V�N�-!ĲI�TɄ�=���	���m�h�@kskz{��ֆ�o���Ѐ,�d7��4�	R��?1� 8W�Cg�H5�����L��D[��{��XN������#��<�Q����O�f��j	����n�q8z� �Z"��m=w~�6�-�:��&p������`��84ԏD)�U�עw�jD���5�q������ې�(��C.��'���2�8�T�pÇ�&��D`6+cf�ز3N6O����
h戢x��PT�?YF.�'ۦYd̤y� �y�<W�ZO���7�b)��%�^����0�����b|Y�.c�%�y�0v܃��qa��sZl��jkH�G    IDATG�!�e%�Hr��9�N�F��ǄM=��3q�ygal|�3SXN$���14Y��ɊIE��\`X�%�u�Q��L�"V�cC�D���>^���9�`.ݑ=}ݰ8�������,V�Z��l
q�ժ
SZ�H�5��X�α:]���>��E	����tf���Dx]t;f�Td�����8����A~y	E�#�$~��d�dØWǡ��>�X_�l�&��%���E:�F!��^c@[�UF�̣�����{)�T6fAs%	�%c� `���6��H�U����uy�t]܂v�C^���.ɘ�-a�F��'S�4�FjF˒����F��p�Vry�n ����3�4a|t\�?�B^?r��D��=�����Q��z��B���(B�.�rz����o�~��� A�#����P'�{bU6d��O��<���%�&l?�4���ì,���ce��!^�4��J�K#]]��hV��E@@�a~�� �I�T*����Gػw��W�tB�cXȈrf��l��*�T�-#�E�)�x�Afq٪�%+d��dʽ�p�rT��J\���[�\:� �l��م,Vf���8Qy�����^�� �S�
5�$�_aT�����X�x'�014�T��f�+e�G�a�9�p�����.��&��/q���Q!��[�� �����}RU����0��'�R�&���O0]��wA�|����^� d3�lШ"T�[Y9��`vF���4��G4+[��&�����������j�pV2��hj��+A���G�<��0���h+"��&f�9|���j�S��jR�{䢤������h9u�Oh�v�����1���0@U
��RdmO��J�E�5/�I���2JFGJ��+�\ӯ\l�a�¬V�	s{]u���Tdt�^\±����]��+�_�O�p���:�&&075-���U}�57�I�)�{v�.��ZE/"�R)�I+���`�Nc��`��m� �� ��( ���~���rb��U��������\<��I���k��ہ��Gp�� �[Z�I�p��p��>�h��rY=|�Z�E�xsҵzV�DG'S�#0Wu��ŖQ��a1X��O�Ⱦ�����M���{D@�՘��\@*�.N%��܁X�Igˉ�/�2�T��?��J9*�2Z��6LF|��0e���f#��4f��Q��1�?�+7��݇06���K����N�G'����ݘY�����26v�T>��k0?5���	�H�u��`��a���p�<8���Q�E�����w���ǎ ��$�����cqX4a@��F6����):4����xE�X�ץ8�Z2�:H�
��`K]=�0�M�닏�J&lUb餀�T^	��㧗���ҝ���gG�^�������蔔�[u:��F��넶َ��ɠsQ�W�cK(����T/�����4^:xY�Y2�&֡(��
�4l�`��YU�O�GG�0=[�.��S�mś�JFG�ܘ�X�M�N�,���;)��bԑn�	�Qc.'�F�-Ʉ��anf��  ��[6Ke���\Z�npL�$��S�X�8ޣd����d�ɉ�T�����!�H�^. �qIy��a���F.�1�U�JM��rã3(��p{C(VX�mF��J-*<��i�,�Y�Ѣ1�w���:�W6�1 ��&a�e�<v��Z�r��ز~-�v+�:���UJ�2e �$�P�se��&@(Ք\;�ɵe���J� �Ê;��9ė"��T��4Q��P��EJ���vsS��j4e+l^N��{�\�#�M���;l}C��|^�4��d�5-"�$#K0�Kc�``-��:���W�y��4#pcd�b�9��2	IS���Q�,���&������6����H�|C�>'y,>;LEY����T����+.+=E�"�\���3���Py<U���S1j��	0��"NK�==э���NM��Ө	�����KD�::U0��1�5a�&�����9�sz�~��l�$`8��hN�|���_�}��g?�̫���u��Rr	.[_AGV4a�]~��0].�Y�B.#�9�݋�D���?A���(	�T:�Ș�9H�0'�r��)���޸cU��̲ ��Yq���'�$L /�.WPd~/@�Q7M����
�8����b5
������B����wF����$������������q��!\�u8e�)A�	��*|�ײ1�`�T
��K)W)B�"�Ga�M7݄pk#�Zv���=��7O9�l޼�6n�m�A"Ȁ�Wt���f��$��*��]~5kqx�~t��H=�R<*L��j���!LD�ѷv5֮ۀ��1�&��>���y)lZ��^�lc�/���.�{ޙ�(T$	ۊd�"l[e��;� +���%đ$�^�-���dn�u���=ɪHX��*`�qB4یR��8с����03>��N�o�x5�C�0�@�F�h����Q���_�n7c)��`Dtf��o������vb~zFm�����߃ǟ��^7����&�s��U��K���r3�dzjJq��H������c!u��,ɀS�jc��'��	]ɭ#�P:��������F�T������"�������\J��nҧH�?�y���T�(ZG�Q���@�����NZ(l&��jQ6T���3����M�F@�1]AH�ǹ+�`�T1�Lcx>�x����5:������$�Q��eT��Y1��.bvr�lQ��q�����aza.�Wj�8�q�H��yE�l�)�7�=��/��M��	60���L�	1f�e�t�q�/K��y�',��̴��x|n�2i�*;��T����T��c&jCE�Li����Yq��7�����=���UW���~�5+�|������Ԃ�=�,V���0I�~�"�f�6*1;��R랼n�q�F���$:bU�Yed#��G�4�*hy�]���L���>��v���@6����0�z�Y8�X-ND�q	=%�I��;-����>fs����V�N�caq�@FFF�J爛�V�=o�!a�^9J�?����K� jV��L2!c;�ˉHt����5y�d�Q@C#�Қ+2��
���8U90J�n�m��*��5 �Y���!r	�.[*L��Y����X��NN�N��S�h
 &�J%�O@ICSE���̦�֕W^)��7��%�'��X��@#S	zV&H*I��e\G�����Ca�Na��o>�=uB/}�#V~����q�� b�nM��9���i|ݸ>��bP����I�}����]i�������o�R5x�X���f�EGНң����`K��tnS�fvz�������N���y8.��ZUĖ�F�+���?Y��D��r#��vu5���H����.�>z�8���:2�
�Z=2���A;¤��q�p��D( �lab�	.���V��ia��S��>6�{�d׿烸�]a���H�㘙��>�~����Hy���}�!����6���f�N;���j:�K|��/ ��ǋ�?#�����{�EhM:��s�x�%�?���c��g+Vl^/�d���
��u�F̏L�P�ê�cdx˱(
�"
�*�^�&ѽj�hq��&1~h�}�3�����3�H����1<��/q��Β�'O¥���#JE������T#y�d}�~�k�h�ԑ
+����L+��q�S��D�q���G���ժ������%2"��o�x�]�A�}�;Q�k�!U��P0��ů�#����`	�]gD��G����9��"��( �)���6�9��G_��&0����u�&~��g����Q���� 15ٝ�I^�L解I�/`�V]@�u��N��"�ę�".��j�
<>�-͒���[X�ߗ���@3m-�d�H�0;l*���rC�h('�Ze��I�׻�(���]b؄ѦCA��B&�����(�t0뭰�u0frpT3�� `2!=��2�4P(��+�P�L�w\��ˀ=[G)��z+�&u����rI�)����XTذ���n\64�5��ue�-�YCv���ߗ�c�X�s�9�����]����2��l ]�		�,�m�ʺč�ϝ�G��/���& 1�0҆����a��݁{var��M�Z����^*u��݌���=��Q����~��ǡ3X�B�QF��a{,�N���+<�(�y�n�:��h�]a��x R�N�C�uZ�b���/�-]`�4��C����_FM��EBe��ې��'@�jԙ���;�@��������\�h�����c�a�ƍ���07���w�_��ļ�р��s��~\p�ŎW_�^Xj��n�HG�}^X�FI������#�Px����ݸ��;���pzQ��-�ϑ�r���G#��tw��^�bzzT@����<<�3Q�}#�(U�ZR�_<X��/5s|<�䣲�¢QH�p(�c�nJe*@���W_)k5tJ��_C�t<����Fƚ2�$3��7N�!���xZ=�����q�� �NUX���ԟ�};yl��{u=����Q�'F �Z�㗬�5�:�R���z$�56��F��d��!�Fsr����E@X�^w|�����=����"�El�؆��:Cu�S���gc� �,4���<r��'�V"�,�f#���fI^������О�.�0�BՈQ[���T�W�
�����\Q��F��8~��h�'��9L�/ �ͣ����Q���	�N�
�,�0a��0�f�,?M��,�]��Y5���	��x�7�c�I���] ��D:!���<���a��P!5�QY0tFm>,D����>�P��#C�<���z��X�i#V�_�{~u?fcԭF��%��a��g�H��)?5u-rKI>���/ǁ��逧-�H��w%�*����4������k��&ca�Q�5����^�z�)�v:����G>�C���F����s3i�B��fB�W�㚀��St>�\cM�0��=E�O�
�aB��Ts�L	�G�cv|v�w��?�2n��V�^�Y��.�X}6�O���M��܄T$��p"S3h�4a�ˋQ�ډ�c���1P4���f�����),W����4qMnش	C#�X�� ssb�%uO��J��F+�	�s~P[�L��u4�Ȕj2>��`���nFK[P�!�RA4M�{�d��y�>�B[L'�`�@��|�`��S�9�V��S�Rm��R7®WX�R����
[���&�����J��^g3���%�U1D�M�א�+6(���^՞9�����6Er(,$�05'Q*�V���"VWq�-d�J�7
F>Љ��W~�
C*���=)�4��k}�&�_�ܶ��X�z5v��!u:��Pjc��A2͌OX�b��40s��>����XL�
�'�Hս��E�1(2��%�ke􅃰V����|�^7�q�m_��B�T�Sr��N/R�<t:+�7����P���������<�禯P�L��i�1=P���qډ.S%���xSq��8������E��1Y�������5|��_@:d�x�M�R�(,���Ȍ�����z�E���OEGG+�����\~	�9���'?�
����4�������go�[Y#0��|�Pn��*�gj3��!��6�8��h`8�DjL�w�#n��F��98�V�|c.��
amN�E�50Y�"e�����a��0�GG{�L\@�Ť��Έ]E������U�fJ��N��mb�w�uc%��TV��"}��تNƫ4�{ww���}�<�t:)����f�l[1�9�Q��ϟ�y��/qo	j=Y�2a'�dK���za��	@vr�ncO�_Ƈ�H�{���0ѐ �_S���Z12����~���͡��6�d6�o0�W���u��~灿y���`4��"8���ڋU�&Tâ	�� ať,��e�w:�Z�i_4(�g٘"|U#��d
T��k�g5vd1nP�t�Ŗ�â`ެV��}��RN蓑8v����1Y�H$���'\j����5ad��
�H��	#�#�x2}�
�хz������n�A��<����Z���_$ ���\##x��ߣ�烞,B� +I;��E�M�[\�D���Omm��
�Ǹ�~<���HT��}х����{��c�p����@KG�Q�9X�&�V|��[P���s8�8;���Q���+ر�u�l�<u3�^e7x�w��M��y�%��E�Ke�)$q��V��ƹ�	�ۃjو��"
[��ĩdd)�����WޔF�Q9!����e4�ӡXTX�b+��fE4l�a�ڔ�&m	v�SC�����ڝ�Z�'�AIk�9�_��N'z�Pg+n���X�,a!������+�}�
c��J*��� ��8p� �q��0W�Z�z��v���<<���eӦΏ�s�=W6��R�����l:�d4��bL�Ȝ�Ҕ��!�w�,�P��Z�ȑAF}����r�?��@�T�ܴ�@3�ZÈ��H�R7�J��Ⴜb�J��+k���у��X��ՙ���ds�9����غ}��<r���4&3�� Le��-:��2��"4<�S�""���~��I���� +%�Z�fti��;4���Ia�<V������)��U�)镔��R�rU"N謃��E���G�o�l�dL���⺏������G$��	S����P�~������ǌ��"q�&��2�B���2N�0]�L!��\YGU,�i��k�c]Kw��y��y|�k����%��]�����R�q�vw�azf�E�F���0�J+�D_ޱ��˨Ȋ�Ğp����K��6H�<S�El�_[\6�d����/|���J�w� ����O�_��?���ss��v��*���,��C�M�0�vbl�:;\NFFY��͟���~�������n��4����s��+��5	ye�G
��|��V������67|�e�����R��/ގk�y��4�͎��xǗa�:������@˼H�*�D��r)�����W �^����ʥ�D�Y��qв�O+�>�,��h�v�cX2���P�E�]�$$lH�%�x.V���̆ ���alY�Zb0,�2Z<h��hF��L�`��cP��R�L�ǘn2R����L��ȓ����;O����0%���񧺗���4\�V�.U���4Fq4���x,�����)���<w�=A���*6ϵ~���~��`������#�ǰzE"�ob��fd�ֿ���xt%�RKД
�f$���A��,Br��Z++ԥr�c�6�xQ�)�t�)�o�*k�h+t�ԥۍN:�H�(��d�U��L,%�g_ĳoA
NLǒ������*:��2&�A.b�S�$�Tx���u�5�I�0��;���p�U���m*U��Q\z�Ű�JJ���C��ҫ���t�օnIe9���0o�`d�b	���gE��y~v^ʭY���̭�Gd>����^����A-�;�:�d�218���k���S��n�,J�҉����|���_���Gլ�!�Ŋ-��o�^���ٝ���p���o��"����]8��0̰Y���N�Z&�oTF�:��N�e�%w+�Q���J��0����ĕ�U�j��6:�x�(Z�F|	�XZ����a�sY[Z���/�^��)��	�Te\��$r`bb\Ƣ��[;��iF�����U<z�p@��=�ڳ�\L���ٰ
=�`22�х)L��hC�*l?�혙���䄔+s�&���ǖ�5����$�/K�%�X���B�\���Z�!,��!�I��~��<v�z�#H�����h�Oe	��*���r�<)��arrMM������߹����Qa���8�'��8�#7�s
[h���O]����t����z\�L	,��v6t1�5VYE�� I�����1Yn�Ԥ9j:��FL�=���c��:����'�v�*1P�M-�D��c(3�)��4F���    IDAT6��h���n�ĚU�����5����.�tJ2��i8<n8\Nlڰ�\=ڃa���K������F��1[��1<>&��)g�9،V������ݗ�m]�y,,��l����i�$o��ᷙ�������~����]|�+����ݍ<=:�h6	p�f�������/P�aWn D*Ý_�*��4�ADfsZ�'����EtK�Q��2NU��B���4�L������&m�r^��x-��w� �xc7��z�;��丝�ig���|ccSh	���ã�<�J5����?q��R?�y>�d!x$���^ډWw�^GÓ�3��Z��*���K�rئ#P��8P���Y�uz�v�q�=?ĚU��������9���$v�> �֌`��d�DF�`�o��b�a�T������F<ƐVF�V�����5h���/ċ/����477!�� ]����ܻ|��Z<pX�\�St��_X�W�;�]�{�9���*
�!u���R����ew
Xc%�[��N�N����Jt�ހ����l~xp�,VG�\c%[��V��%汚ҥ�2X* ��Nֶ�˕��L]��w��|�W�.[�	�jp��y�D"�@�MvO��Rb�ػ�C��I��+6��9atG��h��s�?�����~X�
��g&��TQ�N��� �.����a١��4Pȣ\�IP��f�ά�y~U2]�Ӂ��Eg�8"MF�2eT`25�q�6��� 4@˿�!I���aR���=�,$�ПuaQ�O�UVk����ۗva*��D4������Q��� L�Xt5a�A@XsWf
IѲ!Y�&Q��Y?�
����h��p��ģQ�Y��}W���3SSpX�ػ�<���V�Y�b��M젤��n1+|ꓟ����B�}ni�����~�u[7J����,>s�������D�iD���h[Ճ�G�b�P?z��]8}�)��7!����3O�=�8����P1�8�{��C�B��~I��p�D0r���d���=8�u��m���1?�B�j�
`�kJ�oD��*�Ԏp���U\WuE\�ѝ��#(N>�,'n^�'�����@�����; ������3/���v��r�f2JTFU[������ �X�n�����=�\�Q/��+�y��5~�嗰��A$�9��Ft�[�pw�cs( `��G%������8�3057��XL)�����������0�L�x饗���/c��Ű�Q;�;$�w~v�~61h�'��˸��1u_�����ʗ�����݌��)$Ri�_�~�{sS�YtQ�61��/,`���alr#�/#��	}T��(��Fٔt(����Ӫď4F�|�	�(�'�1��@YɆJd�Z�`����C���M�G�<��@X����;�.�S��>)��}<��(����'�B�?��O�����˘���k[[���<��H�K3��Q�ʵ�#�m�Nõ���;_ށ\2���1�^�V�������VS\m�Z�\^}>D�\^F�������tS�̎chjJj��A�YW��5=�����ￆ_�����]���C4�,E�/��<zV���䑈�ւ����&LN��}�f�*l9u��[x��!F�
`�(R4a�bR���<� J����,��J�y6�S���rV ��^'�[.2�p�����?�Ç�btd>��Ȃ���O�MF����RF`v֙�#�\���>�+��o�Y����!�͠���H�ǆ1::�X4)ڷl�9_ē�u`9��F��Tl2�%O�^��b��������>طk��J�?�i��Y֝ɕ�q��ڋ�@+v��#:M�l�
��;05=),X:��u�:��Q�F��*��r���h2g)�E[����z��e�EK�����@PqU��i����eY�	>yN�Zm���
9�/x�ȐE�>.�\��h
��w��#\�O� ��!3L6��h~?��Z�E}*��.�A@�C��Y;�1=M+bv���R+��W�Lj�?�]u���T�)�172�*ӧ2�$x8�8�=���R-��LIȪ��Ҟ|^~~x}M���`!L 5�"�aÃM�Oy�b���W�v,�����>��kVS����|�z[�!��]tֵ�`�.á� �
ԎPlo5�hk�Z%�U�CC�øfs�q�����L%_���2e3`�s�%��k�vwjo��G�����tc`��I�{>��D㱔�DO��F�i�FO�[A�Pg���R�3A|l��0J�����8}�Va�F���»��a3��
�193�_=p?�^��pԚ�Qx*)�Z�J}��n6c~1*�������O�@{~�B�u���G?��g��hoFSW<�f�:�gڜM�	v���\�Ɂakt|�Q�k�k����_B�u�ⷣs�Z�,��!��m�ʉK2�*����em�>c�,,.sX@j6E*����ť�Ut�R�5Q`N�"c��i�7��6[��M��F�K�Ol���V�0?* �^� �چ�=�^8py�i�h������Py49܍�z��l�9h�4�CW�:��iijx^z������*�r�s�J�CM�LK�uEW�edh��7�y�F)�N
X��%�/Њ��p3�QT��]���z���tV�f�m;n���S����������-�Cby.���mD|�	I�#��l�$	�&��t	=]+���08<�\���{w�\�֨�p��]ݸ�������~�ԝd-ut��
�:2aea<,�K�a�/V�h8�kFȟ(�U2���"���si9�v�Gw�A%W��j�ٛO�./^�Ë8��X�4�����V*Y,���blfF�s�^�b!�ˍo}����O������+c�&��^�����҅����xw��q�;ލu�+�ㅗ09:	�ծ���&a������r��2�lר��>�b:���a���T8L.�xX)���O�@�!ąm�Q�ݮ��f�ע�O�������ى���/���߆��r�j	�]�hn
���!�ESs+ҙ�$V�[�����߾�;�P��^#{��2�kh䎳jc�i%"E55�P-f�[^�m�����Z�̌�Rtq�C#x�wO���a�����L���RVX�xlc�3hnj�AoFw�J<����tt��g����.ގo�[��8.���k�/���YP(�N�<ަ���
����cn~:�82�N��ݘ��$@��dE"5���I\|�v��e#ҙe���K�T��-�E(؁@�]F�d�����+U�}^�N���3�f��|�J�B�Q��ǡ>Yy}��4ܐ�s�"	�����#��V�I�s�x�حv訛�#�\��Z�E�͝Lb����R}��O6���1'����\���'__ey�3�`���[�&�TR\�Z�<�9�L�R���#�J˸]��������:�ol������硂6F�`�$B��bQ���f�=0��5���$@��??�����$�N٬��g�Dv0�N����5'
3��JF��o~��r�bq21�������00U����?����nq�{�Ȣ$����Tq��f��x�i�p�e����^�X�\e�������b����Kjh�W��j>�V.N��2��F�(N%O\���=�:�ՐӔ�di��+�2��π�d&�X��Ə��P^��8{	�2����4��6~�:8��	�le�!�h�t�E�KbqN��1~�ݾd��ٛ?��\s��v>�_#]�e�]��kנZ*�n���(�y�i��^	ݓQ�VI�gOO������r����t���ď��)Z{;�h��.�W_���y'f1,����6�<.���`��v/��X�ڋ[��8��Fa��=-4&^۷�����U�Z��Ug�w�'L���0P�Ek��'��:�Fl^݁�N�  �n`fj�:O獞2��LӦp;�P�dztZ�����XN��EC?�;J��Q��ݔ�Z�Rl�6�@�+X�L`t�P�"�։���K��D��GI���bD� �uy8�FY���
z��kn���N����${�ı9Q�������
s�Ѻv�-~L'�i�J���<s�Z���E���s��H�F�m�Z����+V`�Xa����������?-�q��9��m��7�x-��؝����|M�Չ\
��)�ު^�"h��ӄz� �݉�hTF��|�7Ҋ`0sD�3�٧�%�2s�~��/Q�$�k�jĐG�V@Q_�Q� `���9V�L'��Eh�((o�[ۄ9�g�8r�l�n��0uhH@�Ck�y[��E�?��O�E]X���8��+5S�����Xx��u���ÀڎN���Ɓ=��K%e��v�K@�q�v`�1�@ �fn��f4�<x��020�&�O/j���&8�n��I�Z�c�ZH�!��cزjj�<\f;�	1_8����3LE���O�Ľ��T`3��p��w}�����؇�?u�V��+���u��H>� [�V���|	�h}+נo�*,Dcشi*�"y�i<��a�j����H���]e#3J��qt�2��&"gLI���S�ο܅��ފ��!�,���3��~��>����##�Jb��;0����+V#��"������~lذI2�`�I\u�eX��?�鏅e�v�{��}���C�H,��T�7XQ,(�i����"4ڊ$�� ���	~O��att5#_L`|d ��|\��w{���q��Q�)	�w�h&��P��f�+f,ɒ+��֌ޮ0�g���B��;���|n�C�䙹na�ʵ�^<tjj��N���,{�f@$�Zت�DU8�nm*�VN�)�0�.s�	[j5,'��Y:C	�Xr9�,�[��{l��H���0�* ��k*A�"a�L���|�f�2f�;�e���^��]�9��5�����5�`�ω�#�R���ߪV����7���b��A�E&�q�ٌ��(�	7K��-����E>�����w�C7[��A�&���#�����s�f2���{�c�?���@3����<��:6�����A_�7\s����-��I!�MI��J����ٴ�l���a*ݩn��*�\�t:}��\��5U��:,�2ja�F9���ș̙�`@�n�b�������0O�օ �N1E���lX�ž¨	�H����bVjHFgѿ� V��PIq���ť^�7v�!�+��\H��D�2�g8����� )�rAR������J�3ض���$iL�����è�(P��ނO�|�Z��u�Z��нa��'0�rfp���&�l���n��c��LȤSH�x�������FĥGۆUp��Io�jިL�z<p�S<�M}m8�2���1;��Jf�ܼ���c2K��g�y?]]\@��^���M��������'g"�jB��}�%ˬ7m��$F���^H�9܂��0�����pX�%�mРbb%����#X�_�MkA��	��ڀ[��	#c���N�3s���?~�t����遣+�E���!l��F�uDƧ��-Iiz�9��+Wc��UH��`.j�w�4����Epl�_�z\��GmO�^�)+�b�ΗP�򔮈�5�G�ɈiD���X��P;i7ۊ����]�����L��h2�7�3��	��&a�.�KFw4 ��W?CN[C�cBǖՈ�3�	+5�6�~�v����Q\S�yP5Y��A{_w��8�#���B��I�xm�f��a��0®&���ԷN�׽��h	���?��/��\6�P��hp��`��~�Z�\NL����ӋFldtM����\��#C�{\
ˮՠ5Ԋ=+��b��=����PU�幜09lX�y=�����Ò9`lU�����ͧ¦5"[B2��Mf`x �y��?����%�G�1ข��a|����̣������ddƮ�P��<��M�x��w��mơ�ǐ͕����߇��a͌���/��=��h�I���{ACS�`���!�D�-���Ț#v�-Flz-���W����=s3\V
̋�d�صg�K	@gg'��r��������	�5��ҩƐ˖E`n	@��`�u���~���aj�<�l���/~���aLO�#�#2��g-����TE�&�������	�5���p���3Ȅ��mf��p�֍x���uv�������g�-T09���R�	etF��j�ybz�d��KX���>'R�&Ƈ�|���+�(eﴻ`����,C�� lͪ��}��q����!�Dώ���5�Q�+��C��}��g�z�h�j�K^�`�YI�@�,�c/Ƣ�u�����\<q����z��K�Ep��#��A����dF�@��.�}�9�nk4������ĵ�{�?�Ϗ�ɿ�9_M�q�n��S�E�/7�|�4g�ת�h�׎�P|�%5+a��U9���lҭ�r�j���]���CLSUL���x��z��oݔ�8�:s��p;�pز��cX���uW_�&�,!�s�d�����ШFI�ڀ���|��LInV [���-�K��!S/�es �[���Z6�6<BU�0<��*���?�`͈�xB�B�yM��j�d#�l8IM��I��0R�.�Ka�,��"�s9<�6����:��"�r�&��L�՗_�o�Q/�h�~��D����j����1�!Y�w��-���BC@�+,71O��pXN�L�_,$�z�&����ciz~�!���{���oFd|����YLxm�����5�<V�8}#B]�@TS9�I?��ܖd�s��ga���ӂs�ޤ�3���KC��KɸضiI6٠�34��^4�8��E󥜐ؘ����ο�Oa��SW�vj_DA��"����!�ri4�[q��O㕣�(����I�[Q��P�c^�ѢW���$r���~����ҳ����052�J�"�s�����p���-
�醽+���	�}��=�穩Ԑ�-cin�BYFe��:�����܁�|�~�z��.T+93���:���+lG6n��������V�ۉ٩!�'��V(�Z7A�85�j��ȧ�%lܴ�P���py��'���/aǮ�qx������nݶ�֬�Ų)����[��ֳX��Ӱ��(��g$��8�AH�y�j����Ըe%X�Rm�ք�2p�F�C#�C���}GPJ�m�F��X��}�~ƹfө"Ѩ8�����w�)��j���2��l۸-� Vu��;�����(F&&141�|�*���Bn����hq������RK�05:�v�����[�F�����ގwm7~��#hom���<j�
�4�����c����@�aj5ɤ���a���p�q�Ǯ���y�whk[�/$�.�#���l��P��i�V���"�x��g�?�ji���?���n7�z��~���q�{�13@�dH�Q2`�0�%��[5���]��<>�����-Ls��:t�P/���'twwc���0?3+l��LMP�`xh.g2�,�{���8p���������w����8\u�{�`p�?�˯�j���O��|��Z��!P�-C�TP�u�8������N���-p�Lx���ƺU�0��t�v������c�2����Z"q1J�D>���&�H���R1�hdf�I�^�eRA��T�mA9�PrB������?���j4�.���h�3�H�	��k�LB ��~@ 7:1.�$G�lq SD�?�cs���H,�C^ Є�A��-��ľ}{���'z+�_	in����E�+��V7��6�ٹi%\U��Mp{��2^���tN����8ep����[�Qms��ɉiia���m1���b��U��]��jpn	"]R:y	��Z��~,Fd��V� 3���t0s���i��a���:������Y�F��s���q��]�z��/�v`��%�����jm	G.g	��ZV]��q�&4��I���*%C?�=��i���C!忍>,~�QǓ��:��N����n�20ԁS7���e��t���PnC���b�����~T��&FW9��    IDAT�$��歀B�hTFF�j�զtG�e�
��b|pT�X(�b%�T����t�)2�EriI@X(�$�?7��`8,�dR��8�Å7��ܼP�|��Y H����)��t"���^��'�`o�6�֬D�=��#���ScD��W������旖%^Ho1�&��J�X�h_ۇS�=KD��TFn�R�,�}�ˁw���c����y�l��T�
��9�Q���`4��IW)d�I-�+2���	_��,|tX*l��-��
 �xXz�����G+��x|B�0�	km�ݿx;�F�kCk��g���Z(��ˈdr|R ���l�[��n�ッб���3����, ��Fpm7̝��3��/�G�X��vj
ez}�8c18�&l�z.ֵu�k����?]]��T��5k����/G8�����f�V@��W_D">M�yIe1H��tNY�" ����[��\v�EFF'E�l��`�����������&�J��+��	��D��������z)�0�$iFI��qW������_ V�d0J?"�Q�V� [��
��.ḹH#���-!�i���5����	VV���57adtD@�/� =&`�.I2.���:�8k멸��K�2�?�ls&����8~��3����h�
[ɱ1��^�������rcrt]�������o�+�<rH6&�]ر+�s֭Y�7^݁-7���m�D��������x�w8:Џ2#6��պ��îCgȁ���qL� ���r����E�2˲9�]��$\�B�^|63Z#��I��Yg����><��3x���a5{�L�u��)5���o� F�;M6�Z��u�3��A��s��Z&	]���Oۄ/|�X�+"�JbϞ=��sy�p�<�NH@0��h�`v!��f�QZ�6��)^W]})���A�\�x��f���7����d����æ�0�ј�t��E,-����"R�͠`��� :�Z��D������_q!͞�5Z�cw�?�ӷ1���h<�/(�:D��U���%�=�,+ˬ�OΡ©�B�tC#ݠ���$TPd@Eg��q�A��HP�%#��Ρ:UN�N���ٟ��gw�˼���g�a]W_U}���	�~�u�{�k�t�0P� �I�.L��I'D$Ϙ:�?V�6E�gZr`��:�B
�� Z��_�+�5�.����g6��0�>�,[��a�C!a��v!�5���8�d���1������y�ɐ�Ig�R�*��]ssfffź��R��@�m�(���a�ۤʟ��J&l-mT�2a��=X�r�0������f���I�LLL
0���P�cjj--��*�gwD�~�~���۹�Z���,��/�������������l�|��-��	�9����a��3a�)��Y�Wa/�9���'�~}���+�/�Jvg���(��0+)XLet�6`fr�tR66�J���rl��ʊ0_�Յ�<X���{IQ'#��bcԪ&1�t)+���I�}:����5�A_��Z����:K���"���0�Zq0�@X�*���D_QafU���p��,�����F����#�%�2��7��=a`�O�vjƆG	�DgE����m9R����L�!K"�4�\Q*���^�B�R���x>>
��?H'3���(rCA�+��)Ќ��1DF��+:�v�
����#ƪ���r��z{+^z�%�7e,5��b�r�8��,"G+������Q��mé��	�M6;�����y8�EѰ�#��KC���pB�ۥMt�mGĈ��!�=�kdԦFu�>׍0a�_��"����PJ�v��{?�O��׿N
�q`g<S�XC0��M(B%Y�Җ��]* lv|R�dz������_�}��M6�v"����v��"��!�lZ�TT��39�yw�f<F'z}�X�ҍ��,�v� �MH����{�Bs�߼��Z���	ڏ����&<��}0��R��� P3�<9ML�����ȕ{e��\
�Ɂ={"_V�d�rL���3OaxbD�U�"$�"f'�kmkâe��w� ^x���h\ҍp%�'#mF1�?*j��,��D��&|�La�����"��t˔-}�h�k+)0Щ�hE��6�,�������d*.�Ћ�����G����T�n4x�h�x�n�*���4a�\�q�Y�H��m�b���� ���Ղ��6����W��-_�R6/�l�������7����w��T��������|�b�vv!�Є�@@��kU�����I�C�`B*�s���It\x�_ah�D�8�Ԋ{��|J�#:�[��J��6��o�qkV��� �ap�
�"Y���w❭�t5H���<��|� �ӦM�0���ð��u��
�˦��b������k��6���}�*�4�aT+�N	p�hi��3�j��XD�ՙ��k�����wݏ��8|�LR�E��/�'.�^x�9��ℓ������/���M�w�btlR�qs�U�
'�6��X[�[�Nl ^y�u(U���hmkD{�fsW\~	NٴN��R��t&�����x��o!�*#69�����v5��.������cA�e�TH#�M�P�lhv��>���^�L�٢�d֦�:;�e�v��# #�"�"-Y#�狘+��Y6�ONm�S�?>9!@�]���q��3	�&8�~hm�"��?�7kS��b���&��U���+�}�g��n�K~�ω`��{Y7>~ݦ��O�m���<�������K`Ž�����?��������xx��N���k�⩤�/|����s2��D�N�444���	�L��O:�j��r�o*;r,�}ǯ��^�>|����ͫ�1Ԕ7A1��(���2��� V�]O}g��,�8�QN�%e�J���-�u(p5i�u\t��X�PW欳,v�I�_�n��
tz�S5+q@�T	eՂHIſ�y7�aá���h�$�Hw��%��,�G�-���&H�2��(Ѩ�h9j7��M?,2U|NṐ�kg���(�R(IΜ��BQ�dg�ӑ�����!e��݃�P���|c�:8e�i1�f5�T�^�����`S'�y8�|�����(�P03=��XO>���������bߑ�tS��b*�
�h3#ch�,V47�3���E=�Be���0�Rc��UaF�2Vàb�����@S����h~O�.9J^`�� ��&!�L�Fz#I���*ߍlz�Rv�w=��>4cs�N/*�e���	�e���%���Ñ�CH���v6�#���i�6":D,��jM_���M7ӱ0�+N;�+�+a��.k��6N�VaF��2��sH����lĉ�V�s'�Z�R!�x,"�lV��h\�L:���F�����Z�}ػ�]DB�0��6l&U{	�N�{�HeK�5�`��uh�����<2�����1<��3�gR���݅�/-�ѱ1��4y�xn�k��D�P�(��
�&U3Yu�%N��N��ЖTuir���,���������\GF`��(�R$%-E�Ӌ�=�o�FxrNtVn�S������cr6��%Y��~�&,@"8��^qV��J�5���nr���_���ppl�|4��x��'X-��SWJ�#C��:&;͂���ޏ#���iP�ˡ1j��Y���n�f���m��͜P- M���C���6�q�����)-�CC��t�4�#)��#����6�[�[�2_]/Y	�I�ş�"��E"N/4�S k$�C�"���QTPC,�ƪ�k�9:=)��&��^#(�"�.��kף�'�r!��1$b1iS%S)i��H�N�z1��@Q����y��� I�2����	�ŀ��9����j�����n��̴��vK��z�*������r��>�y��}N�>w�6#�{}Xw�2���sh�ɬ�bD8���}�?��ҹ��x[��'��7�N=�$8]��1rh?�ĢA:��ؼ����55d�!��f��� ��܃���kĽ�{:ocK��7
��^���,C2��C�V�<�D".?#���VDP��w�d���R���s��LJ}�����x�3�5�V������$n�|��hZIݥ��]�w!���|����3��N��P�K��n�!��*�UO���N��g�z�9� ��\�§LLOa��U��&�5f�w)
3���?�*L�ޙh��>���v_Q6�|�Z�j0��dy��,%�(�S�T��F���/fh���H��Uq�ט��=j�Fࡻ���＀���2���v���z�&X̀�R�נ��k�D���Jw���5�TP6�0��ট߃ɚ���(PWc���aZ,/V8:�4 Ü0��L*���R ��30ڢ,�u��t�E&Z�a�L>/��������d)�����]2�O��X�<���l/p����E���������$���(&wDC;��p������F)���U��*@��c���d�%Dk9�!-�����7ۇ�	и/����n�y��YկE0rdW#�Ʈ�E���d�4l�mYwHց�~Q��������S��xy᳚b+6_7T0:����|~�ȓx��(�v/*����y��`�ٱt�j^�����}@ذ3��$ �\)
}�����}��!D8ۚ0p�d}fD*��1٬¢�q��!���)f���"i��=�O+���W?{�-Y���C⽴oߐ�0�B�Ї>$�f8���xxM~v��:R�9C/��$uW2Il4Rv�ӃT����A����P��09B:_���B:_��O>!~<��{`3p��砣�[, v��V-�G�\>��H�-����lv�>�!�Z�����8��_R�4@.W`��@UEtf��qV�i���ߤ��,.�k&�x�y�u�f���occ�ϋ�����K�}�^8<���*�,NX��j�~&�\�XB�C���km���>��М$H�����a�qǡ���g/�D�7)���V�����>��HB�Ί�]4�a�ڤ R���
Vy��a69��GM�9��#����MN4��r#�a�E��b��)<��r�{���{;�t5!�+��Y�J*q����Ccx��71�	�74�op@ 1�OӉNشI�4#�G���3xM��@1��Ȥ�xQ/�N������	�{q�e���	�t{wnl20�u$:(���ڵS�D��p۷���v���[hl����.8�_q�$��%k������^x��R �GI.�H'l\�_��6�𞚊���	O<�&������BKSN���lE/�xͧP��`�g~·cع{?��L�Ά%���	�7�;ؼe����(*9r/��G����N�$0�]�ײ�f�� EzZ��rMZ��>�,Q~L��F������ͅt2Y44�$~��vb��%�p҉�:������1�5'��u��~�&�@������h�7�E,o׿/~�f��.����٦�2V�������[&�k��1N�L]������[R�ߗ�XUk�MI„o�~�~�ݟ�˹����#���Yl�`"puy=�`�]g�}�ߔ0o4�u�/������Tܭ�|��R5�R�Ԕ$T�g^�����Y��5m+N+����i���s4Z�AUӃ���A7d�!<��
Ԫp�0V
�T|��+����f`�d�H��WQ6�1�)��?��5;���ĚB��`>�fQA]�D��W�M����Z�n�"V�J�0v��S"zl�7�p������%4+/�\6}ԆA�'��?,y�E�_lG_���D7�^bdu��&����TsdCa��@�͋NW �{�S?�b"���� Ff��u�6�9�f���0�ۥ=�B2�S6�$U[(8'~Lj9���`��8u��ה���M���#_�^�;�&�ue��i���Y�h-H���+?��T;���4�#��o�Z�6���ؔ=�$fa*rsk��/�����071�6
Z6L�Bh[�'����R�q4)Nl\|.���0sD<CSK3����CO��t5���Fxw"^�iE�ՂZ�<�Ϗ�-�b��T�y�#`�"`q㫟�|�)�ߥ��wr�DD��{.�:;�I&��D����cǛ���r!!��l�P@-�3Ó���s#S���}N:�4$�%��Ő/0��!�ʣO<.Y�lE���NCK[�LJ9��L��	�S�|��� oЬ!Ȅj��x/�]���e��`L�@>�\Iڏƒ�b*�ٱ	��|Mtwvk���2\�^Պu=K����1=<�h]J%b���^֏���_S3jj	��	�����߈�}�\dBQT�Ea1�ʯ�m����፝�нd �v̈́"QXk*>z��q�E�F�ZL�٢E��,��w���$J���\CeR�eҙI�0м� �J��tPl�_J"��4�`&�؛BFCI&)���p9��s���n�6}��<�2l'�lv�Iz@����&�o2Sl�����B�6�/�߸A���Q#f���`jl�T�Z-�~�4yp�G�����f�a>8��_{c�G�=Y�a�Ȩ8�wvv�ɩ�XT�g�j��I�Xb���wmلxt���	W_}�|b|��6��=�
~�˻111.�� ��'���mp;�'K�-����~���p�����M-f\���>,�@��1;�X�w������46:%�����߹�[��G7�f�V��\Sw��S<���p9�}�����+1�<��ܔ
�x�5�C�XҀ��]���e��^Zd��m�p��w}�k�V&˗-�)�7���R[��(:L!�5�	om �zT������M7,�	��M �LIf���%;���n���9�i��"�~�E�sGK��	�~niϜ��l�h	���K�h`�2��4���=Vc����$@���
�Bv���h2ٶ)l��>�*Lء\��;�����_�hY�@�Q�q~߀@�A!P��$LX�@s��V�V������ڛ�Ө�_U���m4.զ'꓄�,jE��0Kd�����h���~m.#,�P���vIŀ�ɉ�h���o2802��@#
�cLY&�>���ȉ��
_c�	�Ƞ$�)d+%y\R��r��d�R���j���Z��r-[O�񡸐�L�"_o��0[H�j L{]�u�E,��I�*4�2��ߥ��XmT���]��@|x=�f4t���]-�)d{
d�2&�s���Fe̗�p4��Vo���*+����}'��L<�|:�݌��#���dq���LOF����X���"ƘlQh#��h1���t0�}�`R׻��]�+"��S�az;Z��g�w�����Q����T�����5Vo� V�ۈу�1b|v�aK]�ppߐ��-+7�����߆���f�O��ua,8���,��rV���G�gC���ם�v2A��j��c�j@~.��L��Mf���8���$� 
፭o��74ZT�45�vprtn�n�	/��4�(ʿZ�����!�**�U6'A�	VWV�>+ƦfQ,�rXS���O�$���6ɹ\�?�ǅɹY���b��~�/Y��e�84;�-`f��A��U��$��5,�a���,�0(5���M��C6�	,]�M�Mg�sxச�]�H���%��fF���sI$�Y�i�&#
l��Y�;P�^���\C�,:����E6�?�Gf'ѵd1V,����v�Fز|>}�ň����B����Σ��ɭH�hdl���@�f��+�u[)�n5j^Gl#�����0Z͢�Ke9�����\N#J�\v+��կa5q��"���=�jū�lE�f�0o�Ã|���/Aݥb��u�j0�����O�Zȋ�M�c��8�E☜����	����0�!�JHv&Ewk ->4{]���@�ύG���^v�%\"��?<�� �+>�)�رs�	�ca�Aďk>����Ũ�������'�������V��{�Y���#F�-#���L�}�Ǣ�^����     IDAT�*�4~��[�͔�r�Q.�b��� _�ʵ��i�����[���˯�����v'�gB���2s��g���m���ڑ�s F�ݿ�9}�w�99=������d��	ВM4=���&�Y]�J��.��?�{��y͉)�������j����B�-[N&lakQ��E�g2O��i[�������B��,Z=QA�&g���CFt���R��ϡ��%���I�4�ެ�w�a*�6ޯ�媟��٣	Mv��NO�`S�,0,`R��]���M&�VEQ�V�s��˳����[���o�\�h�	B�k~}���0(I�T+i�9�*%�j�e�"��2J�f�@C�>���=Y�u�7hf�������4��t��.�!������x�U�K0�r0 /h�jF�`ǁ`���=H��	�XФ�0��|��g$f���^��� SE[G;��Sax����Ş.޼�2�)-.�Z8M�
@\��>�h��yx���˥��]��E���.���(�#;� �ڠR}���pH���D��Ќ�l��1t������]p���ۜp�
�m��V�Z�`<���y��F��Lf���P5���|���D_�Z)��ѽH$'�je�'al���YT8l��_O"V�␯j���EǜO��D�օ��>�Sg	�t��T�2�؎���PgW��}o�XKØOX{�O�a�9�{��$2X�ݏ�� y�q�{�0cHb�둈�PM�p��5�E��p5��R�(��|%SM|��n+�.#
>��|qҪ&��u�[ ,@ӿ��
md�c��L#`���ׂ�\s=>��6����h����b>��S��@�a�ۋ��n����I�\I4�-��$�'yML��e������'���;�@�T���u��SO��CN��wjŪ����ep�?~�� �#֮�D|����)m<a�j�x(�	��)V��ѯW2fN��j/���i���Kp��X��/I	Ó����,��w)L�<����Ɍ�sT�RŌd}2����]Bԛ;;�xq?�3�0�h�8p��Ӑ��KT��	��~������p45��-� 'c]�p|�|����׆��9a��?������
*`w��JM*&��Y��D�YE�V�2T� �3YZ��}r�5x=v�Cc�g3ِJD���H���
Z=������s:=�&sr��{�h�_���b�}��) �|�t9%#���5s�S�bE@Q6��(�mR)i���\���qؑIE�[��������	�V��7���o�o��v�܍K/�ǭY����o8�Cg஻~�p(-���������Y��b>��>s9.��B�{�`<����#8C�j�l0,E���.�tcaAN�t��#�h��jG,6�+����Z�S����*f	�~챧q�w��L� E��(�/3���ƦMk�o7�+M�������O��������T�r�sE�h�������a��և�tk&����&M�i[�i] �<�0>F�[�F�61�0�֤����@��Rg�t��ض@+T�����3V�������� ���45-�T4�<?eB�Z�xi��~��>�WF�&d����1ɍp�n	s�E��N�ݵ��d���(J�
i���Gc������Ƌ�F�*Z�I(�(���@-#�RˢZ̋��WVǩDN�CX�7hգ�B:
�Y�Ԥ�|-�ƒ��O��V*�ڪ�ࢩ�݊|&�E͍�����V����.�ł������8槜~G4&�H�k>a� �vju ����V��ID��������%��T�hkmaZ�vH֫�Be,�år��#1G5�z�k�-<Y�u�Po�iL�"S[����O�z�]N9,�j����$ײ���%�]���~TsE�۶]Ĥ{G#Y��>�g_{;F���,�ц5���W��ω��^XÇ�	V���y�M|jh�ԑY�
��Tx ѝ[��]VA�V`F�]ٴ��6/��6-}c����k�����8*ꠊ��s�\Ů��e�2MO��/x��j����|2��D�l~����u�OX�ݏ5��q��5h�������;�	0A�b7 ����c��0�f'�vY�d��L_��&V˕�59P�d0`�����_���)"�."_ȉ�.��9նf�qػg��$M^�Xy����6JXU�>k�׎�L=�Y�\�����u6:��k�
e�=8��FCPN~q���	'hɄ�v��}��[�y�Ak��>DKI8��p��"�'�%�	2`P��hm��E�g���j����P��Ⱦ!a^�����yc�6�I,>���Ɓ8�u;
�4Rd�VQ�pp���Jő!xP8�-ذ�8L>�\(�3O�S�I��$̢�PQ���>�8�
Y,Z���-����4�#>��11z.�C(&^s�\���>�%3�ep�%��b�-��BV�����a��:��)0c��r2����aa1�U/�aW�tؐ�k����&$�`nA!���j���5iR���Vъ��7(����f��&8]8�nDc����|3�&#e�\��K��3G��T�����3���ea�|.3�&>����%.��s>,�)?��-H���ĥ���.Ł������t��!Ɏt9}��R+E-�o���~��$�_�o�����'��l�הL�}�Ѳ�4;��˺���*�s��cN���@�����C`F0�_�V�F�EZ!�e:rlbK����]������M�S�_�?��(+��?�{�G��+li����ϫR`��á(<�4L;��>��_;��,��_Z҄&a��]v�NXnٲE��a����^c��]�J��̖ު����uF�2ޮ�0�)��ݣ i������{�1l�IϘ\x�P������0m�������Q���D�[��U�n��EQ�<�Wa����?}��/��|e�3��0z�0��0W#0�h��aQihX��l��D�,|.��P��/Tׅ�NC_Z5�}��}YH*}��4w�~�6&җ�/��l<N|�g�;��A��\��� �08�}t7��}�:��{/�J���/{�\\]0;,��L��
֮Y�����H�XsC#b�0�L݀���l`t��mh�ꄉ%'�ZQ�)�&�RM���f�����`�K肋e��lR�'�~^�֬�	k�ᑻ�Cj&$��6���?��{X>�[�x�p#cØ�k6��v*�<vF,�K�Ł�V��/\��P_�B!�#����w�r�p����B�X	�D^�,B!���,ؚ�ۨ�0��@��7
�B��c��3�y�+�$�o��T��/?	��
�Mkw>����t�GйdFg永�/��*~��SH˨t9hTeLǖ'���a/)���a��]H�H��X{�zlڋM��.$�%ĭ�L��9���($y�FMF/mTb9$F��7 5�ׯ�9�lay��f�dS�ѷ�}'ctdD"x�n;�ٔ���fL
�j��?�JPe�j̀"�q�&��p2��D*W!k&��������Q������7���E=x��?���=$I	&��j�|�-��]�%SҺ��������\Z��<>o=bE,�Q��X�-��8�g?��,ڛ[1��O�`���!��._Zlnt��D�_��d�0����wI2���ɸ����nN�|

�$:�M��W�^*�"���j������Kp~u*:/��+׭��uk�������'?v�����f	�rC����O�DCG7�f��`�6 �V�Y��zX�?�t$�l�:,�H�"�8-82zH��LZ�.RI���V����{gw7�8�X�L�>O;���"�Լ�h���r�����,F�lv��������԰:]���q`I�����ɀ�R�!�4U��֨�3��%��H�D6�*ّ�^q�7�Eima�JiG�gO�e/Kf�سg�dGnw�����ڎ ���	���D��G�A!_�E�{�5_ī�����.q�g���@2��LA��e�ה�0#N����;ȯɪMOOJ�l����п�L�����F��UX�.�Nчr�F��2���� x�������!�w��#E�Z@�FMJ!�ݚVJ
Q���
��cҹ�'}�^��Pf2H}oӴ[ڇ����5������������D���#���19�&d�@�"�7Gs�焨NX�����C`�^��^ =�����&����2$P���M����1�LЋn��_�g���αǨi��f�^Հoa���Ω]���=�:4��X����H'V�0�Q��æ�a�EaA}�p[X�*<v��x�^5���KB�ʢ\�8	�XI��ZA���-�����vzQdL.R���-��X>�E�4�2EhPU�;�g��w?�y�ô�0Q�O�0�����0>D�0V%�ݝ0��Ȫ%$�I��)Tk��n���p������U��ܹRE�qo�۱-��T�!"fa�
���8��Փ,\݆���h L&��ރv끪��~<7>�R4����E�O��+_��M�ؽm�\�ss�V��'ho�;Ј��<�m8�n/j���{q�E����t7�$�������r�:���e���mG<��Q�ʚf����G�p�[iSR��鴶<�1�����i�uzƙ)��,�F&x�>8�*nV�V��г���նs�������kx���ڝP�&DB��`M�b��_nF?M#g��s`/���3"���+��7�3��%��4�1��Gz5L�5ۑ�GېJ&�f��z;��0%Y�?}�k����K��jC4��3:J��3�kxj#s�x��{��H�&��Zˢ���`'���Ս��y	��t�ftu�Iv����m����ˌ�ի�â�>�^��lO��|�'?���B`Q�-�����-���L��&?	S��L����Y�R��8�N�"`$9X�b��d�ɖ����N�6�>��x��m�ih��,����N��'d��"���;*��a�ܸ��d�@o{;>p��pݧ�Fz.�\Jc�8+fq��@q����]��6>3�F#�/�՗^��CC����6��{n�f��G�ar8�t�`2*h���|� >xʩ0V���c(U<݀�P5W�«ϋ^������b�M����_���
���<F�C��9�p�sY�OLk�}2�3B��0���\P����b��"�/�@t�!��oQ�H+��%ӟS'��0^c�s+6��jj�Uʧ��qล}(�bPK9����ɏ������s"�·���)���ݗ�`v��!	�m���-_�;n�f�&��_�
��f%���iժ�hmi��F��7W=��J�����ʾ��ي�pH�;�{���������IY/��*Lfj�
d��+�n��FÒ���@,B<6����8֯Y�?����wbtlX3I�}Hv y?$�Ǩ��+,έv�Jښ��<;�̴BR:u�C����M1�P�t1��Z��p����/�b^�Kޯ�b�ڌ�8E���^ۗu}�nu��U�R�>�0��g��B��:[Ȗ�@Hכ-l'��pE�3ZҰ��5U�z�i�B�M�ۜ��up��ihLKP�p�N���'���8���oay�o
�M�Ԏ��r�Mo����l��keؐ��m��ciO.����)y��FJ���SwN��5�Q��1*�/|}*�=�A�BC�Z�ВdȈU��e%��ec'�6������8Uņ}�'q��ż�C1a����X�+�S�����l��#�T��J��|^������V�ȢO��807K�)�.2x�H���s�&#���Y�R�\�v_	�7L��|>t�WD�Cf��M�4�.j�hU���3��ΠN��ჩ����+���~K6V��ИiVh�#�fL��Ԇ���p������^iǐڿ��|]�~lX�\*���`�#�B>)ZN���J�Z�Da9-ʲ����T�z��t�Z�5&\�3��8�A�&���齈�fMcղ����!Z�l��Xs�I�%����;nAHMC�Z���s�;�mj��7��u����.@<�ko���#�qxj{�5�gw+~��٤0�<ȸn��&$�zP�g%�;6:��J���N����H������A�-�.���,�ǧ�}dd��jB"�ݮ�j�kA�Y�uh������{�6l@*�G�N�6�8�������4��6b��}�{O� F��l/��
���MXP��#��T9/�x�?iq�kE�;͠�*m�*׬���Ѧ�gK?pX�&hfض��������_)�@�?����8<�n`8��#����O�P��	���"���RX�f5�z��7|�r^��ۉ�i<���������~ѡ1����T,��8������ �G��14��];��+/`$8+�;۟�/d�X�|%���U8���0s��`g|Z_�8��m{��|S6�v�VcJ>��\�qX�'V3���5�<�4�93M!��D$7�����?��dM�.���W�p�y,����El1�;���0%\�4�&����\�wQ7��Z�\9���q��Y8�&�9�^�aӺUx�H��1?5����񹫯A?5<��mj
���/�dzxl��]��:����;��FP��'?�?��'X�|lv����V��_����ذv-����v��I�f5!�M��ۭ�������s�:`��p���t�`vF+��#I❷w�bu�)��|�l}�{�7 �������ǯ�/q+��*���b,{ph��M���J�P��d9�^�	@c����V���hۨi�LӉir�BQ#|�������@��z�)�aPɈg�t�_<��&ή����`�i�( �k>��I��u�zk�lO�����d8"�m���L�{[���h��'I�����"ʹ<��{[�<�u�?��¿�_��i�����F��ٿ)Mؘ��~z���ց�+��ե���ŦU0f�p��K�e��3�0�0Ԓ0�dҠJ����J��g�M;���_qA�u�Lc�P��f�MxlԖ.�5(VN���-Ȕ*0X�H���O��~�yO+���#
����5�ٌ�i(A?h���@��yP����QV�2]d�T�*Vp���xߺ�"�<03��_{QT��a��a7�5=T���bo����ɚ�L	���۶�@���!�?^�#��\��X��r�e�)D�搝O��郩�.�6�ah�!�3 m&T�x�� ��r���-]p�����q�g��CE	{�l��O=��������y���U�D�B���*U0Oj�(�j���r�9w|��D���.��B���G�և敦od<��P(L/�1��E,Dxf��V���۱r�)ذ��j�����Eغsn���h^��߉�����%�|-?Z�^�]s���D�Qa����77��ׅƞ#!��i�l�p켾
Q)���j�Z(!6���|f;�l�ƪ���A��N��E�l�Z|?f�C�y\�������N���7��#�p��/@*�đ}G03�bw����H����2�?=�l,�Ӎ���ݱ[�}�leK�4��<�����y`t[ѽ��J�rN�X�*���z�h�VE�'�[��`ƕA�3#��O� ���5+WI$��omE)��[q`��hq6b��׮G_/b��0�o��&^x�LL�ʵ�wv��W�D[c3�6Z�D@K�A���������^�D��QmO����x��uG�k��];�-pjf�C�Ʉ��4ր��V/]�Em�"柏%�,�qhr[�����1T,U��C�ώF��J	�-h���n�"����o��68B!8]-�Y�FV�&̸�kA����l��R��)�M�(k��`�;d���0GF� %8�T��& cۊ l6��U+���.��ĕ��6�?<N:���3����[�{�;���}O�(X�7��$��`h�0n��gȗ+h���7#êKE�ߏ��V���mM8��U��g?��脖Bb�`��~�#G��ڙ�יd'a�%����    IDAT��.xpp� �Ca+=n���������pz[�{h�
ԗy�=�|����[ob��!����~�Y��V)�?�C��?�=]�H$"�����s��	6�Mlj%�_��p���"y	�1����:j2]ɳ�����l����H���=�� �:�Q(R�_C��������9�"���%
:�g��M�<�)1n�a���~ԉ���Z�Y�9�Pk�ЗSo���i��{�k�M��\���~f��z��٬Ό-{�~/;�_��b��~�-���)&lBU�����w���<k���fSK�ilY�Cv��	�>�\Â�JV�fM@/�Ƀ�ca�;/�&RG��&��bXz�u-Ҿ��夅ֳ{�0̚�M�$�Át���Ɂ}�Fq����l�"쟋H��>ORA�0�Ӫ����Fd���5A���A��GA)b>�R+ï��q����<SSh���Co������R|^dwG�ȅ�S��/�s7D� 1M�����iˑ��>��*�l[|�F�aG�Q�PE6�����ƪ"-a#L�� �A�6�w�����"1�\�fj�.9�c��%�	�C6dfr�=�$�vN8�8�������R%- �z	���H�\��:9�u��ѩ&Dը|3_wz��i}�6�mi��(QwA,n����̅&��ՃT,����X��T�s�%p���8���뿄w�ǲM���h����x*Q�E_���N,]2�H"�D*��Q1�$Ȱ7��$K��$a�|;�E�7���Fmr� ;̪�H�#�b�`��A��G�h����4��������~�/�l�Ǒ�G����I5�y�i_����œţ%�4�q�)���>�[�vb�zD��<����"٠�.��V����>'Vo<^�X9N��UaH	��xq���EU�i�Z�@o�9���bnjV�oV��xk׮E����n����X�h1��8TڛX�t	.�����ؾg^z�e�����d�;�b�h3���W��@G/saY�l�pr��s�ǉ���#�|��1x}>y�==�>�e����!�K����4F��x}����Bg[;��0����2����#�$f�a��n�;�������*�j�4�#.9�lXs%���}�̤s8q˙Ȧy��q��f����j�`:4�݄|�L�S�W&[��ьH4��P\r4Y�=��	�/p��٤
E5��V[w'6l:	�J	o����(�H'B����༳>�Zƻo���[�b��m�� �G$I�y��Ó�s�����pyq��#�J�=8;�������;?��C�þ����sϠ�ч������%qw6sf=�Xƛ�����
�6��Ũ�h��֠ +�~�U�����f'�pzp�ŗI���_��O݂D*%CTM>)&�}�?���K��x�/���_|S�e�lh�?4����v��	��/iE{E�:ۧn�G
�d�X%a�8qk���c;����V�X���;G�OJ���`f<�6�]�c �`��\�;�=����^�I׆	���N�i���P��^�J�R��)�k�y���L@�g8��k��;�e�e�`0�d4���a#y�������&.��Z)�d+)��1�u�r�B�p����A�5k-��^�u��X�-Zݐ�D#:mY�����5�i3	���WP+k�w���-��[s�"��v�|����r��r{��qۃ�b�ֈ�D��ԝ� �oK&�43T}���V4B��]fc����C@�W����Ͽ�6*no���Į�i��ew�������P���Daw}�L.
=D\�����C_A���2!%�f5��#�F=���3�Z�*̋���S>� ��G�G����V�(;>����54��ӟ���~�B��c��\h�u���$b�y	�X���:�"����m^�]xp���g�(�gݸ���U[
u�E��ր
�8�Wʪ�]��iq��3T���^yyz��aé�Ƒ�S� ����낷+��%�0
"�����$�S��B^4{�]�kB+����j�ӧ��S̿ύ�z(��d�6���O�P��`3��0��UA���Eߩ��W�A��aG.�#�f�f;V,^��˖Kk����;Էp���֢�E���V��+�2�g�1��.���T�M6u΋z{�q�՞�T���S�t��촢jRQ14���Q�|�B���� ��㹐�f��/4��$��i��p�����0j�hl��؂+/�\�6���#���gppx��y�*U���ZFwg��ɸ�s�-�	�
l��Jy���C(T�;x 6�C��MV�ℕ�����p�XL��L� ��[�w`,8-�%\��/CGs�����7�7ۄ��'X��*^�<���P��e)!�L��Eͭ����:8�??�,~��s��+p�9�noD����*ZZ;%(��`>:�� �{� lEҬ48�5�ި��������! � +R��3y>��Dv��AA8�@ss#�*'�`]�y<p�/���m3��=x��'��s�I�û7n܈g�}?�������o|�=���j�F�d{Mtj�H7n��:���v�W�/��&��Ї095�o}�[b�pҦ�������^�U��/=��l^M~r�8k8�Y�t��:�0�AI��X���ǝ�h����&�þ���F��t:\�����=�֮^irO�{�����o�Oo�8&�r)�s�A<��"IĢ�g'4��H`����Ә'�L��+�:g=��RՌY�e�EU���"&�l?Rv�~�J�w����8��D#��(�_A�!�������\|�ĿQN�H��][p! �W����#��l�We�� l!+����� ����BQ��w�F����@XL�宇�����ˊ�{���V	��(N?e9�3����ρ�����MM�Xc�{�NTaGUqK�f�s?��eAʬ0���R��d��w� qC��"��E$�n����r�bx�[��$�����?���A�݆(�˚��΀Q�S=���[�vȂ&�����H�
���0V˰拰fs��X�? �a;��?��I�?V�]�ž�Q3�m�k�W���ާ�5�Q�*F��G�&�#�d��L�|$���,��#FGr���[V3���I{P��̪9�Ś���JR����ľt�X�ڃ����o��ك�HH�8��.��Z���؈�~�6������4��d{���X�(�v1}�R7�mע?�u��@TF��˦��4��	45�M�x��y�ۺp�nMaA�~��N:��7�H[+��cbv_���aj� ^+:��!U*�b$�0��$VF�0a��Ȝ�٪"����,�U�bNک�%�(#�F���f�Ń��/�E�ZVŖ��e2z.�C[�>�h�ha��$��C&�&�cwわ^�uk����^�h���Ŏ�|X3���I�8=�P���N�H5Mb��.2M��A���)f�� �;\�F�$-V��,LA���n#_o�-Eל(d$��'�'�P�S��Qv�&'vN'�h^���/��v����9,F��sa���g��ſC6��H��)$Xߵo/�:���i$24ȅ�2p���O㒏������ho��\�B�&?~x��84>�
'���[��فsN� �t���9 ��6(:�ѫ�f�d$���n�W���fǊ�%���6c�� 6�Z���Y�j*bq�i�[xg�n���Z�\E��c�WM�>�Gq׏n���A|��B�s�EN<�p��$�����KO������Cs��.�6��׊������X�
�IL���H� ��m@Km/
b��ڡ%"A������e(�,��7�`Ͳ<t�OP+րR㣇q�}�a�����O��| ;�mǇ?|�.K��/� ��"���{C��d�
�ٿ_���\�+?}9���.ff�p�ڵض��aڷo�[����Bg[ �}�p�U<���x�&(�<؛��e�,S!h��X%��k�hs!�,c�ʍ���06���>��#c��tyQ,T�%��; n���I@b!�jre�u�X��_�X8�l:���x���*�'��XԆ�8�I�X,.'�ƙ����X]cy辰=��d�n:F��+�2�`�J�$[�'�_���.Sa�0�0�j�L��(E�M����#�PX�_�����s��"���}��-M�,:
����m�>}��Sr�{���x� ��S�	����9��ȟ������s����p�m�v�O�aݲ#����_O%s&��,^]�ȕ�0pZ�d���EMah6�;8]�eTi���,+-����	8�i�Y�(�7j>b��F�TVI�D�H�����d��CG��G��{�0;�rk|�����'�23ɤ�@�HQAAT@��i�����P8�HS:��P��л�F��dz/��^>��Ύ#���]������̞�g���gݫ���9��|^iu�r�Ȇ45�D���*LF4�7@� �J#��"I�|)�F�J,K���&��d����3=�P�\+��%�T3Е��2ޠX�`�7�b�ɽr�q�,��2�J�u�[���]a8�pA+YA�TFl���a��)�7 �Qy:��Ak�h�ҁ8t�
jt�r|N<���Qй�R['"�B����>X�z��I�d��m�kK/�O��0��zdy(�,�އ�� ?���+��NҒRM@\]x�p[�X��2s&����� �����w߃���@�8jg��>5��9m(��x�pߚG��sW.���^R�)~&��JޙNt��tR���4�Ѧ! &��[�)�1<������F��R�Ĺg�%���v��rRf�YN���}V"L�U��R�� �	@a�wCC�m�&��f�C��mv� �|)/�V�E�4*�7�T���uBt����-���Ҫ������rbl �*+���SSsԻȢ;�8�$���pL2�,Ofs�9����"��o'�]ði�rb'ðd�\�`���A����m���l߳�� R�"tf�(�3��g�'��9�M�O#�����G��!�����x���0%r{>*����+��N�[7ȶY�b0h�݂��q<��Kx|�S`��ь֙?��u4f�֡��0M�[g?�Z�'�Z�<�����$��Q�����q����-X��L��+.���G��{*��t��:�x�b���`tlH�l��LN�`2:a�y�d�
���+�;G�mtG�J��p�㹖Ё��cl|RJ���^��hV��B�.;��������}�¢���|���ᅗ���*�����ї���S�ŷ~�����ϡ}nv�?(ND��C�Z[��]���;D/��@C��$�d<!f��wcNK3.��h��ۯ?�Z�	6��TV��|Ved�ȮeX�6�)��[0�Ob�' S�bˮC��5��rR\��He��4##�t���+�T�Hg&�����c�F$ �:�c)��?����E�ļ��zmMⱬ�S�*!��� тM��1�q�:pRϖ��O#R�,��L�cg��ph�*�>j9�]}4�F�*��'Ъ�0%�VY3yؖ��)�Su^V5^����IU��ʘU��L�j;	�7�}:�8��{e�������'}�tr��c�*��ք	�8���(&�;]iz��Wn���C��V�֢E�4���z��3H:q�%߆>��u@�2�p$�3��=����`�D��9�RFmJ��IM뾒蕩h�57S3y��P�\"�ᩉ�B.�aH�q	[w���?��-ۑ����%��p�C��/LS3k&R�"�0�J43�u��L��E�W�O���cg�WZ�H���=jL��-5J���z8~1��А�(C�+��CiyQ+�7=j�Hc�m�[��O�B<�jw�E�&C9����ۑ�1�p:r2���M��(I=�
S'9Y(tf�c`��)�TZ�sKE�V4C�R�Lz��x*u���fjòHg��:<bbX�l1������X(�\(�(V���T�� ���\!�S ����-E�|Y"/���/@:���("��zz19���Xg-|u�4��pZ$�v�`?�^�,jg����1��lB&�T�0�I޷<���̹�!M���"��J�GTd	Y���MD��{�����"�=YC
{��+:�H�bv
SჼP+E���M#�;{���{�&f͜���^�3������RX:�W��^�"���	5՘�`9�J����>�d�t"�MH �^D~Ȉ��兼�d�H JvJ�ELI�.U�ĩ���������.�\�fY%S��R�
0��J:>C/�,嶣��MF���>
1]���s�n�=���g�S�!UEa�:�jl��+�t~混c��=ص�C|��ϣ��{:`��=�����h������/H~!������=�Sr-�a���'��&��BK,Ē�q����{���$��ށA̞?�.Ɵ�^���nhM�B�56aEG�8�;xs�Xs�}��k.��c�C��+���t�ڡ~-��J��d���Hũn�#����;����H	��t��y�4���v���ID2I�Y����r.���^�b)���P�P�s�_{��CHf�R��˃�c�v한7Z8�ok_�P,�X"#�:k�����3[�I&M
��C��ի�d�lݼ�]�X<�W_�}��{���Q_ð�
��r��Tt$Sf6�d��ġ��Ak�b<���#N��9�l؁��� 2�2&AMt���~	}=��@Mm���$�kl��s/<���9��
����d`H�5�'�n/B���MZ�6TT�im�t)�T��U�+��#���BF�F���S$T����*{�1p�,�I0�?Qe�SNFE\��
�
V��Vݿ������#B�U ��� �k�t)��A���i�gU����'�_կ�j��?�
�?�%����2��Ŕ&�?'1(Ui���Wn���C_��<�T!�p� �|��Ж�ރ�/�&�!?�,tO��I���'pߚ'0��V���!3{�V&�3o�Rt��!(�7 !E�[J����L���FH0�"[=;�DF�II�\sY9��j�1�)��3�j����>���jފPS�H	�#��t�E��,��bDZ��� ��#�� �U�A8��
���bO@Ś�d
�l	�� ґ���صfgd�Ȉȅύ��7!R�1�̀��㕘�#TZ5jjk�J'��fh7n����S���u�֥�1��u6E���:��at��H���Atl62.��<��橵+��*3��0�V-��e�B�/�E�G�nۼ6���2b2Wt0ȩ�h
��R��V�|�4:�u�B%�Z��4M���X�k�#����'.O�y5\��f9�Q�����$u�왒t�D`��$���h�;㘐���JK�l�lQ�w�����2_����8 <^7Lz��j�y���;"O�0f��|BR�Siz��^�LdQ)�aҚ��k�����ĤT�n!���׿�u�vuuKP*]��TJ�#-vb����5��P��r���ק��?G5�F/�?�L�wq����z���\�¦�Yh_��v��,�{_�爙'f�ٌH4���!S(��Nb|pXw�Lr�N�Ǽ�64�Պv��`���t�X7��XB0-1a1���A�Y�	�����1�T�29�ik����:��n������#�z=�,[�9�ڱ�͒�m燢��p�k21{F<v'Ar*�Ø7���㢷*�����T�"�c#hq���~K��'�y ���	��޹hi�+���G�\�GC����*hOe
�԰���=k���F��#�S�蜫檣��d��x"%���^Av,Y���Ft����H�Y"G�Â|8�/�p,~q��0�x ���.�&aqX�>��[2�V�����Q�7k���C��Ȥ0NC�h�5�͍���K�z��D4�s�='��UG��Q��M�0�ׇ�m�p��.�V_ě/=���q    IDATZ�v��t��~�>S�H�B� h�*d�)	��*�=w��9���!�z���#{jw8Of�b�j��}��q��Zx�>i��f�0Z����e�U����ܳ�pp�hu*��9�3�Sr�|SR���po�r�S�,S �
Z$ύk1�~Z����l6��f�)�8��O
�s4lE�f��g����/#�5��2aՑdu�Xa|�.�K�C�L�cAN�W5aU�4�	�lH��M��P�Ӟ�tpV}�*S��H�0_"*��GET�*�|������:;]�X\>J�q�u�q��Ap`.<�L��AhI�"0��N�a���6��^Ō�EH��(��"ZEثTU]�JN�"F��d�V6-.A�d*�{
��p�0(�SL@I6
�n���M�-�asz$ހr5
���$�ec�B�xq���'�%H�P���Y�Z%#I����Tz��CO�J2U�nNҼE�*��u�"8<&�mZߍ%�t:z� k�3�H&M:"e�W

�	�F&���zd0�\ˑ�c����� �,K�ĵH=�?T�X�l@:#g�*L�"���d�(d��J���g�M6�l<��'����W�3�K�`s�01�/�F��se=�qnX6'��s8�؁\.�UFw&�����(ymRh^�
C0�Q�����f2�a�*�,�F#�ل��((�x�R� s؜r��m���mw#�� T.!�� ��Am�H�o2�o�w�a�0�NC�t��bϡ�d,��:�rS�lZ�Y�29>�^+j�Qv�v���<,V�0��}�����P��d 6@ɿ�J�l.�E2��� ����d�1�Υ�/��+.��J)�0��B���^�I֒�sd sp���p8l(T�e[PP�2�i��EF�>#�̛�!�d��6�gJfM��:�*v+�d���&�09���
{z�ǒ��`m^����;�4���~�x�X6��;��}��NU�o��#
u5�tN��d�F涷bv�,	�L��Z�=�tt,�|B�.u�s��%2�s����5��0��+�>
F�	���cuL2އJ��d5.��_�瘳F��c_ޗ�|Zh&����h���W_x�{�E���kXp�
�P��᰻��e�l%1]����Ǆ?��y��GS�,8>�x�ؾo��Nƽ�s����7�Ί�/�Be4��ko��iC��^+��=Ff	ayG+���2JNF���b�X�R@��v�O�����(g�����_����f@�C��f��c�u�\���b� �D���5�����Տ���u�q�_V�s�vd3��9qHrv@ى8�*tCs��ʚ7���?��Q�:e������e�!1�P{��oM#���i��.���f�\�p/�l>7�ӟ���u��%��qc��0��ὨR2B�cKIE��	d�^Ȓ��d���Gޛ�xO���=���橕u��ĉ'~+���-�3�U�B����?z!yo�:��x^Xu�X]ӵa�>E�h<͙��U���k:k% �cگ��)��2���*#W��������ΪU?_�ه<�+FT�D�ѿ�U��ڢ�}�>��y����F��8����|o���#=��g�Gj|6�C�yx�N�T�ƾ�>���;�zj�7z�W+�'��Z9MTk��⸚�Q}#���-)��+iU�$�������r�����)������*�X���e��|�a�ՠ��I��H����"�J�xYOZN٤�"[L�-Q����+�;؃��.�X0�7
C�䭅YF)X�&���Tt���R^Ɗ�r�\F:/����t�+��ac,��$�X�K�T&-'9��F-J���p��;L�E�j�������=��kF&���و�l��D8P��
"�.�|��'��"v�(
���F��(i�84<*�C�I�%���`s���С=r�Z;��1�LY��Z2ӡ�l)�h:-"�lQ�<���Z�>"3��e�ԗPa	�Ռh<��A�S�X1��T�K���L���N�������t>#��M���P��T�|5I�v���E#V"C��u�0����'�0;]SU!ʩ3��IbFc���J�RI��3g�9���E����1��Ȩ��CL�f�O1S@1�E9��Ek��.�^�[6$�� �0���ec�g�(Ӊ�ߑV�O����t�2�j�x
(d�b�������&A�X%���C�(�����1*k��B�Y�U��I����HdA���e]��&�M�ύL��h�VgA�BP��:�pȑ�����b���<�e��U����E���=S�E+.I�ܽ�ܫdfkj�h�Bx�^a���FG�$��b�I?lF+j<52#XǮF-�N:�派�G�Z%�m��;vH�9ǒơV����c��-�ޤF�RF� TUg#C���,j���׎������눅#�}���-GcC����A���尦�$��<�xZ�m6�=��1��?����*���M�]��'��V�s�G��4?�h�k`S�Z/��`q[��fX�@!���=;�A.��0٭hniA�����N��cR^�ē���Ftv����x���u���C4��nƖE��l!:)Ujܿu	��|<|3�����B�-@�!������!���A�Tf0��M.c<�ƧN8Ѥ
�mځ5O='��#W�Ċ���<��� �FC��f`r"
�ь�/��݆�^t��������f�I���dT4>%�zo����T���zE	"�mx_+��S| �/���K��:Ǥ�l	u��B(�Ivٲ%����P�gEVI�Пꐜ���*x�FOTG}������$蟾�Np��R�7j�?��M�����~_5�L	_�߀����@�H#*�n�Z�c�F��J�J�H��ǿ�;�'Q�y���nٴ}��Q�8�k�w�s&���a����n;���B߾=0� Β���ӊw?؂����i��M�RtO
��G�'6-���@���ݐ��%񻇁[���^tbd,�ǊF[OK����7�o.�l2 Ԅ574ʩ��޽2�\�x���	r$v��ꕘ�j�L&�p�u{�`�<t����;%پ��z�~�����k���W�	�y�Jp�T.�r�c�xꙵ�8m�S��?����K.B>�@�ۃ����[\�>
$l��c��W��\U��F���o�7g>��{l�Y�d1V/^���{a���r8�L�M&a��7/	�srb,���C0������c�h1j��P�Q�d( ��,�ۻw��fu!�͈р ��VؾP"!���׀�Q?ٲ��N�>��R
�A��As ��&/r��Y��^kD�:B��\N���Y��!,ik����<�tF�#q�����I�9�T~�Q!�Mb2��W�݉��I���bX�v¬S�n�"��#3�Q].W�M�df��C����z}(@��J�X�`9#Ya&���;=�����wRr���8�n'���lRj�A@&��Ia��kk`ՔQLFa����h��\/Z,4t��9VAg2���SA����D�q�a�a3�F�c�UA��Xl��}�)��S�+4�i09�$�J�OU+�c��"�Q���e�je`3�p�gN��lŦ��������#�b�!���!�k!���q1�t,\�e+�������`t`�w�B��F�2at�q�(;%k�
9�J{C�"�f�Gq�8t�SD-e,��S<�ı7��`�	��0Hz�	�DV�Ff��X8sn��/1�y@��C	��C0�YR竓1�^c�kE�1���!��Q��z6�|Wp�-��P�_�a�o�}�j!�+!0'��=̊!f�I֛��X*���R�bɐ�Z��}�KM�M��804 �잁~Y�7RWS�pЏ���6Ob�1�m�E5�{�$�~tl ���K�{Ι0��Ȥc�����.���s��X�p.�.FG{P.$a2�,Q����rs��.�k*C*[B��A{��X�x�o��_��U�����m;�㭷��y���0�](T��4hThn���?����x�/���G����V���R�my�T��ͬK���R���D(�\"��Jʯ��`�}r<H1_�قP<�3gɚ<<8��N;K-Fׯ�Y��WK6�ce��W%2ܻ���UGy����r����΀U�A��G�U����R94���0�5řT����/@7�[���>���8+6�	�TT�*��j�F�J�RtC���OV�����6n���֖:��N9��n���0�K(�#H��c�K����İu�&|���������Q.�8�2\��>���:�"�,}t�J��b!�+��Oʱ�*�C_
gR�ΫP�ǔ G3{Ŕ�U�;+@��Y5"�!'^�RD�Y�"�X�?w��K� uM�����ϟE�7��cCR�k�O�'@�Ն����M������C�̓R"��1NX�)���&b��D��a��^�|6+�#n�F�K��.��%0�B��>Ԡ�ق��y��a��m�Ȧ�2�jkkC2�MM9GI�l�^z�]<��k(���= V��^�\���[_���0���:�	�l&�G�<u::�Ȥ�غ��vϽ�4��@ *!�,nk��w�>�d]��ʠκ&��xܵ�ڊ���,&��q���kx�o���L��-hdSl�𝯞�|h�\���}M�h��i��d�PӒQ"0̡�W�͛�����S̬��l�`��+:���N�&�A>�����!��6�ז�,��h8���D���bY�)f~�N���X�xc(�R0����\��M��"	?B�,���F,WD,�C"���d�M����B�ωx8�ӆD2&6x���F :���+�*0�mHf
��H�5�&�5l7�xX���8r���8��:�2�<^6_��1F:pl�2�el?Ꟑ���v���e�K ?��1��:�}K����ᨢ�!�1ۥ�/G)S��d��H�Y�T<�B>%�P�>�q���r����oa˶�r_ۨw ���� ��O�̡Va��Y8�K_���ɱI�Xפ7c����:SHOו�����N������=�/��V#� �0�㟪h��d�q�O�s�.�*�b�G-��$��2�\0}�(�bk��w1<2����%�3��c�"haD!ϗj�No���E�,�Qɛ~�[�)$R9�R)��}�װ�@�\�r=̲�-�X��u���\$8�3���kg2�����˟��c��б�9T�OL`��M"� ��H�����?w	:��-;�b�j��IQ��mC,���|7����C���ԊPF���a�d5�Tr�B����i�F �5�H�ɊH8�Z���1ح6��vd
��hQ,i�m�Ȑ�������}��G��߅C]��]�����:�uޗa4i���~/<�#~�����D�?(�n��JE���b:��	
��,��B)�d�`�I/:e!��{Z�P���V�qF���0���_�",X�Z�x�������Iu�H&I�f�<��,���՘�*H���52q*�|:#5����Or�>�?=�4&��I���"��p��B�T�����Il�<�0a��Pi~��j׫T*΋���6��s����[ϻ�����,�I�V`��͘�A�'V��p^���N6mو'^xf��ڙ88<��݆�J�)�/�.K����)����˓'a���[@��>�\$n�'E�(�
�p<e�	��"k5�����lUV��c�>�* ���3GJL�������!^��2�У�/���^2���21R�B�RA�B�^�C=���F4�k�59�Dp�w/ç�9��q���F��\�F�XydUX��;>�݂^wj�0�����lA�׋�u*4.D�8��������$`��R�Ѷ`.���T�ڗ��7�ޏ���B7S�ː�������6�Pg� ���j���$1Лd��g�k>�tr�� ��}�����a2��/㦫.Fbb(���k��S�D<�lV)�5YLpչOE�E�?�/��:j�[��?"��7ήq�?�4� &Ry&7���P[mF��	d�!%��~�ǟ{O���^7�&#�k��ݠ��R��W^���aNC3l6'l�u"�ey�z�Yd
DsI<��3ؼk�DqʈQ��b�����e� � eRk�s���Ԋ���T�r!aɲ
�=�����c9vT����i��pˍ?E�(�2��L�#E D����&&��?���!�{���ꁾ�^����E,�5߿�|L��H)�*��pC��Ș:�H�j�!��K�����#O>��ׯW";2)�z�	�g���^��İw�Sy�j�e����^�"�KI*7�d��g^xѤ���Ē�B&��桩փ��:��㎇N��N��{���mb���x�w�1�X�dBI%/�p�b\��`а��N��(��ڃ�#�˱�Q�����_=���h��~�5rm����;7\{��Y7j�x/���,����SP	�����=2��r0"3T�sHr�͠B)���gΛ'�=�~&���D�q�j��gܮ:h�FI�כl�h��cR����ob���8�o���O��F��<�g�	��`,��f�l�U�Wc��-X�����"��a���ww���ƙ����>},4jJ�޾m��&�����K.���}> �#�QU�߿�l��~7�v���N+&��p�l����y�u 
J]�Q�DPc����@�lӋ�JGE���1��^t�nv��P�=�$�f��������s�<c&^{�-�jk����c/X�!L���G c����"�H+`%_@cS��)ޏ��<��kע��&�+�J�*���*6���+���(���TΤD��K�Z���}���H�%^_���<p�	[�p�aVRd���$=J��V��cU�V�D|�|���:��>r�ph\9�؜ꡬ�;e�:@U_c�I�������_;��� U��x]�ǅ����Y<^gj�fW�+�Z�f�J����?�- �@�R���zw���,n�w�2�z���`�d@c:�lC����FO_7�t�h�ݎ����Ko�����`ث�Y�C�s�
e�>��Ƌ��E���i�����7�r�O�ǈ��sr:/�&�)�V�x*)u �
��):�2%��:�Rx��,o|E���`�*x�O����<�: �Mh�^ڱH��J*� �"pe65M�N�%t�?��6��h���sp��'�vLo2�R&ݮT�P�L��D�B� �E�m�v��^���3109*��/�\�=f�A#=�^��h���X4o�O3�0T&`�?�_�v��9ŬP��kU������퀺�G��p: �I�N���0�&���v������B�D�lf��N~w��0�ߍ�xG.=!Pt�,
z�ͭ-H�0ڍx��o�����!؜u�ia�7��#�3Q���*f��Y
���\v�zC	(&�X�5���o�
[s#zF'�w;f3*��3����0�}��kd�<�t����=R.���!]����݉MnAM]#����=�6c������h��u
�VR���2n�.:f�2���ǰq�^��NL��&�p��hon�e����������]�&��p�K�e�!��Ťߏ�<��۾����bR��-�pD�\|�yغ�}�mmÒ��EKTH���ؑ�D�ߎ�W�\�Rx�>lض�:	J-1K�l����W?</?�.���C]M��o:nK���=*l^{�M�E,�G,��C�^E�_��u֙h�zQHE%��"nn2�[mnؼ5ML��Co��7ވcȪ4�f����i���ļ3:0�ьD8�ۅ��1,]�X�m�
MV�#.���J��5��j�&�8��U��w����Yc��ج�<FbJՓ0�4i ��w��B�� ��!��Ak�k/C�-�4�|[��f�	�����b�g�����[��Y�-�0f��>��P�@����f�>zV�h��j���0:��� 5:a~��X�&q�s��l�L�%�xh*�1���ŵB    IDAT�X@"Gogzz����o`�GbѢEصg'6oق��~\��Kq����߸�P]��h�7W�+�&���������5�A�ԑ5҈X�f�KTJ"�����8V�Ǔ1��i9�pM������Ƭ�mbPb�1L�_z�2̛׮�456�8�TR�T�h�H���2<�����"��
��$�{v-�>�FG�^�@��\|�ša���N�#+���A�T�%�D�p/�B�Ä����Ugg(��x�I�W�����?A�Z�H]��E�Ueq������lY���Su�S՘	�!--�p~�i��0��8�斜¦3g�EU0UՄMEN׃�ߴa�{M�fk�j��*�J�	�����4<�ֆ+�ڰ��G&���9aN��J�5q�j� �
#AG!ٚDCã��Q<����$j�O���(���>����T��BJ�	�SR3�(@���I�<O��3'��n�n�bZ�W>C*[#r���s��%�]�$S��s��0�ȸ�s� ���&�$�P�ζD4�ņx,"7����Gv�#18؏ޮ^y��;�҆�D�\���$�%S�c�K^X%�ł9�p�c�x�bšVJt@,�S�٠�K�6�x�i�y��h]؁�hX
����D��ϝ��>}�V��H-12�/�#���ՈTƏ��X��<��0�����"�ϦƯ���6+~q���7.@Sm�6���sS�`c�N��l��w�r�p65!^6���K����Z\��3��ip�7�Kg���KWb|t���"�;Lpz,���hlm�ko����>��,���hK�7�Ǘ]��x?.��R\�ݫp�	_�Z	�xN7��LZ��rl׾�"���.\͍��
Hr3M�P�Q1��/�֏���>,[�
ǜ�Y�ci�U:�]^8�6���d*i���=<��Yh���`��B;���[p�x��Gq����
����(hd�1x�ȥ#��xb݋x�oo��#�^EW̡��?��՘��C�<��Ym�ַ/��j�e�ʴ��E�\
�Y��7�����D.�֏��>�	��y����7�Сq�2�19�1�;��J�H��4�y�l��C�W;��#.]��+����l�FFP�+�Q�.�%�G�7i�e�kM-~z�o1� U� �CWLC_�㼳����=�|�P ��pf�̒��ŉB��迦N�w<� ���	Xm�T������՟�u߿N׵��"��n?:<���Z٨�A?��z�l����WJ_$G��+p�8f�J����b��b�"k�jaq��~�jȣ,���{��_�:��b��tOR�&&�rNک�dr`N[�Z���l�	,k_�\$�7��p���K4����$�ivX`�8�ƺ5kP_K)�򑩔�̤a3[E�Fph3ꑈ�亴ZM��蒦/�<f�	�\w%흁�	��M����{_ƺti�%���.��m;>�����	������,��@ .�N����X~D��^s"B&�n�y|Q#%��8���ۭr0d�A�#c�����{�m�.����.U�U!���Kg~�<�	>����\�y=�̈F#p2f'���$�]VT��p8m�=F�y�������P��0sY��5�TFi��"�I�^[
X�F��X@�h#K�u����
8a�wXMG����K�.`ɽ�����v?J��z���}Q��v:-��ǵXUB�
�(`ȬL���ǯ��(�__#V����UinQ>������)��'�Y��a-�t�l�c|p��Z�R�ח+��t��*�T��;��?��?x�o�/������.\��s1���*�U�d8�X$�ٍd��Q�����?4�Ɩ�
�!�����|/r�()H�.�j$�����M�9T�0��ݽ�H$���V�`0(7?�N�dq$;��`�/.*!�ӎl>#����O�FxΜ9S����R�mZ���b	k� �}�4@�$�i⁾~{����C�+��y+�5�V+YD���).��h�����񩼸�lz�Z�g}�+J��$��P^��`?<N���(�����SϮų��Cs�l&K$e�eą���9g��s�8��g#a����V0�
�p�-x��2o	���	+ŀB�Vmg�|�|�1\r���8�>{����D��(�f��/>��7����V�RPiM�$��ը5�1N+~��[���D�<>:.�d�L�3�V-���"�}�Elݽ�-s0�hs!���g��z7Z\N�p��p���g~�C2�����#p;t0�5��?��Kxs�F��10<$��&��P�^|����:\�����4����k��x�8)\ו��KO���o{58:G �
�g�·��5h%|�K_��7���~&&'`�١3�
�Q��A�.0�Ͽ��$��Y�����<Z�q��~��]��/�7��.�����త� _J�P`>\	:�
�?��ܴ��t^�V�I�~u��ؽe���p�e?��?��o#C�2Jd�p�k,F������-��l���mjP\����_c�ƭ��onê�G�o�7��|�j���$B�I�2P?k~}��>�
%d�	�A̮���9'�^m>�g�Z��p�� ���sa��eie��K�uo�����BAK�C���0N:��겫Ez%�#{���DB�a8R*0���Lz5B�(.��Ja��l���	<�<�����F&�DA��
-B&�5�ܸy1X�a��v��on�o����9�
�ux�A�(���2���k��$�b-�f4���T���/!<��^ǂm��t&#�>����p�?��v�T1xY�7�����ʶ�TV��3�-eʺ��-���v���Q!�O!N�Vh�����~�ضS�ot�nݹV2/ N�k�|Z��wj�e�B��0��߁�z�� �a�+�
̈�à�	��1*�Mr*��d��9LCp8���Y_���$6� K��Z����ϯ�gO>A2
���N��^b&���|&�b�����Y��v���<��x|ͣ���͐���SB*f6����@�s�Ai�HaTZY�MS�t���tM*�|�du��Q��C��S#z0�t�*�=E���c$$V �T\N�\���4��H%�0[�Wtld���	t���:�tnZ���#{�[�?�zӌԃ����ů���R'a�ܿ��z�M6���ȟ�MPf�'��4�g5�������sI�'0kŊJ��F��0�G�0濰�/o�rYɤ�e�a�y�1hk�`��&�sq8�q�Xm>ɐ��__�s�^E�P�<.d.���y�L�8�Qr�㤝|,���LD�����d�<c����ҷU�ϋ�_Ǔoz�*�E
�7���z��Û����<-j��(���*?/H.:n6A%��M��9D ǋ���� ���ʑ�MI�+O��IѼ0��#F�z	+fw"
a��8�_Q4on*dӌ���X�y����Ë��$�	��V�Y���1����6f57Ih.��L<�\>�ێ��Ay�V���+��8�^L3���Zg����a疭���bт�PU4ߠ���dP�9.,F��?��
�Ո8�[��8�ґ �Y<v�Æww�������\�l��tM�f�V"$������kh�ي��Ȱ^�j�����d�x� vlކ_�xN=�4��ydrqv�������Λ�ǟ|�vJ5;�CI`�QJ1�f�Zf������v�6�	���E�M�׬���<��lۻf��O�e��5hr�!42��＇��-M-⪊�S�k�ojDT�_𩧟��%C���a�鐉�q�܅0B��|?��'8�ӑ�d`����HdE:@�,X<���M��`���h  ���	ߙ���� <2���rn���X��|V�Y���:�^��#�
]uÏ�)����Qq?r��3�����_�n��z\�݋q�W���[2縘�U�H�������]�ݏd��`:%��j��b�	�:��|2^y��u����.��vZ1��M"X8��O���߇�+�¯s���a�dޑQ�l�¥����!�"f�F���jX��%{��Q�C8��}#���$�SSǃ���8.:�����d�*�DA�jZ�+nez�n��rN6���A��W�@"WCGZI����2��T9􊾈�}���V��Ӏ���I�~Q^X�*��it^�V�̛� �h�[��}��l�n�
Ah4��a�YجF�s�*�2aO�:�AR�<LV=�4�.�����1o�lт1#��`��P�n}CØ��*u]G�<7}���7cp`�H�lz�MF�<$��6�?�+ݖQ��V$)�mN�6�d ���{!�cX�Q���D6U��5#��{��;�[6z���y%/2�����g?{"ɵ�$�.K���^6z��d.�y�`�{��|V�+Z��<�<�������q�W;k�T�j�`�k��S��xT@83��J�a�23�j�� ׊�-|�s�k�˯�@6���]����:��x<>�
�a�Se�J�YM��+��V�d��;���YH&���Q������2�M
9Ac\�Ӣ<>�8FYU�?	*�j��f�2y��J�"YK:���ɟG[��2q5+ݾƠ�gVXG�� ���Ly}.�Sj��Ν+�;��d�E${Ƚ��C��d빗�a���U�~^o�����yQ����8� ��g7^�ʦm�k�fh�:��������c��a6�79���==x���%���T��./e~M�HY���(z�f����b��\Z��9a_�������{�DGטFho�8n��LI��4Gf�?�O���Q��+ P�����j	5`�XX��q��hl�������� ��������;���Y'D���<O^s2�:�S��rY�9�:j%���W���C �(岒�C������PW�� ��1B�����xv��8��_�I�>��3�(W�w+�9��bd<��[�b2��nF*����jw�nrJ<C��G2Ə.�n�fC]MS�d�����2Žoh��~��(��h-�4̟9��b�Cx�P*���I�<�k9��zK`��14��������R�F�7#hoiæ�>���7���ނcV��������,�(��a֜zlڴ���C��ȗU�&r0k��w7��P?6�}����J|�^GO�J���lm�o����w�b�!!ĸ��N�U������A��� ��{��]�F5�v�oߎ��v�1��!�!�
�f4bq�\lzo�^�~u㍸���-���c,4��UNI�[4��]���!$J��6��k
��Y��]=x�7q�/o��G#O�}�p_m\.'tf=L����(:�lAa���U��uc�k�7n�u?��~�k��d�H�<,�a|椓��3�!�N"U)�܀uG6�������<���fq�5Ի�vٱ`~;L+b����t��[0�OAc���S97M�ys���.�G67����8��2�6����Ō��}�=h�ӊ�C]��1�N�����0oN�_ ���O�!J�x�QP�j7"ap| 7����X�=,���Ũՠ�)A�*Bo`�@�B��-�[�r�#˝MFQ�s�������{����'��݀�9m�L���G��?܎b.��J�V#N�??�:uc�ҥ�#��9[�1�J�ܜ�v��a��1>6�?�u+l�B&�K@*Y�K���m��`N�<�̞�����Jd =��"!�UR���)Yj�L�".��l�{�@�.G��lv�]��X�xXʩ������ю|!#l���v��q�5?F<�V$d�4���(��H�"�����|�x&jS�E,�X,/��J=W2��J��A 3�j=n��T������o����% \ں�	�~1��lݰj���\�X@$5v�7�-;RBv9%�aomm��/\�(y!�}��.�l��X��`~b5ɞ`�nZ>�0���v;16:,��<�!)�f�x8pU@V.'���lU��i����
E���ى����I�j�������7>�Nd}�){8��{��o>~ou�柭����\�z�>7r��<�X��^���٥�L�Z�q ?�'ǰ�y�3�����܎�+T*{�߀��_��+��z_�?����n�{��a��Pof�[p�Q�1�΄94�� �#N��W���v�lq�M{3E�
+��q���?��E@a>�,~=O<YW��&s����bN.^j��pP��㘆��3Z�rr�V�I�?���X�)ȯ�{	�x���PU���Omt�J,���R���f	^����K���%�|fE������΋�s�l6-ϟ@�|V�0��j4a��+e,yʉ'�͞HF�� ��!nF�:��~���Id�X�j5���+�tu�ٵ���Y��7�х��#��\옯��Cv�������px�$�
c�
�
���Dch�و���T܆s�H�����*,�(��Gq�/~�x��3�6�"!9�w��D1U��G��O>���N��"����>�4h�%���%<����"],#�禤7uy�=Ø��W_���9�*H��/�Vϣ��Z�8^Z�>�@F�F�]���ᅮ�C��C�C���G0ļ%:�4�42���0�R#�8֮{�\Y#'��J)f���zD~�y�qY�b�*%���`@����N�ŭ����,���`C��h�Y/�`>F5��:�A\�58��FB����.��(�3���փ��	��CAk�h $m�LƊMn/6��6z�/�K,_��@D��\6��MqIP��ۆ�ع/Ѡ���	��*_���l~oz��E߽ '}�O�6��~�fŲq�b�\�
o����A8��Z�'$3Ԩ��u{���}p?n����������Z,;b��g����Dg��o������p9=S����X���蘷H����r�Q�>�;������-����<d�Eї�bqa=y�_�d~z��(��i�@�Q���F�F��\���q0w�&�ӎL�"�$�Xi8*e��U��2� ���F��(�܃px5n�Jyx6�{k1gf>ܺ�<�&v��Fm�l44�FO�/]��n�C���e�aq����??�Վ�y�i�
���%r
�Y����r�DpX.gq�����V�K�a��Eq޷�G���8��S��_�6 �z{E+���0aN�k�C8��#�ӟ�f-�j�ѧ�u�V��w����{�ףwl�!?���d6`��W�ܢ�(2����8���A8;�{oeW}�?[��̜q�I�CB	n��\n{oK�:Ŋ\��C�X�[�R�X x �>��9����gz��k��^�[�7keMf�}l����|>�0Л�q�����7�c┉���uڮڱx�b���Po?����x��ՌfL��_���3s�����+�����2���.Y^]V�M���EsK�<����x�u�Q��6	N�G,\$|��/�qR�H�{Y����b�1�MFZ��t_5�@����o��f���eO�s�N��ǧ��$F�\�{� v�/^�]{v��y[�^ޏ��c���^\,J�n���r�SE�&q0�RHq�kkk��J���K�f����~[�>ޟ�õxǎ�yS��$�C�;���!�n��5�\!2u��-Zz��(��m,4�x_S��r->������������������p�4��b���x�����=�Lhhl��U$:B��F�8���Mɪ��-Q������Dd���زi
*|d�i�l�
}̊��lr;8;��#O~���I�l��B�ڥ�Z�y��@ֳ�����I�����(��,?�&S�$��5"�&!~��&�1B?������b����&�\�jke񡲲��Q�M�І����δ��I�*���Đٍ�6cמpx��g���r�<��3���1����q������~&<kX    IDAT�ֆh(��U$:�L6��>��ݎ��脃[6�`�d���%G=�HR\�9�\�h.8�gV���.���SI<u���50ǹ��#�,�
�ET�BH�F�"�@Ux��G�m����5�MhFE�'��Gc&ʪ7�z?>۰����^�'1�l�]~Y�/�跘;k���XEqC�yA�WZKUTze�X}�CX��c���Cdp��jt�QSY	������v=�w��Y���p8u��0�:�5.��*�߹��+��\$=��j��t(���^�d�x4*�%�� ����
97��]����;�u��o:�rPԲ����Ћ���rLlm�s��IEN^P��EltԊ�)x��7�eo;�0�I�7�n*�n�X��t7�|5&O�(�ذ�
��)7��Í�h[����`�Qz�|��~|��'����5�U0JyL�҆t&!�C�=�QWTV�w(��b��>q�O%�(��a�����&qO�\x>��ݎ9�MŌ�1c�\ܳK�av^|�U��ׅ��I�$�����̨�g��ك�Y<�8��1yR
���Ō��_!Eh./�]����+�#�	���<b�|�rTޙe�޵�on(���F��oٱz�0��`O<�J�2$�ib�.�3 .=j1�9��.���])��:,�Q
B�
�'v���7>Bo�(�.'&���ѻ�@Uȗ�9lX���x�gQ]W�P�������(t
��(.`T�.A��)���{�-��L�;锉�x�~�L�.;f9�mX��0x��a)p��M-'y͉��+65Ǭ��n��ɢ�15.�*} 7@ȿ��Gq�wc�������mC��\��Xy�-����=>48("�,rT�OeP �M����<�t������F��ɢ-�^!}�t�S��\K�z�Ru��xqϽw`����G6����n���,��e̙=��mm-����S��&c��9h0h��B�{'7,�I�������g�Ը�ĤI��P{�r�'�/��{�T	l�V��g�ɚ�Ϸ��F&-Ql"��&�%�Z�d��B������G"��.�8���	��%)B�dR����.������;����5�/�,���e��|Q��}<NKK��~s���ӱn�:y�}�v��E0���.|^a�`�ou�y}F"����/x�裿q��e���u�ڣh����]���ଢ଼�`�Z����0}R-��w��܁�k?��]�RYE�DҶ{,�9' L�LKl������'��CF�ǟ��h�P�Dɱ�+y�g8\V�ǌa��;�� x��+�C��dU4���ʤ����?��a$U,��i��E�^fFr$]�i[���'�e�J�OW{qR�"'*��x��D"��&��[��~��	 "m�ښ��+����?��q��xoo��0��/���6`����·��>���xw����Ftt@�y�O�d�\���̗K
���8�;�=��Og���_��#bv�ً��:!�{�c0����Ͼ/�"��KUH�, �$sD�������E�]�L�&L@dpf.�͎ƿ���ftv�ǣB1K�0�NAuM�������;�ɗ����!DQ���ۦ�:���@�����0�!y���y!���TL�6���0n��!,;�L|��z��)�A91TS���=�D|�b�I�E�B��.O}�D��K���_´��KG�S��K���A7Jx�g14<  ��YH&ݪղ�H�ϗT�����䳯���SաX��:�c��}w߁�͵ҹ��b�`L:oU��p�����=<��xɬ!9��ء"�QM�����kĥ� �EM[���½�3���8����ǟ�@���
I�U��/ס�2�X���9�u�l�
�T��W�s(@mU5�����;k��g^ �k^�������j���1���_tF����"�hǮ�hm��G�x[w��dX�C�S�5
BR�04z��YXv��8��S'���N��j��Mؾ}+��/J��h�5u����T�PQ��B�3�#��O~|*n�}.$�ò��J�iSh�����]v�(�u�}Q�����$�P"�hG@o��0�6Ӧ7��VǢSi�"�uU�b*K�C����G��Q<��;���vJw����
�it�ŗ���IF���I�0�Ja4n';::*<4n�15���ظ��K��o'&���T�|�	W]w���,9�\JԻ��o^������zDFiy��郓ٞ�8V3���{�U��TA�ɧǳϽ�eǜ,ƩY��ށ^Q����d.��"[�I,0a��ܶS (�U)JTU������#Q��&/`��1�) XQ���^x�M&���lj�
?n��F<���ؿw'
��p��ǈ�pL1��_�bp�鍆��&,X8�*�|�歗��i�Ir�-6��m%�Bǡ��m[���$�H�Z['����h�"�#�A�,h,��s_���n��(P��6����_���-������ $��Tv��l���>���}��������'������x|ޞ�4��4Y������3��`v��E���c.�O@ȿUW��c��v����3���뺭���������ו�u�0�3����~������CWx�����(J�(lF
�5�2��ܚF�������*%ì9e�D3;�����m\�c�/%<�d�F-�T�QHZ��qޟ�4���]2�vX'>Or~�ϋ� �'���搜<�5㸋ρ�|�,�nq�H�'@c5ȅz�HU�R����`-9��B�8� �nP���(v�m[B_�;S*!��!�������z<�Z�5�!�n�i���	��E�&�ŗ�����;�P�gC�h����D.Cm�?:�?p�i�"��� pdtP��i�DFF����JrU���è��G,���[��YSq٥��?3Q��I�ɑ�'`ڑ3t�������Jd�,M���	���ʸ��[�ӽ�K���3BO/�|�j�1D�d\u�]���](kc!�n�*��]6TW����c�*�.�\�@T��Ʉ�[�4L�0O<�����xlݱ_:TvME*CUȃ�� �����P�\n�wY$��c�{�=��/��~��7$9v<7�B(�Pp�eW����� ≨˩+p�u����ˤPQӄ�oz ���=�2�"�72E*k-řC5���[1��	H�Gd�gg��ɂr�t<)�H�g/�}�<���yP�ء�3QQLg����p��x��;���~����b��1�zQRt؜>\u�����m>&Vg���*J7��ꒋp��+��v�ri�)y\x<��Q����g_��w���/ƣ\|9r���W��G��X���z|�?����u[�@>��3d�E�:��������PbD�^�P ���!��V˖.��S&���Wa�V�?}����D�c쎻��\���~��R�#
�g���gM��ç	Xa�7��]H�h�R���V�t�i�Ӝ9�F�)���b"�r�M�4�u�a��T@42�)S����9�u
�Ml�Po���9,T+*k���k����a���4q&�{z�j�J�{�u0��	8F"���?���;v�����*����~lڴ	;�n�xI��`��**q�.���3���P�Ev5ݎ��۱��O�s�>�55b�)�Bg{;�o�*�}��ðkw;
9N�_h^��#���[n�*�aL}=���~��'R\���0i���v�o�݇:�����\L����U�J0�kks3Z뚱u�F��1[.�6x�u����	�gh�-�-���Uu�&z�U8�?���(f1-�ų�:[���ӡb˦��y�t`��_fc��H?�Λ���/�;d��DK����i��Y)�yN��	�&	p�g�Ԗ-����$`�#v�>��#�<q��r����HG���S~~���p��G�9/QUc �]%>=:y<���ʸ����.�p�锌����2���CEH"�>��S������򨫫�\�`0  3�#�ځ��
D"Ql۶�-��������JA��? 1O|<>>;��,�ڵk�X�(���W�3��e455�kkk�L���Z���op��ws�7hO�D}- ��o��������S-��.�T�
	(�t��ˤp,�C��ы�2��d_E�&X��$�:o#9s֤��S�zA?�r�0���+6���嵪U�9��L�"����H��\��<9(ʈ��R����-�K��g���vZa�B~�
bfg�h� ��H��TK�Z���ɫ�2���FQf_��6��3�ј��E6Ckc-N<a%�?����k���#���CR�~�n^�C���
���!�`>_\�'�<.�<�8���sP�&�S�v�%�-�L"ˣPV�a�|��FĲ)�[H���
�����U4T���e��5�~�+��c��)�����i�T�M��\���(�e8i����VT�<6�|%<���صkFG���\?����|F���V\{��X�nl� �c�NC��i��N\u�o�(�Ԝ�'��^i���^=�����#���?<���h,�MCeE #�0cj+���_}�>aT�qDJ��u5���)�����껟�#[�����0a3��u���s�D��I��v:d�y܈�
���A��Å��	o��9B�&$�9Qr��9hnJ�K���P�߿�V.��h�_�	�
u��G*���D]�d�q�q�CϢ�3̀y��d5lz��m��[/Fm�[�I��g�P��/pz}�%QUӈ�o^���Z���792��qI/�)g)9����~�7��ӎ|.�l:���&�X��S��D˔�p�#O���;P)cR.^(�`Ҩz0���,?������� ���u$Ǭ�����Op���ɕ������.�Hb�F6�9s��1�X<g}�tTU��o���K<i��G�ƾ�n�h~[Rd�Y��f����i����QF}}�:-mT�ص=r���ذq+b�R�ܕH�
±A��u�ǳ���J��4�h� l������F#��(��^�nw�����˯�E��%����={��o�^|�tZc���%������%���ҥ�K����k�N�Z�@�8V�z��]E&���W_�o�B<��{�<'���/�e�v�N���c��;w������"�z��(.���=�WG.����V����p�H9���i���/����������2y
��4�`.$#CPL�q��eW�����F)v��R��̫�.h�0�Eo�����-@�G/[��+V��{���U{!������
���&NlB�kǞ=[఑��GttX����v;m%��K"��iq�QK�x=�4�cǉȬYs�3˝��z��	Y8qo��Iгc�N���;hii��=�tr��8�9�ɱ�r�z,Z�@"ո߱1��/��vÖ/_�3fH׋{����y�qu%� �>��TaRL@���whh��T'Z�9�����bpp�x^�_�G5$}��HZ;��h�D2�0����0;;��x"j�!%�K�#���u�eS1��*
�t�lh�S+*��L&�_����G���4A@�T2r~�/Q.���n��97�Nj�r�+z�$�����s���L���'�^����z����NF�(dH'F���$	�D�3�4���Bd���C[ ]%�
��u9�	̨�cw� Hl�2ǝ�I�&�fw"���m!�-k�)Jr9.d��Do>�b2٬��ɇ!��z ��GD΋��F<n�<.����uL&��Z�|���}B>��+����D!1̴T���;�vڤ������
g~�T�\q$j�H�.@Q���C�x]6U����x��ϡ�*��8��He�U��/DP�G��b�"\���������{��p
�x�=Cx����D�;)_6U`t8&uuȃ��J������kuE�{.RU��b09��?�C����t^3�JI��Ԅ<��ظ�3BC�eC2��U�����	_��޲|��`y�/�"|�g�8�S
����0{F3"#�P��H�9������:a
��J�y�p����m�Rt������\�lS'6!����>�$yj��re����<M��H����E�^��� _�չk.©�Q_冊�|�AD#��s;�0�$p�4!�t��\ϻ�:��ʇ�6K�X�y6E%�b)���W_~>V-���C�h�8I��|�QQIBM5���'^��?S��`r�ʹ��s���p����)�L2"�$ռT���e��|ϖ	�q���Wއ�F��������6 %��#8�g���g��Tb�İt�hkۑ��T5�a����?
��>o�5���D,R�ťy�7�A,2����+^(����[�[����ٜx������J-X���A	} ����@C}%�OoÊ��Ċ�G��uY�~_�X�|��z�}�Y�4�W�;=_.�d��-��o�v�~K� �t*.�������o��B,[DCkj��nh�ҡ�a(�ٔ�ёt8P���̡��3\q�q�K��#H \Ƞ��+Y�_r=���CE�LD@$��w��.���ą��pdT���(m�Fsk��;����aw~߾=�	��[oJ���h:)��������Δ�l���hnj���(��&L��pm�tGv�ށl����2)��\�����gT�y,)�<f���b8m䉔�;�{�>��S�|�X���1��8�[����bۗ�"�T�s�(�����yT���B,�|>��*�v��5��TL��#Y�q�X�ѧ��0o���%K������3��HZ�cT�g�Q�e�T�1���wo/7��Kp$�Z4G�mV��p��������9�!�\���wϿ9s��y�$	vq�dO���V-!?��{I�������^�r����q�����ۑ0�����0-����fQd���H$�ɓ'k��Æ7�Wb�X���ʦi��D�MMM�h4Z��r%�ۭ*�RTUU�u��H$�pX�f�Y�4�Ua����`.�/�t��4��m�af.�͖����j9���,��u0ҩ�����<dtt�����7::Xy�@�}Ѣ�[2��$c�1W��?\,�d2Y��\��R(x��i�כ�B_!�}- �@Ҭ~���yg���*�5n<�Rƚ��/GDޜ�ЪA�<��V���k�ѣe�H�&κ
�8�Ovn�(�|`穐�Ř1lIs��9r_�!!B�1^&)'��/�F�e�$�c0�(�If}]t��#R�D���:>Z���D#XcI	
�A 3�G�c�:��#\6Z��'�ɨ'�Ҹ���F.mH�!G#E�.
���n��Chk��Yg��U�.C�9�Ŭ����J%�%O���=��l��m���*F��t�2m��d��sq�Q�����p��0���{�����=�D����v�Ͼ>�@�@��Kx��VB�߆������k�ń�h�L
~��.g#����s�*�7,(����؋e�Fm-�rӥر�+Tׄ�g����mR�2�rh$o����N|��6ؼ(k�d�94�1����A*��+���9�M�붉�$�zev���5B޽���p�}O�l�G�Z��@�����YL���$�r{��(�����ɔ�����/������{�A+P�4T9%���G��X���ԲMƻ�5���(ӚE�₋o�k6��o]F����R9��K��W_�E��Q*�Q��,���0>/�ܞ ��&��G��C�����A��E�O^9k6������ua�>�:��>���qt2��t����}�Sx=�P����L&Kq�<�b����|�18�;*+����ҹ�0����f���s���݁�|��]���#>��Fo�>�Z��fNF��ķ�y�v��r�µ���ض}y�(���*�ny�1E�a�^�&f��������sx�Zf׀��M[�a��=����A%5����MU�Ź�C[k�>������q�o;w�ǚ?E��    IDAT,N[
�8���>�2i�Ixym]���Y�smb��U'R�}t#~������FU���a(΢���^��j�l�h$��8��t�/�9���/�HLx3�MM��bRXrM�C����O��&�P��*�k�A_-*t=.�$؅c��r�gb�S��ۃO?�S�M���a`8�D&��_�+���P���$N\� �\}\vS��јxD�Ƅ`����|��n?��ga����E�`32�Ӡ�<�|)k��1��E��A�ِ7l(��X~�Y�H�'��_������\�L&���a�y���a��?�(+�ǆ�{�c�1��itw��n��g���f��]\�y]+�t���p�G����O��ְc�������"��@�V+UV3bL���r�"�<zM�yW��͢C���� �E�c��M�ʆa�%�(�����*��g�BQ��R~����JA����Z�1�F��(
-���%�T2<���̛�=_��U�}�uEOB3����%��J�0��4VL�PU{QSբnc���mf�^6-e��WL~�M�PP����`M��V*��r<ޞ��(��.�|�_���_��ka�	{�nz����j�;_���譜±d"*&!�[]#ߩV�D���@:ˇ�z���%h`C�]C��<Q9��ŝIYA��P@<��}U�'v���D�_�:o���;�A	x�LH��g:��>.�c�������c�Y,�3=�]�e|V�A��Pȿ"#������nb�iQ��̱T0uR��˅$��+�j�2�:�(�U��q���1
	�#�i���:|�v�NY�\Q�v�	�RI�������ۧ�$>Z6��訌�	�H�K���x��O0���~i�'H�2�\r�k����.O�׍\1�x"&��b	Fr8�7�a4m"^`ڪC�i��U5�\tb�c�ރ��["leE>��"z*@<MRmο�|�� tw�ÉB��n�*-c\�U^w�yX4
�A��n�#MJ\	˂��V�����?��������"W7�"����b�<p�R
F1%]rRt�K����ћ΅�/�=���s?�e'u�p�:J�^v[���V��P�eS�7�^CQ�v'L͋�/�|�W��X �$H���d᳗p���ܩ����B"��
Z�������~��q<��05?
�&�0�Ut̀�V�S��ޛ�Du��h��� �ހ�02������n��܏7��^w3(;�����x��$.<��8���ؿo��K�T�ÔIm2���S�6g1�}�i���s�W6�f�D�\.�㐅S/���S�u�X<�8���������aɓ|����뾇Q(jp�}·*�-�%�&��9TV�1��FF�G.<\̄Iy`��ˡ�(�[�9�zg-�y�(� a܄�~�l%�蜳���C�G���FF����GgWv�:�������<�'NF�P��O�@=b�,t͉B��b�`؃�N9�`�9{%�|f1���^Yi�&�PU[�X��Cz	��;�Rэ��A��e��ڋ�+H$b�C^��-͍�Ƶ�J�-�7�c�8Atww
�%'�~���#7�� ��
l�k�r���g������$0�d��eho��h�1<��_�/8����CEG.��V_/��0QD��Gk�V%�V��֝�q�X�b)���L�Bji��B��B��E���5�p�㨗�i�AŁ��H���O��_}]ޏ��fx=�ń���;�-�B٢�p�\*�0o���<�vA1���Ɖ�����eV���)�7�I6�*<`��8�$��_�fΖ����L�O<���,�ea��]��y�h�"K��r�6�-OP�ry
�|6�t�3��V�PE�r�����ϚnK����T5e�J6��GŐcб�0Ԃ�*y�4�s�i
02Mݰ��&?�M�a�s&r�a:���?���w
r3�L`��p�	c�DM���Ѕ���c l�/��+w������δYw�������3�z�+Wb=�Y	�
�:c�O/	�Y���e&������B�9�xXƑe+���0qV�G!�-�.��q"��r�/������4�ᖉ\�H��1>�؉ �
���(��q�0|x
]�-�gM�jX1q���8p�O�����\~\H�70"��]
MEcm>��|!�ǮX��[�	-5�8S4920wp(�w��_m؃	�恌$7.���P;3	�H�����NƒE��p�Q&��fáC������>�o��!b�,���[���KS1��]�c��:�p����9�>�Ъ�yv������hF�S��(jZ�b4�A]�N|�vm؀�
^�<�������T'��5���2yC�	��y������\!�.r�hzʈ&�a�r����h����=����B����EM}3�u������O�[�C�@Gt��CM��H��շ@-&�q�ɎA���+JwM�ŗ_��>�
��R@X�h���t��J�	]�`��W#�²Cw������fjxTG ����]�w�8�K��͜�L�V���S��0�M:	jU,�o���CC�tQZ��6��>aGɤ;����B.����� �+� -׫�ؑ�������pm��Q���zx\M0L�</�0���b���p�I����]���0��%;��tN��.�CO��_]x5&M��R��M0����.�i�Z���7O�i��$�>�5U�c���������K�ή��+���2�f�՗�n_M؏�Jt-�y�O��'�ļ�3Q*$J��H�(���y�<�����,���dE���!�F?��w��B��߉��C����Aߡat��c��}(6(v7`s�����v&�%����p�\B�/�I��Q�Ob��ñj�B�v��s���i�)]���W�����k�œ�}��~���.|�@W�A��Lhi����7����/_&�tTg!��G�nG%�huvd2R�p�Uòב-��;��|Ua��[�f.^���aE�h��ǣϾ�B�	SuJ��GNǽw^	p�-�124*kU��t�h�X�����c��1ˎ@ׁ]Hu���Yi�JI1"�	,G�.���vYGseeŇHZ��9�PҼx��ȣO�������$>��
K�����[�h��"�w�4R�Y�"LC�LJ�_\��cjI~��� ���T��5��p
B�`]Z��geMX,1���/�	�8���r�'cΜ9�M�t*�����a�9�
�A���G]]�:PPl
;YE��.E)8{As��RI+�l�B�\.�K�r���T,��b���rƤI�ƻR����?}]��a�Yw�#�m���3��O��K��Ŕ���ǎ��aTB�[����b���I�s�Y`H~����i)'�G~����JBL�J&����r|��xҳǛ�.�`���g]v�Q��Jg<�^Ԙ�#Ǳ
��7�7�O��:�^Ƭ3xZXTWV���˶rV����R���/��GUP4����a��>�\*�[uV}c	�Mj�P[KY��A:[����e�>�����0��vg�"��)�?]͡���'�ę�����j���J^��+"�+��w�Gu]�(#����bUQY�d�X���>�`�����#f��~�����N��F�\)/\'*$���d𛋮�ֽ��h����	6?�U�˳ϣ�k��}x��;a1�c�2VD�=�� ��&��<� tWT�eŐ�K�3'��k���[���"�u"9��L.��P�fܽ�Q<�����M�d� Õ3��thy��M�D%���t8]�l4{d��]v-��|to5�`�PK�^΢��x�(��r�҃rmx^h�W��v�jY�0���UW߃?���Y�|�_��F���Q_{�o0eb��^c��K��p �T�M�C�<�'�{�P6�����G>p���MD*�b@��΍��(�{_��ݫǇk�I'����|d+'\j����q�������ס�7&v8�~��7���C���K���N8�H��3D�m�
�Zj���O��˖���/��s��i��m�־�O�cO'��2
y[@
v<.;&Om��Y@"ч�G��駬�&�U*DAͬ�X<��>�~�-h�
dr&Je�m+r[R-n?������MI#t�����ή^���uB�>��`*�5�cY���r:P][�B���
�vv� �®�0N=���8q���14ԇP8�}�{p��wc(�G4^�� 4�#�����_{)jB>ḱ �� ;Z[�$��I[�nB>K~�L����j���ۅknjFS�D�]^d3i1[�p�V32�(����o�]�،�ڏ>�'�|J�C ��n<��N��Cws�5�8f�a��K��a��X���/�q��ã�ױ'�|�[y܃�����ОB�H�Xbj�+�eƪk�%ՋXXp�I�!<�ԋx��'E�O��6a
z������R�j��Hs;�V�� #�D�S�\�XtD
�Q�Y�]�xk�|��T�3� QDf*��&\�qK�QlFXn��s�����<?�DD氻��}��r�3m��M�,�����ɍ�n�;Kb<�u�&~]��_�q��n�5w���l�\�V���%�p�8:��XUD^Lf���̢��Z�Ʊ*�Yv�mK�';Oc�VW���c E��-v.y;���ǅ�T�\����=ݯi�I��⍲����aK�<5$A�cU�8��EF�e��q'��1��c+���W������x�����A�in�8�QŤ�H���"`���-��s&cBs<^�gt��͒��2�>�d^~�m��@��ɝ	U��*t@A"ҋ���X�t�lp��-0�9�����/����:�X��:��iT�6�0�py�hm� �*C��1�	7_�;�۽��j`��\�EU�~oX��������!��(�;{�{zPHK'��k�d��Z@tx@ԡ-Mhkm���0��
�a\|�mX��p�`�N贩ȥEݥ��F	�_C��jD�:P�u�̙Ȍ�ȱ5���hl���>�Ǟ�T'm=��!��D�T����o�Ѿ�Ќ�N�d�9]n��*��C��'��/��}���F@�)o3sp����ߋ���6ՉB�
��k!p��5�}a\}����m�y�!'���Y�CS����o��,�߆��=�Cޡ�c�LPz1(��£O��Ǟ�+t{e�Dz���
͏�pky�s˕�:�n�I*�,e҅t�o�
w��>�t��6a�'�⤂X�C��G?�6�;v	:�H1�봐ˢ:@}?C����kq��Jװ�_�yKFA��*7�j��6�Ǯ8�.��,��opH�;�~Q���-�ߏR���nT�a�v$�I���3�(U�࿾{:�yƉ�Sg�s�����N������xoͧ�fLdr*L�%ݷ�?�Dt����a��46��ȹP��J��O>�ƍ��+شm't��K��&L��\��P]S�M׋������.$��T�bG.��bz���~TV���} U��8��ΔѾ�_-j\ ��im��ߞ+ L����	��0�?Xuuu�1��S��444 �N��pm�&��d�c�Aʚe����q��CY�:���!Q2ǝp�+�oف�;��W����L���M�b��0��z��(f��,���洉�P*����-��@��c��
2 � ,Vf"�N�'��ֿ2�0v�b9,=��6<���x�ٗ��V���k�~	������xE+�XH�a3q�K1p�]��qm�ZN�����w�{�",�jRM8�8�������{���4����^څ/6.([�t���p8\p:�� Y�`���ոP�J@��|.�� ��E@���_�o�֞ohU���i��'�2�C�D� ��rA��խ�C�B�,�pa%�[��\Y1(��n����0Q1>:�w�^T��6cdzM4�*�M�@�M����B��?Dz,�{�v��-&<����8��8,�Y������a�c˟�1����A�u*j�v�l�yk^�Oi$��$��A3�ƚ0�R�L����יWz�����[�x#���bi!A[�^�+b�f�\���8:��1y�$T��0��۵���Oqұ��s��q�����{k�b�ރ������1� �Yuu��pV�X���)&��q�e�@��=�2i�,�%#M7�"g���@,Qy:Sp�:=��D��ŅgS[e�-7]��h��0z'1��d��sE����!\v��b�A�^�f��$�i6�p:\s�yhm�@t��0�
ټ��T��.Z&MÝ���Ͼ�Y/ �b	B�T�5�u��0��s	�q\@�벢Z��
��������}�y�/{D��8��jAw�u%��y����e���B��aE��_����t�����O�03��E)=�뮹+W�Fw�^T�*Ċ�Tf��Dv�n_5^~�<��K���	z���S3������Au��b~�.�P8_%�����`wye��g{�q5K��\Σh�P��eBG����pܪ�<�p�F�y��}�<��E��mg;������߀l��&���F�e�M>^c}������Ӱp��{N�i6#G�,��1t���?<�X� U��D����㵣�~_G?��٘2�	5�bq��і�\�����i��'_l����O�s��K�j�>̚ނ���ƌ�M8�9�����-��e�6Iغs�9O�������@%�=7�C�@�vMF���@�^����S�{���W?�i����!x~�:�t����x�K�����O��K��	*��ae���!�̄�&��n޸Ih�ѥ�R<I?8��`V���ǬJ�Dj�$���p^Q��bVXP2�$�C4k
�.]�������x��q�'��RSڂx⑻t�������!lٶ	��0��µ�A�	��l"��ν��w �ČAXZ�(�a�RV�H�7U�
L����8���^x�M���[8x�3g��a3��Ϳ�A���$c|�Yr�8�4=�q��������� ؍��k��xt,��b M
�*��L !��"��Й�e��u��tr�1�jxSL�-�q�q�q�9n�DW{�#���
���W����(��n����ށ��i@���������5V%M̂\l��q���$uAFO�1��9yB�mƫ�Չ���5�	a���;���p�0������t�YYeBp���	�m��VO�E�xS�]��D�_}1΋�<��.��E��?���?e�6��=~{� xlza�Tyrl����U��eG6���JW^q!j�}Е�Xl�j��&�H��ӎH"���a��ϯI�˔�#�7�m�n���ztx�z;���o��~����"�R�t^x6mE<�,8?b�^{�o���_�'�l��7���ϱc˗h߿7��;�غ�[d�P,g�i*�B2�*Q*���_]��H�p�lJ<;��됏Fa����uKEJ�?;��/��b��7�#�K���1��5�K*[�v`�2���_���'c�i���,�$�@�c�������S~vW�&�y��)��QP���~�B���٤�֜n�����`-���N|�� ��F�K�׎ff�#�#�p��[n����t�UΗ��z/M�	�T5������'۠{�)h�X6E�_��2�Vą��K�������":2�l1U+Kު�@E����1V��9������Q>����2����r4pT��da����gw��-�`w��}��.��:��M�<�htT��N=���8����D���,�n%g�h�	�d>�2�棍x��7��� K��2�R1�\:���C ��c���8l��hO��rI�։TC�#ؽ� �~�e���x�����k$E<1 ���������`ڤ�"�Pʚx!�
��8�3�M;�㍷?B�t�H�+"m��    IDAT;�\5�Y�=:��h�q$�OmƼ���
ɚ�Mk�3i��r#����S9��J�ME����ʆ�NE��F�L�14B���ӏ?�2b��/����:y#�{���]�;�+�X��_7|n'V.[�K�CxșEI8\�]��;lmh��9K�|N2
�Ο/B�����ip26O�|Z|���e����n,ޅ����D������$F�س�}�x����k��'t	�*���{��P�2�ߡb4:"�8���ϔ��b�W�&~��g@+��Fl��e�ͼ��3�f�V�i��"2BGQ�4��c�QǊ%�o��/����aL�83g�����!$�d
eI8��{��iÃ܅���"6o���P�EY���rgQA�[v��Y
y�ұ��1��q�>C��  o#�o�W�~g'��8�"8�d�r�J1U�E�ǽ3_0n���o����r��_�	�����i�� |�ӯݼ�=vB�^N���K@�,�7�Q�s,iR.^��i�i�h�L�Hv���1�3#W�#E0ˉ�9JGl�I�:�-��PH�Ęy�Igv����bQ�,9���(--�;��rۡ�Q��������;(|\�;k1��@i��c`R��T��t�+ ���?:f�RK��9U���WG<j�
�*I�
�eM"����O�᳧K��v�H਑�0n��T�l/��:6mމPE�ڰc�NL�2I�����l�\���E1�����Q���ۅl��_{�;:A��(`ǂ�me,^8]��p�5#:҇��)��2؍ �-�Ӷ�S	��9�^��;PP�x=>$"Q���]���p�u�Jn$��DZ ��n��R��r��V�w�߀�P���BHwjv��s%N��o��v2�m{b��۶ms�	'�&���Ķ���^��߰U�oO�S}�������J��/E���܌�����Pt{X��
�WdЮ��9�f�p�rx�Wm�Zb�Y�-��D�$��d�����)��	o��u����>N����LA�o]��]M�\��2�����xA��{i1o��ny��B��a��kB��q�D~��Hh�K�]<L-���,4EW�1C��B&Q^~
�8KQ�P&@�ڏ�	��<l��W��.��Ûo�-�Ʒyb�w��O{�lҌj��pҕ���^�1	I���8cC�U���^Ɋ�)����vtߏ���T��V^p^��C�_$��j�]�J|�C/��qv{���˥)����h���+�m����w2W��S�$А/�9T��ی���B�R"�ӱ�ϥؿ���S�;���3��cۏ��;G�J��y�e��w	��p����	������u��Gp���[{�ĝ�g�ܵ�
�L�N� 8��g3���F3\v/�I�9W��t���_Uer�,�7&Cf�Q�SPqn̦������k�>�{gEcq���QE^��~��T5v��g�Cr���+�����;>KY�~��fԒ�%�6mZ�;������Q�=FaN�-OT�n�Zȗ'E�[h�}B�붴����þ����u�곲 L%(�g�8s�#s9ҥ���;�ެ>F�8'�k����fh������2���E�.Eƨ�q7ҥ���(P�s���䍫&�_�R��sWr�l�?Qv]����8grZ��zޣJ����5�,!�O����-��t=�t���\\���$Ǔ�3�TQٺL�[�p#��>Y\��	n�
8G�/��������8�m�7�c���SV/A�{2�6?r	��H�kM��`y:��%���~���+��������F����q�zk���{��֏F�V�3-�}_�x���j8	x���S�U�L�p�[�����>i�3���1������d&vCAH��g�.���K��$ȕ��Ӂ�5&����4v8��B#�oE��8�Cy�+`�4QW��.н�+�D����j1��a�ipW�C7�'"c��B��D$dE3�H���f�7 s��M@"M����en�~��z���p��[�jYc���I��yY��y���x�s��4���+�O�OYL��˶z�󤦦n/ߘX=���f���Y�F�iںhӜ�U�z��
 �Dm����W.�Z�i�x�x�v��{�L+gp/-�n&������M�f��:�(�>\;���J�ݫ86���vt_�H?����6�������C�'�aZ�XH����Ҍ�|��t�t��MRUQ19��8��ӟN���p�f��&��Zɹ�UM98\R��s+�[Ѫp����׀� �U�1��I�޴��O�<!�xp�e[S�G���$&�aR���������R?�NV�` �"N����k����M�ݠ�s� �`��bf�NS�/� rg�:{埛�KYF(HNk�G�Ǉ�s����z+���[��̻����F��	I���~�!��*��_�	3��Q�%�g ���Dꉹ�x{�+�9�y����l8R����C��o��x�cSA�q9y9����m�4��/�ɔ���=�����$~����LK�w������ �����Vi��9�UcT'��N��s��c��G���G�/e\�o�_����Kɢۡ�i��]?߿��m�Z�w��h�82gh������z�:�g�� ͸��˔��-�ı��Q�lO��7�qNQg�W��Re9��:�g��������*6�~��<»�&�ɜx\����XV�s|�Wʞ*�L�"���$`���pz
���*��/f��ܭ��#WT��ϝ��&���3m��ǝ-9�Q:H�B��R�?wآ�U�fTm^o;�1��o��B�N�v<5T�Չ(�t���{!�s9213�ճw���I��E[���9-���>�x�=�w����y'y�����~@!Qp�6W����Xސ�z~Q�YL$�xx�C�W;jU"}߁[}<����;��ؤZ,	g����w�Ν�ζ�IJ��	i[��O�Ҷ�t�z;��o��Y��)�"��ރ�~[�_��>�w
�e��8H׸'��(����L��?�I�.WK��)LF�"b�����2��U+��:E �^B���#�Ea�ߧX�e�N�z���q\<D�>	=�s�rgZ��ڨ,�~�H�n�~<�|2}|���-3��GR�P6-w"��"�R	"7t~�$z�ܿ��XQ:(�����7�_����2�J(B���u����]8/[8�����`�����^y��QL�}�\��s�����q��όަd��ND���*[��S�p�2�?+QOt�_pYp
��m'���n?��6$\F��Om4�*|��p���=(�#�mZ�ƽlZʸ�����d�wO�"K��<�N�f\�΅#�W�@#r�Z��M�̦��5�?;(��m�^١����6����-��_p��n�Hʸ��E��S���^�XI&ǋ1b����N_�+5�,� ȘH��������s�c�'B��c�|L�s�$�?8�v�K/�9'�?����&e&�!���t�Vy���(Ιq�}�Z��-J6*�g�ig����j��Ԓ����|:�l�\��v�i�û��5����\��4�3�j~(J�Q:|�;X7m-qtن:��"�>R_\�Ϗ|�5^+��(JHVeC�׀eӟ|��̊�Ș��z�v�����k������x��L	�<�v<m�Y;x��4)PY�A��rJKI��]���XW���D�`>��L�'S�Cl������������*�fph�0S��oJ{{�M΂��x��I�T8��E{<v'p�yi����r�0�A��'D�c{��>�Ǘ��})��ÀrI��)�@m���/ci��I	����!���ysF<�X�x��į�M��3� ��
u�g�A3�}�W�J�vO���9�b8�س�BN��x�c�����<����mJ<�ZiŌo?T)��;:W�'c��ǆ"o$��sM��#u��B#=}��XS��ܩ��K�}��l�lh�_�Et��+��%���+���* ��.Z�0#]��	6gus�<�w��{�)��E�麗eN�Z�˩����� ��G�.��1E��:>�Ip�z2OÅQ�F~aWP"��p��O�_4J�)��[-��N��}�����}������/7_�U�L�md��ty~ ��i�侊���"�&�"��Y`�_�9��A��l�*�\��.���?���sN��p��y�v1��J :p�?�V�ڋ��<���,��=Z�q���b͙����w���V�w����5��r5[!�B���4j��s���s��W�ǧrR_
�o1�ȩ{�3��]8
�ވ19�W��@V}��-R\:W�"���}��1o ���zο�xo��7��p�ꫢa��z��^}]�f����|z��v5��� H�y�a��y3!,Ϛ���vag�A�I���������qU�U����F��D��'��3�e�h��`��mҾ넂CY�\�X�?^�&�[�x~��v<��}}��V�z��	��3l��M�6'�*��5X�O���i�����L�'mF܃�2q�b����<�O���j�Q�x\ƛ#^�{��gnAv"_X����گ�Q������*p��oȴ*[����xGa�1ӡB�'�®t/���2�;.	_%��SD!��(t�p�azlZ)<�ڈxY��fev�{	��궉ٳ�B��a��~��DaU��`�~����]����� Z>�w��t�CG��,����A1���fħ�hARp4��H�R��hcY	�۷i6��W�<ϐ��08}:��@�\�u�8B�|+����0���|U;�׼M�x%��� �`#�w���ч�$ەu�(��������8n~�ptyE���̒v�#V	=�)�B�Ŀ��@�o�!!�55����X4
��8�*��ۢ7o�S�tsB�a�Z���] zt�Jb������8��մ�F�4��,Y����E!t�k���������+���1��p��-����\����`��x�[ԫ������%>>el�XEl�gQ��� �JB�|OD�i��P���䕉��C��#?�E�󬗗	�E\b� p	l��i��o-�Tٖ��M�1	&F@D�w�IAؚ��k�}N��F<&�iz{��>�A��Z�Ah��~=	��¿��yb�$�%�8��8[�g��7���M���y�S'��m���`�����j��
����q�=�*	��`���i�
�_DEHG�rm��<�$"7σ���0����z��A��D��j��� ��������PzyٳLp9��������}�ᇨ�xSl��h�m0B8d!��
���Z��Dw�p B�F�=:.?SV����<��?�fP�4Z.�Ґ��G���֟6��'��4��mmy.,7+j0��ϻ�[�u�f���"]�� Wx�~��X��V�W����u�,��l��Th��u��=����}���K�Q�jU�e��o��~?��vщ�;��%u һ;7�6��'�s9BD�h���׺�߀Z�h� ч�SI*�Ck!�F���#V�a��"��;�\-�Bh���՗�k-�9��s0�8;���{�����LJ�6���о-��x)�7�QM���*o��{�eYF��QXiB�I����ż_ �jJYI�Z��^'�iA���m�+�#��MC�ާ�����0l��j=H�Wz�0���$g�l,-�4o���۶�s��x�8v�'���=�CW�ﴧ��k����Y�}����W~�9}U,����:ytY��23�h�6��x�2��G���ք����W��^f}���� i�W����K����X�3��ln�=��&�md`Y?�0��o( ¶{E�mo[W��`���3�/���	��2����?�4^���n�Q�WH�	����K)"�D�Ʈ`B�4gŇ�O���xN�k��X4r���~�k]��'�:a�T�E]�t���q*� (V��޻�֎� b��}\��?�[��a�����6����$�Mf�]�K ����c~�W�=�4�ţ�]L��3�EUQ�LnY��s�Q=Y��E�N0��6�� �R�B�y�;����؝����anCS�>�f~��ʜ�y��]��%��R�%����D�5��9;�~��M�(�f?�@�Lw��ٺ������!L�G@ f��E�Mjo�P�Z"���I'�8�+�����&hzV���9� ���r$�-�RQ"�an##�Cw���.��u�t���i�D��	�L��!��ܦ��t���}>��n�g@.�B������]@�c�8�v����ЎR4s7^Х5Q��,}:�}3���Q�U�N�?��-H�Uo��\ί�8O(J!��h�8��T��y^y�ڐqV�*$_o8#�٦�D�5yn�e�h��'�viŇ�p�ߤ���}Gs��г���LBn�AYIW��ic��l9�R<_�	ZeD�M�!�Qf��5���v�p/�^'ˢ��=_�H���a�_I��I��#���i#Ev���;�GZ��3�C�#R�����
����>���|���)�#��N��5���x±i)�o�_sOt���C�ER��5��e���e��w&�b_���#�Ѻ�����}���p����ee��D��"���Aw{����I����Z�-,�=���ĩ��3���z�(Ohc5jƎ}.c��O����������O�d=a�\�զ8nH�<�b �A��Mf���G}W�<b��$��5��7�u����'�\y֜�>m�/�y4��x�ч&K����C98�8Ifz�q����5��$�3���}HUa	a�F���d��氘V��	sP�����%�k8���z0A�i�Vs�{L���ڙ�JIszq��8����TZ��W�Q{�_X6tQA0T}�=��3�f�����P����AMN��+!(,P���A��p3 ��j�]6q���I����K�g��ڔ�vfw�����%�^�ų�c9�Q�iK%��䔻w��<��r�b{M{�.��pG�D�:G~+� ;}�Ϯ���� �zV�����r]Ze����"E�}!l�KYH���0d�q�w�F"�.�n}�V�0���4�������@�;�<��$����ߚ�^�PF�/��l><�t�i��y����A�0�J�ɀP��k�ׂ{w#^����tvuHMY�^q�`�[nBJ氶1�a����mP�}�Y	��f���\G��p6Z=G���9�+�BH�*b�QƯBq�;T���9ԃ�����	d��\n<��}v���~O%���U(�$vH��:>�L�MQ� f2� 0fr���q�+��V�ѽ�%7� z����7Dw���x}�J���>y�R��k�KV���.����a>{��~�AA~�u-�|��7�y���6��wr}� ��r�n�X ���ט��_ct�}��C{������>77[>��z��;�6 �_�<u�jɸ�C�3ؓ��x��W/�4i	���p�ο�OJ�o�赆]�HH���/&&��-k@������Aƍ�vD�P��R�\n�I0�BnyH��)�J5����YgK�t#��wy�X�$6�rp%���:��͍r{v��԰Դ[��9��E-���?X��9m��B�wb�>!�H�e�!�~�?��+y�����O�C*�Vd�A�p��tY� G��vd�pAg��ϴ��]t��&Y���Wc�M^Xx�蛌�@���9
9�S��CW(�#�ݞ�2pP��A;aJ&˰� ��z�����;H��YaId���Ƿ�ݲ�p�h���VaeҎ����_��D�&��o����m�A8(̷ljj��V.��y�n�J�BKs1��<�AҘJ�O桬(l����vu���J*S���Ê��)�KܕB��/p��緰��w>�D� 59�4��������rw����Cs#o�1�D$��s|�Cۣ�-�.b�Q�r�1�yQ	b�ߍS��뾋��;���}���r�����(?����t�?T5�凚]�5GN�)P(53��&l�Ȱ��M^��ߦ˽��#�q��_�Ƿ���m#�ִƱ�;�8� ��WJ,&�ר|\aB�_#$ g�Y�A )4PZ�<>�( ���R�G�m��y�yr� ������犸�W��B�  .��� Z�� �T�t�v-@���~���#b���^T.�����qEb����bb����#/��.?N�Ŧ�V�*F���{<.��1Hu�[���N>f�Y�T� ����bW���.s^se�� �j���c� ��� �2���X��cp�r���ϓ�	�H�ӗZR���������l=�_`߀��cVVR�v�\re]\؂5&�^(p�#�܉�������6 ��Js���r[��r>|�d���uF���/O>��S!�'=)�v��~-��$�&&q �-
�D R��b 3���5�}����I�|��q��A���.,�}�=;�v��5E���>d�dE�UN���U<So�Iɯ���ǽ�Ij2剂Y��UA?'��j��
����Տ�9�QkK��׏�
#��[�X'�|B�틧�:���D�Ս�����}�R�>���s���?x�7ZN��'��-���q 7�����Qi`)��,ǟ�?�w���98a��[�bB2C^�x��dk�j�|[7�����VV��Ky; f��|G��*x;7ɡZ�"�/S��17WCL2��QԖ.����o�R�<Ju,�Pv��D�y��;�pb��c{��v�O�D�é�[E��	��9��~(.j/�{�%OI�ɻ�����7�s��a����J����o���׻z�l��ž��.XS���΀Q�R Y�4�@ӟ�{&�[�Wx� ]�^mG�Q�ޛ:� �'�7Ϻ�<{����f[���&c%U�>zV��N�AX���b�����f͕U/�궸Y���P}���!���z�w�#������F�e��ԇ'$?� ��۟�v#� ��PB1p��.�n@Y��E��8BTP[s����慼�)c��겦 z�#_3HV�����[A$�r-w��a�H�sY��,u�� �E^�8����f_�\2w~���t�i#��-�VvΨ�*3��l�(��T<���6�Gy��K���m���� �`�:v�Rɴ�_��˺bчhf�P'���c��:�ʳ�����XL�+!�n�pu��!D?�x��[�2 ���t���1�(���j���S�JL�+\�&]"�$J�P�[.\D�����d�����3�� �'2��M�><N��31<�����'�6s ���� �$�L�ŝwKK��'j�RA���I�RpT��#�(6� s#��0qb��3���U�W&s���@`�H:�#T�7RKW� i�[�CF�N�{�7�E�S6��4��]��-42+$Ў�h����.>f:�s�E�m�tÛ�Q/f`L難i�8��nP�yd4�#^=Q����6=�
�'�H� t��X�h���v�F~��#�8t�������ӎ�o�m;RI��2��fR�H̠'aE뗍!�9&y�#9p��pY�+6͝�8��J[[g�]:�: 2=�q-"�C¤&�`�ɡ��}E�NÞ:Y�}=r{P��s��Q2��X�8�Trs�7�T��5���Y2bg34cJ�8�s��ߖe����4��B���z�Ph%�4�4��F�H xi7&�p���K�s�_`!&���>dc(I�'�`U���k�9�<��^n��£����9��b��
y�:�l7����`
k'���i(t{"�=3S@'�N�PO�Kr�S�u�_��+���	�$3�PB��﷞R�xRP1�1e��+;I�
D)��6�a�:7>���hǞ]�{�lo;BI��\�VW[�d��"-٬g��V0�Ԟ�L�(�"��lY��L7m)#S�N@�Ep4�1G��k�lw�d���oCF
�0�,��}!�~\�X~�X����YS���t�*����kOj�:t�>1}c��a�/�fi�)�X��������0�	
2��t�4k|����湁ӽ���B.KԖ��e?�Ҭorh���)#6��Jv�E��,����Vc��Akp�QɆ��3��P���Q�٩aiZǲI%Y$!��!�c�!��ϷlH��?�O��-P���3 8��+/mM{�S��,q�ui}T3��][�+K��g�_�d
tM�)Z	6=�#�����?�s�,�U�;K�<]Y�S!�����$*�Y��l��v���s�rs<�����?�'�-��rF�GGG��t������fXh��8�k;;��������z|��g���6Q�3IFx@�_�U;'�[gV����ju~WA�����-����� �F/#��.*��&&L/�ʮ?��(&4ȵbhrLzB����=p�l��Nj��!PF5#E�@qD3/�В႐�pp�XY��:������3w �L#C~���b���� bX�Qh���������Z!XH;g�X�RF��s>�[��@%��|��4��̫��f�~&��f��Nd��Y�#[:|�A�%}�N�=;��%���;�7��ʆ��}!އ�c�Gk��O;�V<,(*y{O�Q| h���%���������,��]xo�!���%P��<K2�25�����m �Q��)~i��)7��S�	��aQ��������P)�<���7�Z���������wAcm�*�ۆ�&F�*�M�r�/�p.R<~���q����P4(��~�eC} �xl�S���+�Nt�����qV�Щ���Vv��4樠�5���;�_��j��{/UD�6�Ť/�)oL��]/�FRH�G Bc���X�W�fѧ��-�ג�_(�*�����w�|/�&�zǅ "I�p��]�fz���s�����g����q�6J�ڴL|�n�*"0��sX�c#q�)�(C�.�ʁ�r����O��0O\6�Vݾ(6��6�x30��y׉G�8�Kt�}�q�$^�''+f=����3��:��}'�>�p�����ޝ�ƅPM"�/.��>'��g�x�xf��.#�C=("N��,�q��X-)��DF�e�'��ea)��)("��!�������$Lz��=�׵�G{I9�b)�����E��
k�_���	e-S�C��^����P���IU�:�6�Xo��]ܪ*�8�Ya����wB��"���@}(�m=��M��W�A�@7��`׮,7�Ù��r_�2���#jg2M]��%4��.=�l|�VU���e����v4"qh�Z9�����1U��R3��B���I��8B�<H]!�/��u��Z�>/�x��O�l�\���gY�x�"dҜ꾭1�-�̉��q
*�1u]�i�ix}]�"28�Ά�zi��92�Rx {�ڪl6M���vZ6������\E	�4u��Ѽ��3-�����ص\�C3��a�맢���d����n��Hm}X�ɵЕh�aVLu�}�NW�g(�<=ul�3bE�@ �EB���O.��Y\Kw���kZ��	MO:�|�u�LĐ�['�f�^��ǎҥ��-Oں�S���X�A��К�D�0��}e�J-ʖg�A�g���$�Nܺ1l-
��3��QĤ���������ͪj^����o��zӡr�sx`j�>�u���t�ơ��O~��۾/�vLD����ݙ#�a�� _�X�McL�tS��mQ��]��Z�~� E
k�]İ��63s��ў��W8n�yQ5z�>V !$��ތ�o�a��a�پk��L��=��0�ʎ�σZ_G�`�a��W�E�ʷʠ���3_�#x�*��H�1O]ԃ]4���@�!�����x���-	a�bO\CcjQ�ij��<�&QK�gH�\N�|���M��Ar#K����vA0 $��\�N_�Jj��Nĉ=�W��X9� p��j�.dg<͓􆹚�=M%�@�^;����D��h=%q1�Mx¯c��}[6��zR�쇇�c�'ka�*�_����m��%�C��>�<�~u/.�B<�Z�e;@�</� �m*?�)�}Jt�Sb�JI�H�.���_c�B��;��a�����b{�����e�:�%k��#��G��*i�hˆv���`�8��?�V���my�����qGt��S}˃�J�HN��+�}�
g]�֢2uQ�^FV:�gV��5鋶�P)uo�D���e�A�����F�HE,��㗝���2g�l�rI�!���0=�3�����nJc�������1�s]:���	���ϯ�\�>���D�c-�� ������ȯQT�����/�j�U�����ite��I!CuM�:Et��4[l����5�4q�y��R)�|u�i��tS�I�Lq�Ak7MM�q�&��\�?ќ���T1Q�d�e��������d�m��JI�!`t��X�<������|��c��"��D�%�����0�m��?)��A�i��ZXsA�͉�G�����t�w��H���aS�����ڎ����i��a�K �������	�.J�+w Ic�M�hj9Pj��l��(���N����d�5���ߗgm��� 7�fY�=�(bM�>K���s�)�2�y�$�g��B���)hZxq=D�J�,Ȁ�5��h� �Q�<[�$�2"�j�| [�%^E� � S,#��;�E�qυ�h��c����R�@Q�WϞoA��˸�m���V'�0�I�n!�Qo���A��@���9:���C�;��9�#�:�4`�}��s���R�Ԓ&v�;���*t��%oY���,�����S�e�As)�����48ɀ��A���������71�PVe������:����Y|��>�j�H�^�c���>(O���0N+D����AB0�#�pv5'- �d&#���?�W�H�n���m���.Y�`��o����>���	�X�m�׆�bm�I�$Տ4M��h�����7�ax��W��︫m8:a�����ih[x5��p�`��'�3y�P�$�pE�(1�~3��00���	�`��W;5ͥ]���t�!���K'rfb�}�	-zk��e�6R���B`1B���s��$0 	iHϺy��c�Y�ɿ2���[OH��E�{%	�QP�f+Ot�����ۧ	5�cPC��r��y�q�O%7��2���K&�x����ŊR���uB��:r��Ư7�=s��K���#��jo���a�@��-XS�j�~�1�����r�:v�*��>�%��s\����RS�T�"�|�>��-|�:e�)�C�A���2�S����&��E
˰S��� ���&�������\�~���K��HՁP��"���d�p*��h�����B�}d�
ԡiK�; Քq��m�C�P���\w�>��N�u�ʫ�>6uBX�?�Ǻ�-��6W�6��{h��Y7�mRY� 4�N+��#I���M�Y~DJ�岓ʬC�&��>�,z���J`t-�F{���w��{>�0���aD �bU=� �g� ?@DM3��Q3p��
Zd�!C����/��4��tB<	�dsu#�3}&'5}^�k����_ؕ~r��f�pv�H@;|`ڏ�a]�Һ��x�����(;V"�*"f=��2V�;n 
;U<j� �Yx��IɌ�h�7��5�7@뻔Xei������ϯh�+�
&�\+M�b+V�tS�X�²��$6����$yTE1�&�Xil�<�$�c���jX�bͰ)15<]=Z��j��D|r�!�h�Kj{�F:,hw�y븖4��&E���4����-I@��6\x΃B���:<b
�����6�L���^zݸ`�~����P'J������}
�l��)�Դ$FF�%�@�2�~�$�WК�(:��]3b�����8kA�Cc���+��`���7±>��2̐zb����*���;ߘhF֏>��LN��6�]���/o�,�wSm
0��~�BĽ�E��q�P�'��V�C=&K���q��[p&V;|�` :�\*h,5�ث.�[<ӥH�`^}�x��uc��j��GM���jH��9Q$� j[�� 7�h��i����pQkd�dN�(���MTW���t�1!�,���L�;A�vV�N�QJբ(��!቟�lJ.��z��6�Őbrs ��I�dW#rKsW�K�$�c�x���.I�Tj78jV�i4�5`��Q�f��4r[��b���u4�I�5?!���7���=,�'m�ؽ!�:؎�.V���vTN�,O-j���#�N�q�j�v^h�j��EN'�Bs� �j���]%��)���!L8!��ƖH�IY�@�����}��-jA��=��Wo%����*��ej��.�Tܼ�e�������ƞ3��Q4��Fݚ�z\R���:Ö��.L���\3
�)]�Rw\\����1V!'�ל꞉S�5}.]��,�f�֟�+�M>�C�J)�{� k"/���@p��lNUV͐�<R��k����V�G7r�k$��"_M*�tcM��P�N���X$�.D5i�z���r�X
�A0#��.>7��k(BE�<�1E��gn���i����K"nȼ�*d��n���
��%�r͟	�%]BFb|f�AB��PSM��Na�>�[��Iٝ���Hp�-��(�xRcj:�����/�V���K�`+7��F����S�$ʖ<���?3��Γ|f�:�a�ْ<\r��H YH�a����N=[pf�=��Zo@�t׌3�g��t��B�����g+Ls���ʎ�u��TB�F]|�����r��� �V	�C�Az��Av��؏i$��!D�b�pزyM���|��|��]�����Rfd�V��h���i)f�>��|/���=?�`����f��i��o��y�d�4�徯#M
}�<����m�$ܱbi�<���]:)�-���F��K��	��g?��<���M�$8al�9����0?��3v$�L�Dm�%��N��+)g)�3s����~-��L����E�/���l�}���m�����=Xi�o�_U������u�:��_��Y�/܌��(�4�M�KNJY�N�� PK   ��W������ �� /   images/dabb1173-90ac-46dc-83f0-6b94d38ee5f8.png\�sp%L�-�9�1��<�mN�	&�1�3��;��m۶Nl�}�V�w��ѫ�Vu���]{��U;BEI�	UVFB����� ��"�����&-Q3E|A!+!��ip��M�����Y��oQ��ǏTSX�U��C�!8[#��t�Qh�;s8|V�`6�>h8�������h��K����/����9T�t{u�c?�����=��'Ιwc8_����=ӫ(t�HY��_��#�<�zfLo(�L'�R�u��2���P�Y�n��T�\P�`��.�_�0RFH3_0�{�bz� �'��F�����"_�-�i��� ��?��Q6�)��PޡQ���-��9J��w��<}q�ǩVÄ� .��oS܃�
�����N�1�]�5^tgLb�M2��ፔ�����y�T%�I<�Õ!CW5xt���r��"B�:�$�,2�qs���6-�E񱉇�D!&,!3|"�7��P� YV]���� DJ��?�5�u;�!D�*�uA��Ct]�7χ�#�M�L�,��R6R��g�*�|.��~�ݟJ�^S�i����Q�~3�v�y��ص�<";���uW2PU	+ R���`����#A�#�x4U5a"��a4D,1KD4aCj�#���*"U��"�kf!P昷_"�b0�Ex$�0A*��Pe5�H<9�c)����Z?B97��a��3�8��jr�nƺ�˚ �xt2�p�� :(�px� W�Z���#b����5a:�����e��tlܜhÇ��1�֬>#�I�Y�����XS��"����0�d�1�"Q�[e��I�س�<��a���I	�1�Ԝ����"�"�o���E�;J����b�R��Lx�j�
�u�5$?��%Q@%�qp��ќ�� ػ5�I̈|�Nrz�|�'$�!{F�"co)ub�ɷ�b�֫ %�?L�,��D(����}��}l���~x�`�E>��������_$��(�8$���Y�ú��<�ƳؠN9J��w�55I�
)yO�gQ�Z0��b~7�5�Z@Um����;��<'�O�Z����ۡ�@U;��镉��m�J�8y��1�2~	��_�V����Z$�YTu���>�r�T�P�e���NIth��8�T3ݘj�׮����08���*6��!v+R]�O��� 
�px��p���[u��8�[�~�
�t�����I!a�h��s���w �� �D�\�~	�EH�\1+� ���#�*4�z�@�pgf� ��	}b+W�A�م}Z��3��&�VK)!YF�D���.�,�_fM����@�=��2�O	 VF�_��Ǧ��t�(�C�Z#��;#�",���1�-	$����#��T0�a��!YG�1<��<b�i8C�|K�u]`@	|$��&�������fLo\�&&��oJ���j��!��(~E �e���8�'�|-BAC�Uy4��B�gB�:���)(�m�N�D��J�D�Z���d�G���Y8��Zh$���J�l�Tu#���!t���2�d�nN�0�Ua�V�����>BP���I)�g�ZBl���h�IR�L~��ò��A���T��q%���;�n�A^��
�3��|��	�q�@�!�7��|*v��x�A���
z���&�,_��9H�,�L��*Բ�����<��8 S�ȵ�5�qݍ���*���Ο�O E���'4�Z���?<qs�g��A(z�ۧ��m=����Qf}�O�Rl3�Q%�ƧHW�ؾVg�%���E%�t0C����{�~�e�w"I}A���#�P:���'tz�%Eb�ݳYi�n���,�,cDק�N��\D���������q��ښ����6:Ե%�����=�ɹV�������Up@6q�ܷ�z �9�!���������}��+`(~�`�
�Ƶ,"�8׈��t儢��Pӣ_�	�N�)m��u.�KaQ_,��ؔ�*����@HQ��A)�2���9b�ϠŃ,� Zcր��g@�Ԍ����e	H�,�mw)Λ�*��MG[�m	9,\�?�lm�S�de7��W-V�4��L��2%D��5Wh���߽�z)S�24�&L�5�6�E0�\d�o��L�8�9$�9�����q9��:ؖ�l<�ps&7D��7/1H��y���� �"/�"��
�O���u�a�t
+��@#�L�H?�D�V��PBXB�U�PSBׇ,����H.��u-�SAh�vtV�����ht�Sj���JNjTp8�;T�g��� ���-+
⦍��Y(F*��Swa�l~d^��qqU�1�����ҋ�� �-3��֣�#�P��� �����ah�
����Tpz�̊B�*�s*��M�� .E�u�6(uTΕ��q璽�BIz��*"8u�
���!��>�����ݓ��LU3G�7]Lz��	���xI+�Y���ID�}� F
�g�$	r1�D�<�4�AZ�*?���`�Z���q�7Av�/�a{
�>��q2ӹ�d�.�����w#�O�'�ϳ�'����&fq߃��FhP��E=f\@5��������*["�08e�F�?��|�E��Y~� �����&��]M�{�6J
VZ�.�)����+;�`i%�SL���n��<��	5�:��
+Q@�i�R8;�+$"�I0K����]nv�'��
�o����£�(N�h@����x��J�qs�-VjVWö꣙Pz��9.�V��X�:~n^]���;݄���1�v@�/:�H�^4��H��ՙ�Md�a{l��OgE�2@�'�ik�f9]��95\�W��o���b��!­�#���O�u�@�uo:�G"�*�U������H��>>ѷم���|[�霏b�C�kS����8���tu#s����i��\�<�u��S�^������cr/sCo|�z��h�_���6�z[X0�1�� z��t�-�L���P��ƠL��"��)'£�٠�E� ��WK��&�n9��,���� ��`��ʀ����d	�t)�2%���&^��UD�Y�u�9+'/��imk���&a���ϱ��Lp�����-O'��ߘP�Uc��;�84�*��0�%[����(��"�f��[���Ts� ver�3��I2�٠̻�'f(?$$��9ZQ��
�*E�/so�2��V]fz��|R|$�~4�u�?z��R!��.s�h��b��b}ъ�'�}~8��4�0���T�u�%l�wn!]fmV	����ܻ�L���#����=;����BrD���Y W�T�퐍bĂ,�����Qb�! �K�m�7PG��V���U|��u{A!/��.� i�����S�z:V����+�H�j�?`Ap�RPk�̬�ͦ\Y�k	��n�"���
����"-����,�)!�1�.��M#�0Zi\��^�~�f�߲���Ň��(����_+#O&�?h�k�2g`�l�5�54Q���Q\ſ���������ҧ2�2a�j�
�B@.j��N�_Lk$� ��$��B�.�!�|�>(�p�����T���č[r-~\�}�^����5ӽ�iFK)��Z(!|�kj���KSu�y>X�H��!ܨS���B�+�����Z�2-���p���e7-�*�дŒ������f���v9"�@�T
�H �b3��L�H*���-["�o�,���*��k�p��y�f�M���9o��_Q�ӕ�`���s9�����|��;I��2��p�7��1?�G�,�N��a�?�8(L%W�YO�N�x�s8��|���w��K&f
��C/T�p^X�K�n�W�����A���D�4s�t��n�/��][C�y��&]�z��/����xM�2�2���mA�B ��(�iߓ!�"�)1v��-���a} T}s\]�ٲ�^��R��^�Ua�o��Z(l2��M�z�2�ׄrC��-
��\b�ݕ���]s2��K�(�$�cK��Ɔ���2O0��Xhewb9Dl6��3�<��|�3Q��Z+�"6�w�TUu"��[�y�0��BIXr�!2�Ȏ�֗���T"��]����π�	I�u-�[�܊?(G�l�E\HE�ƌ�H�mx�<��]����t.%.Ne�}�e2@�gp?�
g��gHAZ��&+q{�)h��o��p[�	����^y|e��w���F�ˤP?-�|�Tm"�z[�/���>����w=&�R�q�ZD�r�ƭ��
�����\H���Qs2����)��=����[�>Zm��ՖG�1c���n{(�����Z�������z{E;Uj`��dǹ8A����9o�pu���}鷆Tۨ�갰pT��aU�-��ö�Jw��$�o�$��ppp?��a��4�Æ��9���/�K��B�dkۺ�M����{0̰q"��s�I@�OaQ>Rm:��n��B#�TΘo��||s���:/���sT�w!�T���x�?(֝��0�{�s��1%Z'X�R�gk_< )BJ����ҳ���a�Sp!,9�#���"�]�SԆ�%��|iu�������W�����Db�ŧ�}:k,��P9�.��H�xⷷ�:꜄�H Ӷ���/~tr@ج��#��ؖP�F�%�tʣ6�TǾ����Z�O��k�or)D���*cQSF�w!�D^�A֦�#&��%X�]󓿓��1"O�jn涛<��RΘ��w�!��}�r@w����7;�~$!�Ai�-k��d��S0��q8uu[)@d����K=<:m�Ua��"u�:moAף?<M/���G�Z���U��T�̋JG%F�;���A<��S�N�c�C��7`��T!I_hf��[x���g��D�f��
a����0[�n��Z .�XTY�Ѿ��<��ԶJ�ʾ5@ϡ�㘹/�����`z�+���U�c��t��^:[=|�Wi!�r@���As"�ݽO�&ɸ�P�a����׍�Ӆx�;����+
/'�8�wض���l����Tl+^�><�Zj��k�V�7QvJ�062����J`�(�<�(M@�Dʹ"�ׇ��i����0�C��Wԟ�y��0,�C ��2��}�SCz�)uM��ϘAJP�܍6G��++-�F%ڐ�Z�,(��o�{5�&w7�E�ǰ?�p�hS�?�e�c���Į���FO���2�+$#-�\E�A|�/����'�b���>���ӯ�~������G I�ԥ�� ٴ�1��3��� �E^�<s��e�C��/j;�L��t���+��ʝT~��Z����fȤ>F�]ϡ,;����ϖ����<��N��Q�~��-7��C�.����,���do���%��:��(Ý��������Z�r�$(��~v�C��N;��<>q��u���V"V�<Y��F�+�~�V�w��;O[�f�i�X�.moDB��JN=������[M�����U�TP^��T�����y���0<V<�4�������V�b2쎂�nr�ָ�pB���H�T�G�����x�Q�ϵ�i���!�Eo�a+�~�7jY�DY�_�a�O8�o�[i��.�Ψ��2�w�6F�~BN�CɜWT��'[�LXu*0��n�h�x�R)�7&��Վ�<�@�N#��УDq��#wYk�i�*�$�#�7P�
����aq
o>���%|���(�ʒD��g��W�M�	�������v��������~���8L>��K�2�^�'���Ĭ�(5)-
_(m�>���6YM��_�+Q <�H�V ����B�:��.�AlQ%Ĝ�θ��O�=�Zl��K9x3G1��E���GE�>߁�����ȯi�zG�L~��N\��x�hQ��
R�����yM�E�^��鹧�҄U��OE�Vr�b-�!���G��f���z͵~;	Q�C5�Ѷ.�_`|"|��?�D�銯�^	ΊD<h�l� h�T�o:L��!�E�V[�N�u�R�����y�\8Ub)=�����'�gf���G���
�/xR�I��7�t�';%Y����3k<��_\4U�����vR�6�G��)�^��5+Cn�,�|�8
�xC�+ɲ�[�~�.ٰڻ\kD�j�,��M�7���.JZx�����k�h+l�-����BW���3��(K6��zTqx�B@.ɗ������_z�ܜ}����r�t���R��e��"k��i_y��
��#���HH1L
9���ͮ�[;�su���2�y�J��5v'���k��>�Q��$�"K_/pGL�ꨁ)З}�u��r?��^�]l��?}�<�	[�.��D�;k(���(8%�C�`�B|%��ՈWx�eik���/�췾�f����s�}�cBɰ����{����H9/&aW���/J�J���q��i'���L��y?�������N�S)t��􎹇QϠ?W��Ҧv��߃�9��`.�z��OQ1�,-D��Ұ��HPo�/��]�r�iyb;���L�>i�p��Fd胖�y_��rx3Bg e��#�Mˠ����^��$�n��~g������a�w��y�7�ꆾ��&h�� ��Zsf�!��'��L�R���-׊k�1��]v���9��z��4��Vv�M�}�Ods![d�b��|�=_K����_�*�:cJ���98��\�=���ͅ�+�z�|�N��2g�ׅy_xtU&���?���a������e�La�K%�Ji k�	�G���/�%�+�i���C��oI7@P������H5M���|�����6Jgv*�ҫ�����a��V�$�� �cI�}Sަ36��9��F�[�r�̩�th s��˝�a���Yq�W����R޴�v����*2��[���/A!�y|�2H&��ɓH�_f`A��]k�o\Ư�+Œr.��"7C��������>y��/�����BU|����q-�R�,Q��:tN����&|O^�cݥ�ǒ%��4�b!��[q��� j��Zz#�v|�l��i��9�U�U�vE�P�d_�F��B�ˣWm�g+\-A�MBWs�H��I�a�&�� �*��	Vr���\gBFs�!�B�pX���=e��l>�̜��o���@���8.V�K}��+��.�&�eaՠVSܟ99�^`:�y�Ubid�e�h	��a��?wS��ïu.O��NC��C���;p��w��cE�tPmz�޵�p�Q��T��^�zMv"薳�j�*w����N��=q���B��?{�ךv�q4�~�W%�(�Jϒ/w$�e�4�=���t��:��f;)�?��3#��������>s��m���,)�#i��ɑC�9p�%�Y�ոH4��Ήv���wC�Y����};t(�xDq^��5N��h�v&v_����|LemҦ���m�p�C1�ͨ�;,��Y��u�οsN������Z/Z��F$Ï���Fit�������Kd�����w��{5&g�萘72ݸI���8�s �T��O�����Q�b��.�ph����X��ڟ�D��� �~���f­�O�ٹ����u���Z��Bj�4{�+7������i_x�%���TB�	�{�%�������z�fi�a��5�9�&��$�W���Ʊ��+k���Ni��ɺ/��K����S��چ1�oO���P<�`�����?���ǹ�!SG�_�6��C�u���6r�L�N�5ݻp�
g}����y�0x�^�Z�BD�ݟ�8�:�z�A��ޓ�v������W����WW"2=���0��齔�	"|�
��t�Q�&7���*TP,^�;Ed���_�F v�6��rB��-e��̩��am�1^������Ab�c*E�s�?�͕�Y�ҽ�z]7a1��t���d�q�6{dƒe��H$Fh�o�]�_4FaH��+ڬ�6E���3��2O -!I]X��[���R�I�=���uoT��� ���S	�]�˻�Fk��7}�`�`Ps���EH�n��������B���j���73r�8���
w?�䡧�s~�[�,��H�x�(|,���
>5��xU��W����I�??���>�!,�O/��ݗjc��BK=!{���7ơ�I���t�X;%�����wa��D?chi����T�YL0=Nn�wx11ɤ�GKZ����P���q'^�?&T�����0��@�1�x+ˁ���U[h�M�V�c[>�2���\�[���p�r����k��U�*�L�%��>����xq�� k҈"X�y�M�}�/�{��yG�Ĳ�s��fe�̷03�*V�H�yYl�Q�/<6NΞ���^W]��� ���r!8�Uѕ�"F�~�2�'���U�i�L�۫�9fRaoT[,\t!�q�D��F�.�3�*���ft�Õ�AYW�N���A�*ّ�{Y����rO�-�-�w	0�{AM����'��@f�҈-KbA�$�cn��P[`�ɇo:�	������U��b��#��������q��+B,)o���f�;�.2OHɯ��{���8㳥�����=��_C�`K�^�/��;�^�������h����ӊʿF�>��^7�>��y�'ߟ=�BL|?,�m���5䇣����a_J���X����?M���&�w~ �>�&r��rҺ@���M�j���l��Ky����L�Y��O	��'t
����,Kb��|��=�y�^�Wn�*u<�7-��+��I��^�/W�)��¤:�o�u<�?<�5�����v�?'���E�8�ק��{��l�>��U@�5~�t������f�(�WPi3����Bd�9,$P�`��G�*�Qy��X�Z�*$ٍ���;�\�W�H�N6~w���	�.��)��SÇ 2�l�C&R���3I(J�>���|�s6EҨ��(cfv3��k���?���Lm4��΂	`E�+Y�#k��[D�� ��ٺ.u�1��S��c=�-��م�:>iL��X�a�E�~`�[��݂��z ;�1z��M�5&*A���2��̣O��*At����K�a�4�z�3F��ۭ���L���+k#XeIJ֑����,���LduJ���ҭ�R.�Q� ?�/I�;)�ŏ��i��Jdeö�I4��n��>�<��,�������$e��k-u*A����D���wjI1�Ļ�����(��-��DC�&L��hTP+�0�%��q`>�on��C�R�E��SVE;]���������ǒ�,"�rk����ggV��
�� �B�t���
��Uk4��w��Pm�ۼ�l{w,I��HDF�f�]����0`�0���v�zZ�,V�X�M�L ^�EWG]��hU��g%�9��K#c�9�	���a������f�@�����+A�a��ܤ��ߨ�":���N��e�b�Q��w�,���q�vd=�b����啈�S0��UȐ�/��q�u��KGe�s��r��������e8.�q��PX�3�����g�����%��N�Pe�@��g�BukQ��<�p�Ѓɪ�u�������ml�����[��m�)~����(����h���?\�́�G������B�h6�c�5�y^fm�;��Vn�u���ɸvϒ]�뜇o���rX��n�o��|T���l��5ƕN�Ŭ�ר���~��ʎ�i�-r�)ҕ�7����_��B�����@�5U�n(X�#^��$�03��	�A~�]_o0|��el���֨B��
�����\��B�cb#�v�H9�R��z�4�VϹ���s������l����E��D���:Ը��z���zp��5��/���f8���Z��
+�Mоl>�p�AbgZ�B��m�+�����r��u�@}�� �_9~�Wּ{�Wg>3E�^��Nŉ���u�PŻ,*KJ̖��2gُ�ơ|_�7���<Q����h|N�y��!��l��fDBz}��/�R��~ѧ`��sթ�%�Ii�>4�j�i%q��uf�xg+�[Cݼ
��&z>�4L�ʪ����e��EXB���&�5��m��w&����" ]�Eu���f�����9�w��
�q�Soq�KD}���F���޶���a��6��q�6�E� �v������Љ�1L�Lj�{^��6������O�ku�vs��P���u"G���.On��*���ߪ�"A���d�eai>��'�\SW�ǿ�L4G���y?q�r	�� hI����|
�^mvO�W��*�
H�EJ���%K��@��H�����Bǫ�s�b'�z�f&l����Ɓ#�H��Ō��V��ԇ�U�)W���~a"�ݳ�N�J��k���6U��ɮx_gˁ�Y��ILưw�@Ī�`s�LbJ��h�M�U�5�+\&lR�/
�	��BrOv&ި/��!L�PW�ΖK�2`7o�(�+	���׸V�c�g��g�!�x�h1) �2ɥ8O���(��M�9�O�9��ޒ �a`�R�{�{�T��A)�X��g�.Xu�L:��a���W1�wy�t�x�O��"�?����m����VT1�ʛ�&������5T�TjN������V��DJ]�uF7�pe%M^B{w�*�~�.�M*W�� ���2Z�UGl��������<��$5�dio�'c!,���Uj��-OƑ!EW�hFK� �k��|r"���F��+
��,����[��x�%t�#^�GPTTi�����-�l������Ff�=��v����ީ�b!�A�CM��m=�3�̾�Z5Fθ�1g�ܣ��n'��-U�`��ZN��Ӊ����#ȴ��D�S�L���2Y�4}3���UX�iZ
I4E��6�ʛ�F2Vل�SN�'��Lk�:��@����C����u�C �����Z6Vl/(e��)N��oUh�WS�+�����$�+e���?l�}��u��|I��k�TNA�\FZ��W��_�H�w����qqE0R���Vb�U�8<h�:&��DLo5��Z����R}k�kܿ��#oe�l�W�
����	�\J3+�Qd�PA;��as�ƭ��s��PP����d���q-��I5������7�Cލ�����!2ߔ$��i���,a�e�:N	��>�ģY/�D�_%�kil�t���¤&���!�׭��'/��8���i�u�,���=�v}z�K�U�����He��YL �S�g@L���R�����9����Ðj���vh���;όƦ��-�U�>Ӎ�L��uMA�&���X@A<4q� �k�?[v��H�%߷��"�^|��H�����!�gI�q�4qĪ5R��B���
���b�c錶[��]��D�՘Y�4��mJ����!Nn���j��S��?T�%G������+o�ћ��qT<_o$�gQ=*W8m�}k��0c��N;��� ���FN��O�a6���\�&:�	9e���!\��Cs�|j���![�$��<�(Y�2O̾B,@
����߿�)=��74�T�7�0)S�c���!Fn`�N���)�ٔ���8E��稉�2�R��5B¥.0�D��E��,&��O�E�:L����W5��2%��j*b%ؼ����jDD�~�8۞!ZRH<;逭�%�
��q��ƨBK+�X����R�]"3rG_t�m��L.�x�Sm����$ͫ�0ю�g �& �x̵���������ٹl�<�Ǳ�4����+�>Ӱeio�;�$���[y�a�;e0�����@�J�s��Й`"�{P,2g%8!�W)��O4��k�&����k���J����t�_��X�0�%d�P���aRc�B�9�Z�GGC��I����:����������H�%�2BJ2���jcɫ����K�����O�M�����$���!�D�Fk�F��Q	Nx_���en)�*�쎗��8݄&0 �edJ�'��v��U���K@�.|г�>�/,�!1�R�XIb�iF��ʅ!2�6�^�|�l��n���Z�]��[�K���0z��ko{�gGȫߕî��6�N۸SZ���:\Z۱��`Z����r�Օ<�t5���J�vo��̑�;�鸴���F诽���z��'Y�~�xx���%d��}����淣{2�\�K$�V���j;�5|V�k�_D�06�0��~��w���K�
2v��.8�L{I��%�)��w募{K0(��b�&���1������^�d��m+�U�؂)�섚�#Ku}}��#��UKN��h@J�ï���P0H���V@�_�̧�ʗت�.�p�)E�����8��̯�Ǔ~c�E�~�Z����"�~���#-�4e��|��@r[L	��OC.����ngr�{����Fw4���qg�c�s6�)Dbl ����TV�-���%���9�Q)�m
>�H���h��Zv!{ pA�p=G a��*�H�(��%�t-7�Q�ȫ:��jc�l
��Ue*�<�B����B�2<�E�����*�19�T5X�%�Y����'�r�T��*,��Oϥ�sP��Nd|����!�PA�1��_������v}C�d_��Т�BQB����\��{�Q����8�ܜFǏ$+�,�BCH�],��r��¨���b5D�wpp6K	�]���D�ʞ�D�9�q�$�-��CsG��;k�r�T��.���I�_&}ǩ֍pPy}L�MD8ioӲ���
�4���ꈪ����ˡ��DJ��s�пF��GG(Ζ{���W!p���-�VG�Ӎ��}��{Ц�cB�or^�|d_��������/�ˮ?�C���x�ڌ�h@�rαPʸѴ��q�T����m6l1#!}&�i�~�^�Q�M��rB���h�����%�mȜ�y|Ś��������E�c���� ��җ�0��+���� !{3�c*!��:qe�4���O;۹�����2��W�M�^	�`/�2�Wx�a����{�"aJ�Z �%����;�DB�����`s�ן~l��n�7�2�wkL�����?�x~�G�<��[M�տ���m���o3��d_�]�T�Ch��tsٲ�����4X����V_��U�	�~*����k��>{��Ƈ*��Ȕ�PRux%ɫ4��;3�ކ$�S�}+i��}��]���^�bw���'��P8�5j��$RP�M���Ď�%�߲ �&0��#��9c�b��E��#Ҕt����?�{ޘq6#ƜZ)���	2J���n�Zr�|�^�'�?敠�E���N:7[��Y���K�V���(��g�YC���q�c�g�ύΦ�[N��g���>O���3,�_`ߟ��O�$�k�ͤ�2���8�$ߢ��?ڤ��� }���mf����p,�!�l�M�����wBOH
8��\��}!�'^x���$i������x�n�=fM�8L����t��ʃD��n>j!̇n�A�H���.��K�tn�"�

�m��?C&�)�]I��'G�n�<wP�}�Bg>b�/Z�wF�D�w����V��ꨪ~�R��JƫA��_��]�"O�K8y"1`����l
��#��%�L5NS�g�6�vA���e���xSC�%ԑ9(ڢ�h}�?��?�KjT�9g�p Z��u�nh�r>�fy�L���}H[5�3%�]/�����ْ�4�5��*Ɣ �2Q�L��}�\c>�ԡ�\��3�LdJ[v/�{�C�d�Y��f���T��V�`<U��/5�"�Y[���W����qu}0$���6J�k#%>��-?S�xL�֙T�b�}�8�8��qgW���ׯ��3z;m���T^�׸��3Ͼ%7fK�E�5�#s"X�b����+�GK y�R(`�p��h��Q{m��u�-�f�R'�fK�� �<���*Nk�+X?�p�e7����+~Y>3!>1���-��l0a��8|z�Ydk�	��~�S�6���
p�O���/;\NRs�[���N���{1��\8j4����,��B�Ci5��o��;�IP�е�?_ϼ��w��J�p}�O!J�btC��UB�3�~�;2d�~�a̆v��=e�}���~1�e��
� ����h���<B�(�<�1�|�!ei%I�;PvjA�!�Z���ƨ�R�2����I� ��Og�y�`|��DV���-�L0yy�|�ڛw
ɾ �n�O��D��B�E�8��j� ������	�9a�$�\����P�ow`����C��~K0xТ�Y�4�zn���z�C`��?��(���j��nO�5����
O~�ʂRn%�$+(	*�E��Rr�&�^�ו�fH�qr�������]���cQ��+�ֆ:_��[)1��p�%v���Sl��@Q�����Od E{�;v�W2&?�y��O�wA~8U����<���u*��]�F�(��_�4�Ƈ�2�	��Wq1.��-Ȏa���>�<y-
� �i2Ae'��c�@Ͼ8;T묈�V_"����j5b�s������n8��]m���Ƥ8�6YQ\��F`=
��윟�8�f��
��ϖ.��)��Y(^@����p��*EH�4�b-��pEw��Ֆ��f��$$����HD�H�繥PP�^�З�s�@_1R�'���	]���r$�y���Ge-�1�FOtKm*��ΛW���-�� ����'��P2�,8�J*`��9;�=(��B��l�:ɦ:	�!���]�-N- ,o�Wa�@�ŉ���d_F�#���{f�摞����T�@����M�� �~x�}f�-q�/��F�%�UD�A<:�������J9�T�m�H���
CiΪ����\�����V�h�g���p%�:��ψ�����Y���¯�V�5�Zk F����ԉ\k��}��SF�w�H����7u=k(�����Q���H�Kh���]��9���R-���Z�g��.Mָf���e ��G|ӥ�m�.�Z�+r����L	
�}����M7s�]��ф�qQ��WT;��m�����yEvј&z�~)M6;`8�Gx�q4׸��؇�����	]������]�r��39S��J�N0C�NK�z�v)
�Ɩ/�O"U~Aٔ �s�:��E�G����b�)2_X���`��9��<&;�yPU"�����_s���S?��N�?�}tw�ԝ�M�&,�`��m�c*;��O"�d��R����I�5B:��4~���V��ؙ�����	�Ej]b���f�3U�Lt�Ȱ����߄�q�,q\�|���6�P� �hR�F�"�n���L�F'P���F�x���d�x8�G���(�BY��r�F��"�/wcz�<�7Tҕ�GA�⟹νW���#�:�rHRHI꽄C/S��ԇ��wD�}3+��A��qJ��eh{��M/h-ae%��y��^&���y
w�I$��L�U�הﯶa\c�DWFɊ��-2{8�2�vGV��6FӒv�K?]�DBl���Q�_�B�ըb��j��	�x�-J-%|B
�Vށ؁�y")��H�`]�'H���V1���I��E��huiɢ𕶳��I�2<�IK>�9w��R�>�U��vIȆ ���Ȫ�E��k�Az��H��"EI.� �f�f'Xɳ{����\��
�C�
�m2���L*D�}̘�e&�p��ߵ3T�EJ����)�L�Au�U�4G��P�r&_u�k@��W7��
��c(����d�L|���4���#�r���N�I}�-C�0U�ldA�]��}`�~BɄš��E��Oѽ�Q��y@;Q}�䚒;>�4p�;N~��M7��;�eq-v&���[~OZ�]e:�!���􈥵ա菀�.�0��Z�NJ��2&#�PS�$�sS�/����d�Hγl��Ysb$���y�G����U;x"ǟ��TЋ���8˖���z{,Jޯ"=�5zYoc=V���K�ʖ�c�������/��0-�7��Oǳ~�����EXe�$��ZOV:�]�����c��i��{;tk�H���m����&�+��gC>]w�4ٍ�P�Z�
�h��[8�c�����l�:�bа�6��ZzR��X�2��*~U�n$Sb�����rF��Az��E?�0����1d�͌?�G���^ �Q!����Pv,bj����:_� �W�͕�M�� D���$b����ї�f�8�!����T�>z�W���k�_�Ë�4^�è�T�}��Q;�!���<���u�)��=	�L��h+��� #@ܿ�����"���`Oud����"<j��8�e�hoieC�H��'��(�A=����/n�@��Ts�j\#��(P4X�pZ�qn�7���$��G�t���MTF@N�7�`U}�o��H)r�\�V���`�q������'D5��ͭ��%��o�V�@�ݸ����w*�H@��q��̈ 5D9�`��
��fK�;/>�ߋ��v��!�ё���hG{k�Ũ��=�dY��S"�њ�CX��T�������Ei/l~�����֤!��Z�e�hjlAo�L/]�{�n�9��Ir�:
��s��Cs[;^:�{�6��<��� >t?XuNNEb�鍌9	��pI$(���===�?!oC��;9.�ER�W��E�6�ߨYL*��ᾣ8r�
�"�,Y��"tn�����Ʀ����a.�۳�#�������840_K@Od�/D@jp��r�ip��)��%�P�(u9��_���!.�:��#������ڨ���{2����A�)������wQCZ��BR�4i�e�TH�J�BiN��&�JQ�j�iFm�����""l����}VI�06�=3���sx��qpxN��s�4�Q(��b�J$��7�R�o�����)�:ĤpZ¦�,(����m�z�Y���{7�v�k����@qah丂J!���#�a�>4oh~{�w.Z��+O9e���d�'_���O~�bf�/�Z��$ǡ��2_zeh^�XgC���X����x��o՘�x�C�6<��?��5y�eKy���k�Xcϑ)V���F�j�#O+z�X}$t��Й�"}Mh��b,֦|���E�:@y��*Ι���A�҇�p��2HX)n�⑑�ST[��E2��W�.ִly�Y�v�@�E�߾�{�1�L,_<����1L�,px��}}Eܷ�9���##тj�`�TB���
hmk�'-춎��1sO;�ݷU#��L�܋��w���X۠g�(+��	�����$RIzb����6��i����A��~ z�j�A�*�G����Lu��5#�ej{Է��!為h��O�
$cG���y|��ƹ��9n:���8i?��#mOe[��X��_&��&{�'���[Y|��X���qǆ./��e#~�U�L�Ο��T�T�j�r�jlzl����Qƒ%��I�~��1��Yjj(�H� �J��]xU�
V._�MR�I(G� 0%a�tQ[Sc����	��]��+���Ӽ����x����	e#"JX�tf͙�߿��K�ԅ��Fz�G�4���9j���e0&P%p&������ʿ�H�#4~�p�.� 3f���nܸ������6�9`E99�ǠN�fϞ*Sz���ػw?����N�L��Ck*3Y�F/^�\.��{�ؓO`��[�k��l@��yVGF
�S9�*�A�&�n��֤����9�A��'��D]�Na���2�7�ho�1HE�&;�R.����_��zD�ڿR4mp�"e5!Rv��?r��)eB���������	�5֞B;�〮��ͭ ,�1t�7H"���#���F��G�y�s�65qʐ�*#�27�JJ���`L�(ĕ 4�̂�҆ʀ�����}�E��sO^V�f��gw?����_��H�]%�s	v�J|�İzȩ�Ђ���/[��e3g�!O���G^���'�����]S�t�(��2�.8���K�-��s�ek.���3f�C�ǿ�g�C7b���'��5�$T�[�G���ᧀљ� �t�R--=;�vE�K�9��Ƶ��(�&̐�=�QH��7&nP$@�7(r���By fy���W�?bd;gV`��T�.t#��ᥗ���g&��F�L�ރ��V(*E�U�9�����<k.\���C�1��B�`��!<���xu��B��l��##jBK�����6w�k�,9�<�|�è�)�Q36t�G��~0������hU�N#�I!�6 B����б2�r�vM�m(U}��BՈZXRbʝ�O=#�t�Gs\�����u��@�Z(xŭ�a1w���	�uڇ���/���\��&���=�x�'�\�W��N�o�L����d�;��ֿ�<�8quȺaI�r*��W�Lc\���&G��ꝝ\��%��s���E��SıC{���{�74d��э͛7��u��<�-�i�dr��H�l���^��s}Æصs'S�<�Hi,|�ZH�[��,>�w�Z��M��~	d����7&"Z��+��ܹs9:��j;w�`j�0M��)�������oꚮ㡇¡�Q*��;��CR4�ѓ��3��N=u!��w��l~�>:rS�uj�I����~��r
7����b;��4p���J�̐ք���	��x��ʶ]�9T��p�$�n�FE�p�i5LV�Ǭ��2|��%�4ş'�5�ߎ�ZDu��Ԛ\"�ǘE�� ��ȕ;����Or��v���-�6PM7� ���8ym$�e{˔<�S�`Z��^Փ�G�őAM�&���U+Q����WCp
p���E�Bs������X������E����ݬ��f]d#��B~��dC�*.��PO�0���ՐU�Ց�����>t�]o���DI�{��]�����J�>_M4C���(U`����T�N�n����gްlf��O�2���n�����`���WEF�T�dƴЁ�
�ͿޚM<��3�r����=z�샛7wo~n��g^���TcǅU%5�h��I�I*��ЙN�k.��s��\ u�^�M�R���0�M�'�q@��i�;"Q�-�;|O�4	QD��X=.�DCH�2�P��Qs�>46d���SO?���!�j@�⠩�	����d�8��� ��65�36�Lu|�'�n�QM�90�}��p�Oa��AJNH}��T'ݒ�6��v*�!���Ђi�`���ֻףzp�������%0��Ǝ�JI2��h�d:%.k�:NG3�A����F��r�{r�"~�@�f��L�����T�\8	C�ι��H�S�����K<�9�>�.����D�~�H)���o��>���Ll0���le�A�>��;�輞o�6�����O��zLH���t9�ki��s�=�|B/j��#�*0I�[�#�o_s���0�������ɏ_�ŧ-��}�{��m�܊l*�S��Ē�hz��5�\����~��,�c���oKjq;�ı�xA�Ӗ.�(���Gƍ7ވl:�F�Ɩj�i�P7��?�O0�=28�{�۷o��<.E�t�l�5��O�S\�V�T��oȇOɧڒ�MX8x`3����s�=�������x�)ޞ�BjΔ`��?4�w��J��W��Y���^Ǐ�f�mC6qʤ�|n�r�袋���hj����]���}���W��5s�jCU��IP��惜���1(����l�9P�'�Mf#G����`�娫�f�H$<Q�.����ǁ:���FmR̔�?����e�5�v{w�g�~Nz�=!���`@��XGqt@G��SA�( ��K�J	!B!��v�����yߓ�s}����I9g�w?�]ֺֽ���b�A#��C��ƀщ���6P~F�nS�l�#aW�j�1\RcQe�W��g���rUP�"L�Lբ4+�^I�$V��Ŷ����T�j^ �@@}V�VU&�-]���{![���/��>]��<�*�<��\��m~�o\�M��u����q�`���[뾴c��OM��p+R�*�N���Z53�*<�\d\{��K�ϸ�s%��7l�f�ֻJv��D����D�*����Ys>S)��V�f�Y�w����p�)��=��>OGw�Ю���b�<�j��,�V_��R��LMU���ć�� �!��	"��UJ�5)������:�>g%�R�(�`��.Mf
��ߋk�ɂR�.78	EV
0�"pU����^İ�z�C~$z;�r�?\׈-�nA,�5 ����VS^����YC6�����#{JU���@o��ǟ_�O�u��
�W�(�(te@�a3��fG�ȑ6a�����zx�m(q�ͥ2�-�ēȤ��Ȳmli��_�|.�ة�8�v�j����<��4IT���@g�.�C�3݄�M%n�<�$>�j�U�Q*��ֆf\6e "0Ϗ͝�%&���ӷ�L���I�3�]�O_� r�?�w���4Զ>�F��`EA��J�L �9+aY�q:�~�����Rlp�yN���Y��0��XRՉN&c�"�@���s�c/� ����%ȑ�ΥV��T��f��R�7����݀}�~�j)#	��b��EȦ�x���g�>1����R'��c�].Y��o��$�w��(�UXHz��
�_#��h,%�������#��[����ϯ���&��Sn�{Ȥ�{���X`Qv��*�B�7��떳"L{�M6�y���зlۊ[o�U��.8����(۳k���=���}7��ήn�����v�鲰�g�B ���g��_\~)b�^X���w����O7sΟ��C�x�&w�ꫯ�wo�A�h�yi��~�\Q��hrbؘ)8�ы����C	V��*D@G�:u����IH佥����(1y� ����UW�ӹ����@&����W�1.���sˤZ)���"Lm<�iP%/��ht缋r�e����(�[��iE�My�눒�����wB���I���	�J�b.!�ՠ�u�����Ջx���A���Ī�u�) �#�������j�l�xR�'*�MM�kl@4�P���A�3v�7�ȡ��D�\@�L��8��)�bЌZ�$+�]�*̅$|�¦�̾��sgm������a��!O���?wF2��y�L-N��j�Fhu�`3U�[�o��ٳ��������ؽ����	�^VI�%�ZM9n++	C�R.ej�B�V)'-�J�f�^��K�8v��osy�e�f�̜[ɬ�Me��O�
j�S�J�: #�I��egV=�ɮ�V�ޮC�<���e��n���J����i� �F�P_X���� �?x-5��:�X�	�{�<,�?{v~�\��x!�-S�"ErX��WC0`�C+a��x<f��8�L����V�7r�
�8��]�y�}Df4��EIXд�U�	�6;lf2�lZ�4�;g)���o`v�e~^*�c���%����E��Z��&a.P#�����C���O�dε�j;���m^����ga6���p��E����y�8}5:ڙ-���ҥ���7)oh��	���w���w#��멺L���BW��5���R����nd�W^7F��1���y�ube7�u�D-��g�pGy�3D(q�ɟ:��b�b�S0�*X-����9繭�[�[	��AƢ�r.k��f�?��-x��pp�'4�B!�ŢE�ce`{�����#���d\^/ �r��x�_|���N޲�=���*��8��.;������R!�1c������&?r\V wuu���A%fX�2fa��_����-[���n{W~� ̪
".����믗��P��?.?����fA�\�n���f���۴�����5�::����P�}|$��2&�"�O�?�8l\���ඟ�!K\�9��$a�]%"�bA^׿��X�x
���.ٶ�pP�Y�(j��_@Go��eT�pd%�r���T!��(8�%G^t�SšZLdl)7,W�Z�DY&WnV��˦��8�<&�<��, t���̳���n%��0�
���Ha�s�eX���׫�i�'[\v��Ț��JaB���7>۪��bL��2���X��E��ل����.ŀ�,��v�4Y`)��Kb�);Xd��fOO��w��x�~��^7�����X���L(*b��b*�M�b'q����ŮJ�b�!���ۥ��U5�J��kh�����_���F��o��������ښ��ع�6�;4�fv�3�<�~���2C�f��T�_3�o����|����Ǿ���?V���|�.	]g\	� �>r�Y�H��,ʥ�$5�X���|�<d���ӡQ ��?TZfHx��� �r	~��<H��g�)c��*eU�.�e�ftS���UT�pH0�Pz�9�BL�2�<49&t3�ݧ��t�>�F]Ѝ��F���]�������`�J�D&��x4h�"*�B!<N3�.ZZ�{��)6�5��Ďw�![0�Tg����$�
J$�Y���jlmhliF�b�ɮ^�����;X��]0	NND����֢�ܨ����J���Q���s���a��L\�T�_���_��g	���F�9����lIvq�$�\��m�]�G���C��Gf���f��ϑ)�C��*��u���"���5� �稾�}�����M�G��\dm�°�BQߵ~�\�`�*��tM�oͤkS3A&�t)Y���1H�sc!���)�|�P�HХm��}ɐ������I�?nl�hL�"̕~tӍX��oس{'�[����$qs{����j�� i6	k��=
K��,��h� 7l؀��m(��fU�YaA����6�����|�3����.���@Y���s���j|�k_����e?�я�l��&&p&�;��~��2ƺ��{�w�����StЄ�E�W�e�.��~�3����܅�n�I�r��'y�����e�]x��7�)�ا{v��w�'O�B6S�R*�.�NJD�z䑇��y���W�q6n��ۏX:�	Sg�/]�?��0z"I��22cq�W�uʎ���?�-����;��Y>#oS�����Yq#�F��������܈��ȕ�����5тBQ�\;��pHB7�]&t,��#3�J���}�a�A:o�5���T
��_8����
t?��M?c���#3�3�5e�����Q@"k�a!Z�\D9m��l*�T,�\&�7��_�B�tJL�8Za1�0�5��bD<�����9�s0Y�:PFcj��"	*c,΄m���l&Ѣ#/⽟�jox���s^8��������h���+o�۲�ӛ��.p�B��)�3�Iv�%��b �췙z�6~鼉~.R���?��[��[v��N�Z>W�"GT3j-?�Mt�)Kg��ĊV�Yd��)��Q�Yf �n�
�Շp��č�Ř	YM��T��{ơ�"�aJ0V���dg�J�U<u�.�2��w�!�3$��X��Gy��d�D�L�tJ��nE&��fF��G�@H�,�Xq��{,Ҽ�q��r��U�\�1e�,�JKB.�.����&�\���p�T������C*XJ�ʵ��dY)�IJ�xnTs8��q��.�k�m�6�2\:|e�{�x����M���f�#jX.��IL�f���L<�
=��K�����Kȃ`�RGZ��ݦ���yJ�x�dn�u᠘xpcW����$cј��^բ���/.Vgdi?K4:vvO� 'T�3�a�2�DV��	�)����D.�߾+I�tszqȳ*��jU \�<�݆�r�B$ɰ�Uݠ�-�j�ىH��3(-4K�O2�b1���Z�ږݕU_2��O�XE����� E�P�����-E}((c���9��B�\F�\&��7�:&N��)��o&j���U'Lș�1��$A9v	���]jI����I����S��TƉ#��L�?7K�Ё��띝�%���QI����H�|�˘>e�<�+VH���$EcI���qhVY\t�2\��q�*��R!BwEnD�M�ϛn���G������x{�fٳ���d"�ӡ�=+䲂^��]�ɓ'q���[�iHfX|�2�;w��7��CR\��b����Ĉˇ8�ҡu�{ԹP����ι:��3�eR�G�Z[���xEr�Ac�y�	K!ANzɗ赡��N� vf/������{WE,�`��a�e�L9���y����7#�ϻ�s��0[��	���̐�d��    IDAT�x��� ��
�~��~�%����%a⹦
��ɢ�J!��+p��aÄ��'d\C����	&��:Y�"z)���D�|�"��XS���/�7�f�@�2��QJG��X���pp�̩S^?{���1��	�II�H�;��Б�ol�<gߑ��k&�<���.���hA]}X�'�&G)��L��Q�u��x���>WB|ö	���zE��M��B�� wY��Z��fق%ZJ��1d� @0a�uCJ7�|E
��(�>h9�e�}�g:�3qY��_�d�)�τnF�T�K�)-$7Nћ�Ŧ>S�$��$5�M�%8� w8�y�8rɘt�C>$S144���X�c'�!�IʥK�2�q�J�����*�;t������U9����0j(��Y-�a��E"&��V&"}���!U��r5XnT�6�=�%3�o��%�ŦCC4���7X��v�O�;5���"�Ǣ�AG-E�ʶ2xcV̟�����`s��Fp��!4}hE2���l3��f�t.+sA��9CeWa��F H�D��	��:iX�nq:�g�V�8[	gbO�ad������&�?�uTB��g~�U��s�unB�3�����X�?#V�vMf��t	�T���r:B�Bd1��|�j������[*á9�ֺ�r�{T*�ē�3�°�Kd��ul�$ౄ6:c�_j�����ט�Y3��g��-f$q��u��?�91g�R��25�:�����e.��玝���|N^�����fΜ�P�N�-4i���a�r֬�kNA�),Z�]p>NMwkּ�����+�&W��I�˯�Z6����?��G��Ȇ�,=9��MoE�0w�Y�1q��Ilٹv_ �@@lomN�<�w�ۢ�+�U�%�b���J��-z�� �y��,g&z2S!�L�7��:K�|}}���3�P�A��K9��͢��Ӣ�gm�4y��נ g�/ce+��3\��N�Ю�f�r��97SIc����X�D��P��jD�:����ſ��B-�NL���Z��<�)�?Sr�(fԽ�ze��5UP���qi�B�\�L�]��=��0��d,�l� �ǃ@C�8br	����e�d�U>�Fq��6eG����\
~�͌B2V�Lծt,��kw���nm�q����h����wj"�U�k�f[[�ls�����$�B3'.A�.5�0����ϲ��\:��~��I�׿���杓(���BY1$t�$���K��ʩ�3	���dT��|Ht���/��3^�ҙ譗���>Y�E��I9���̐��lvs�$�
�6<��)�%e<!d~��yP)��t_W��H�b��:і�fD�}ȕr���2�#���.�����U�,�T�ve	$&�SU�������B��219�ֶj���)��
��;�3i��NI�@b�i�!���/�X�瑔ڰK����H|��N�3��G��FY7��� MB�~�)A�g$���Y,�q�)~�^��;��4	�'�E���e�bPK��v0��Gck��}����A4}v'Y�J��?v�dE_w)�� D�T���;%{�;��>�-k,��b��u~�u����_ê`A"0���a��ՙ�s�4��I	P"��D��l�o���j8����G�8ggd�.J�&�E��Й�y�U��\Mf�u�4�TḤ��_�Kuk(S�[)A��D��\6A�d�M.'��gK$=V�M�r�[NΓ$Ji�B�+���A)�����q���	��*�fH�&�!ÆJ���?�^�b�֦>Y�&�����=�w��޽[�/��Y��rv�W�������������w7�	���y���|��a�����
X��߰e���S kei�d'q�Ϸ�[n��\��_?��lx��v�v�K�/�uܣ�n�h��Ĺ��4J!݄1Ѥ���2$&|�����;��u�2�9�T�9j��Λ-�(�����=>�B~T�V�(i�Vp�^E��i_%��P�kr2��z'Ji�~��pb�"Y�g�ZA�p��,Ks�B��+!�v6q*�(�6=]HB��eY
U��z�%w�\�b�Q�[�7��L�ׯH�e+[I�[%h�*��<(���U"�w����f8\N�:qZ΢��9!��9�>+�Qb�3�|!D����sv>��,�����$耝�B��J�R�f�\�R��,����VO�w�V�j� jf�7��ɳRrV2u;r�L9��V������7�?�a�W���`U�΢}ᙄ���L�4=� Cw.����nїAJej@��y���I.���Vۤo�Rd�~R����c�7�y�%�' #��j�S+�U��iG��V��Z�\�u����Rଌ�Ó8q���\� aq��@P��wv9p���B.�G>}�1=Pӻ�(.k���E'�j���rM$LESl�x@�Yv�&�57\�R6��Y9*KT�y=v��)(CM�'DGw�\NXPj}�"f�[��sxܢk�K[����W	WUK4ڈ!˽�t��%M���v�t�<�DX��9e(e��4��������h�����iX��:X�-�JY�n����H�g6�c!E��Й�H`Qi�݃	�*�]�W�,.�lXPI؎�Am��
	)��=�3�9��0sp�&p3��|eZ�֐�E���>!\q�#�
 Pr}��<����&����xP$��ͣV�&	0\���ɕ@��A�M��%i���'G*n��e�8� ��^�E� u���U��x蕏 ��R���K�2pZN��B6'�_D��j�+y���e�A_n���%�p{\�=�й>U�4at������A�7)�m�y��L�A�򃧩�fs�I�f�pqK�*c�aÆbܸq���p;��ߣF�<�B�9y��s������on��W�`Ǯ]rƅ��,�kTL��+���ӧ��[��+�蓃�ٹ<j��$�]
��Y��ֿ������������.��$B>{�j̒:'^:z��T��ds!���Y$����!Ţ&���T��X @�~��Ȧ%�a1Ɵg� TB�S�$f����k���~U܉�S�(����0gB=��;hr���C,�����ϒ[ 	7�����߫VaR�ĭ�)��)>�U _���ml�:v{�hnn��Bn	@�T��6���66Ib;�3�ŕR��
���4G)�*j"e$S^T)�S`%T�#�JY�$��2��D�v��ETLuj���"�l���&�\	�s%����7~P�w|��c�?�����ЧL�G�N?�ȗ�|�U��*x�$��{�J������8ah�uM�?�6X�,��^�_���.[��7����L4|� \v�E��8��Ja'�Rʡ\ʠ�),��z.�����r�K�<2)���A�����������Sx�����a�	�٪�,yI���kr�2c'��$�F��pp�R@��u^]w� ��ԬҌ�CA_.��	ϓXR�f(�
�#���E��Q��uQ8�a�@�29#�$��m�}���h�aE[}A��ZYUȜ��E�gȺ?x����-3����=h0<N���L�$����f2����m!�5����
0��k��Y.�n,�KZ��
B!8O(r����"n�@�z��Ku�g<���kLq��ᕠ)rȚ@�żZ�nS�i*�Z����	;?S��20�ǒȈ$�2���P���N�lH�r>Xx���g/�������<R�_���g�˔[��[��Ƣ��B![�s�y4���S��Ύ���~>�EM��t��ZD!i,��H�T�o�U�`H�b7&�F�[lfaƓHĢ�����fe��7�	t^����\&-�Q �;)|4Ս˯�l�"ɗE� d��:�	�v�ۣ6R���HIm��f�f�IƢ��"�L���AF
v֚u��Y�:�=x }���rޫU�	�$_�U��ѣe��r9���a����)w�w�c)���
��e<�k�U����)��qH�pM:]AE<n�OL�F�9`��طi(ռ��|B�s�\��ht��@$ǐ�av�9��y�n��[Aĉ%㜑����ExV|N}�CH�6��l4$.�8D.�9wb�ϸz��O����V����VM��.>9ƨ¸�|J�ο��E�8U6�%1>�7;�#�X�[ ���N�u;z�,��ݲ�(U,C�ln�3'c�$Jz0�._� �9�KY���X���K"�D�J��'UF6�Q�X��0�.�����Τx]�n�HBh������.�7��5C`��9�o�����Ȅ��r	F�Yd0=S,�C�OH�Y��E|s<��/�3I��BI�/V�R��ŉ�=�����%ܳ�ѓ;SV���S�b�A��A��.Y�L�矍9���?��tg�5�H/���Xr�8}N�R��Ί�x*G1K	VǏ�@<���^�
L�1;����y����_C_<���nؘ�X��,B�ʑ|�9_Ռ�?�L4.2�	t�*2���8�"|G�/��a"�tLLX�ȳ���
[ɢ�X*��9;Y&}aiqH�H&(dR雄EM��B|��т	�x?��z4��9~�BA��XR=/U]}9���BfW$�]p��56���Y�I*ET��â�w��xm�6<�j�>�t$�SE�i	��L������N`\s�B�����]>��|��8U��Q:mr8���0�T�dīذe>oz��T��"+�\����>f�	ٙE#Dm�v.�P��64���1�q��_�"�h��L��A���l8t��z�i>r��0.��rL�6MX��`ԇC����t`�:����x��pz}�?M�o�m��0Lv
r���#�\<	����du�٬<��T��>�4,D�u���KQY��-������+tH/������i;��)=�d7�!�hj[�Uى�5l(|^�3@�����"���h2�e7�v���]�]nA|xn)�c�a�j��BO4�H,����2Y����M�T�L��7n���b�lA6������Z-�
ʈKPO.�tJ,8���u�r��5)%�,,��ۦ\�ؙ���&�!�����C��N�S_l����B��n��H.M�p��1��45�RAe�*r\@� �-g�gẗQ��=:z�q��q���ğ��n�^��z/SJV�͏D�{/�Ro.�DZ5I��Ig��1��Uf)_L���M�u�l
8��<es�^�X,��v��vt�(� F�D�8Ƒ&�dd}Lf1#_)��r�D�x.�B&)�+��<;.%��XE������bp�<�0f4�ɘ,y9��-J��+H'!�T����L�!QWx�>$Rqx<>�eNoTy�[`pX�
A�����ώ��<'Z�q�B�[M��J�|��ED����;���/Ο�����cz���/�,����Vo��Ʀ��38>U��P�}i$��[3�ˆ���W�	v-�L� �$)K�f��l�Q��C��\�ǹ	��7�؀r����7���ӫ'U��%�Z��8o�,�;���(g���_�)�wc̤Q�ԊB�	�� D��eQ+���#���m�.܄��'�oj�������ĳ�#�*!���QM:��٬�t���p����v�\ұ��<^�d˄Ҕ�3	V�,.V;�cvM��urNX��߯*B�a��Y�N���)2���+�I�'T/�'��m.ň�3�"L�n��_�y�y�>\�t)&�/�t�� B�cw����;ҋI�'`��H��=s��$|�a:q
=1� vѸ'<����r���"�� �d�ĶZ��E�1�j���. ��<�
))���s�p��C�,	V�P�\����e��Tũ17���	��j�:G�+5��Y`�\��|\�`!�x���{Ɣ��<yB�=-R?ݻ���դ�gφ��A�P��˛�A�*w]=��<���o@o,�L�nh.)r���.����hN��D1��qnB��4a_. !��c�"ύh�p�0��z��tC�e���aa+E��9K�5�#� �J���Y)9��(�n:���2��46��� ��.�c��9G "Ƣ�2K2�w��X�iٱ_�lfL�)��4mvyM��ڇ�^׌O����Y��sHg����H���IQ͎�]e�zwJ�"\2�s�[�8�{��s�z@D��xvK�'�JI
&n��n�=t�8l��M�K6@TFE�������Qݟ���fCS,�oÌ�1u���u�tw�O�>�M�f,�šc�xg�Θ0j�,<�,�.db1�9��{�9@��[]>=v[��/T'a�)���^��P t��d�8Z��,#$���3 �X�B�����(�B9r*�R�} W�svv�2�q��$7B���sq��I��4�됻�w��-�\>��R^��H9I4�x]r�x�Ydi�|n:�z0dP�C^)\��b�z�	X���N�SY4���Gd�c	!�
	���EQ;�QU��ץƝe9s���r��>9v�Ѕ�"�O���˦$r�&2s��R@�a��k����������w��eǟjZ`lZO�$[I/�w�g&��)���~�6u�u��rټ�Ej����ʋƤ/��@�,�3�e��YEQuFR�9�Б,��`��],,Y�-L��e�-��/��Ϫ֯~�
\p�98x`7B>��K�F���d�B���T]��N?�\��gP�s/�BW,��g�Ť����u芦q�y����,{k_X����]�D\��:,E���-�êu���8q��`+zx�Aa.g+"i0k$�@�d����h�tN�	�9^6�x��(HW��<Ov���4��#��xAY J5IȪVF>����SD�O�����ŗ��cǎAO_��<�A?��9/��O�xW�L���p��)%�z|:������(��F�[���=x���g
R{�N�`�J��^ݼ���X���'~D�)DxY�^�T` ���p%����Y��������G�J"2:�alt�Z���C�*�I�u��3�̐�>,��|Ś5�ſ}�L9�]sfN�����'�2�S�`6#]����Ǟx\f��&���T<��">�TU�3^T ��9�	��f�z�(T ���^~�L�y�RI؜j��ʿ��C��H�qs,$��I�����1et,�xC��p��L*��.�)ϛd-v�t�}	] Q}�P!����'��)Oub�E0~�G�����뾎{��=N�:�I�#����C����g����$9���{�C��ȯ͜9��@o�W �'�}At�5�&,�x,!�\�z�p���Q��UHp�hٌ$y�㒐ƄM���Sݮ�w��B��lm+�Ld'(V6�+2���i�-���<g<�D2���_��[�.�V���<���~�ƺ �����������X#[.��/
4}��p�up�lVP\�H&�T���c&�mD;:����q�n�(�Ш�fA2��g�ED�q��yOD�r\�C�V>/}�)�\�E�����UB'
������-���<���,�{i�ZQ��E�k�����VW	'�>�n!W�k��	�Cpᢅ0�rp�-�KDP�)�"Q��˂\���%Y����p���a��	�Fz��[�Ԍd6���(��24w ����壝�
��I3D.Hw/ϵ�qǨ,�(�%�'&ABX�!{���yH���8R��n��������46"�C�JA�����9oф{綷G�?w���ڸd��([=�9��>t!��	�/T�����"Ro�JF�פ����&�i3��͠�N����8$�Z�E�	B&1*i�U(�QZ׌@����3�A�(�V��u��X,;�E�����?ߏֆ0���/b������h���tWO�Vu<�$K�N�l۲C����_^�T�]�1o1���3��7�߼Ͽ��!/F�N	��k�����`��)����.���2�\��}	d*NtF���Qbǉ
�ȣ\��j#�B1_-%
��ټJ����(�A9/�<W���0�P�}毫��ϋ��BJU�>1�`B��t�J��7݀�SG��啘<~�u����    IDAT
>r��dr92YY
�"+	��3c�Ǐ1��a�ۛ�k�a7	��6l�s /���'�/]v%�Nl�:N��ϖA��nǚ7�tM�D
k����5�yX�Xm�d��Zb����YV� B@���	�RI�R)x=.A{XȈ��1�	���J(WA���jq��Ht�w�����){$��0H��z�^�e��W�ݎ�׋�\{-&�+���i5+��:���+]:����sjmG��O:.��%�~':�p���BZ0�o�|3�ǨQc��sϧ����9kچ��vb��I�]2�tZ�t
�־�L2!�
����@K'A���jQ�"���(c�LtG솫,�u�_��Dֳ�J�BW*��toz�� *c�2�N�2!�<e�8��7��o�M��K.��l֯��i3�������U�O�p�	��ύ��9mj���r����`Ҝ�x��j�f�p{��=�Q�I��p+5��G�!�o���p�"��� �e�DV
w"��}GԲ��9Wc"���Y�e��#���֭Z���FF*$s�`���BĄ_��mx�Ux������eҘPU��un����Å�_]�=�`����oA��B�c�`�Rn<�l	p�p"����lƩ�(<��
}�u�DK��y��A�R�A����+	�F��CM4R���H+�J�:�010�*2Z#�S���[�y�At���`�k�d|!E�[
�|����pɒs1c�X���c"ښ+�H%d�.��X�����=�4����?��G��j�1㧢}�(D�EĲ%��nb9*{4D�1Aq������b����= 1���"������9:��n��Z-�:�az[̄�j$􀽖�Vw�9'�;��@�w��e��ﻯhqcBϋFI�&�fR����rU�
�Tw9�B���|V�J�m3#��"텕�K��'s3Vw4*��<[�]]�{��,e��`L���ofq�I�Eu���"0i1���sb��I�����r��?�Y$�>ف�ӧ	C��	��x�*�F"xػ{?Z��P�b���/����ƌy���o���#���/��"�s�����Ǽy��bs�ǻ0b�(Y+y��~|���+�_FGoUG��.�γ����8�~�}]�(繀Q��	A�O*vv�	&f^�j'�U1�1��B"�	�<;K7�e�'��K�*)��\>��Q���?�����O��]y*�N9,�!&���z�g �����S�p�E'W������f�z�q�08���ឃx��8{�9��W.����nxf�=�؃\�w�l�sv�����ӋW^[��~��z}�m|�@ E&���d����L���V.���"�I�L4�Iy�G䉆�[��(J�ґ�_4��9�p�������$+�ϙ��#Z>�k�^��c����ݍ�p�_�O�܌M�6�� 
Lǹ�Xyrv�3�	�Ǣ}9l��c�ۺ�p#���"C�ß¡��p�����6w��7���Yg�����{	�<T��D6���ttvJ���cCYBB%?3�b!�j)�݂X<�B����fs��9)U�W�%���(����J=-��g$��,�3��\Ȧ���1���wq�o�C�c������.�A4ƥ/�"�E��.1B���9f�����6qj�)ȓO>���CP��_ ?�$��̓1m�m�!xi��8k�L��4����>��׋��m*�Hc�{�!�� ?�&��:e�#GE���S�6�݄��J�iH����gI�kH3V=+3�~-���l����Z8t�l��;nÖM���a�Q���!n�X���ijh@WO���a�<����V�����j2/�y�P�,N?���ƣ/�BӐa6dh�
����8q�$��S�2�da4l�h�lv�ڻ�ty��.���,Xg�\$��\�Jj�;���=�����Jm��i��]�j0��/AǄ�eH��/i%��O*��p#Fj�o��Xj|���0hp�t��{$��vݛoa�;����ꫯFKCX^g�D:�ģ';e�%��5�k6��d��$ѫZ�u4<*���S��,.E[�ʸ�����t�S�A%q�(B(7��j��6I���I��W�UJ�)s�x�T
�ˉ���ߟ�`�}�+��~�_x����`�/�����O���WJ���E�(�-���r1.���j���@k��7M��:C�J���8��+m�Z	I�lS���c�!�/�U����W�KX�t	�������an��71i��ݽ[�h��J�2��ۍ�A����%pc]X$:=�=8�ܥ�5ࡿ>��X�ˍ�/Y�??��&32�8.XzZ����Jq���1|�2T�'N���[?���.���l��c'`r�![&��!� �<�4��j��t�E ɢ��i,��Hw
��@Ʊ�Թ[��
	�)���^�K$5����%0��p�"����
��V�ӵ�|G���s�Lŵ_�
ɾ^?tƍG��Ȃz1�'L%���&���aР!�<n$���S ���1l�d|z�V��&ڇ�ƹ�'��:��T���̖]E�jlnA:W�K������ol|��nG�lE��D�Û	v�K <5T+�%��h��t�u!�)v7Y��.jΩs��@�J�a���Ը�:	P����Kl��5�p�e��\�����}6���3i|��#44�j����P*��3��H�(7ߥ�2e��>ݍ�6	��
n}�)q��K�/b]����v�e3Y|�w7��1\�������_���H��t�"ƳM����^
�%�֊X�����r��)�G�6)ȥ����Lr�ܫ��ĳ�|T�^�n��sK_�����<a,�Ϟ��V>�l2-H���«��$>��&��N�0)��6��6��`'N�B8� ��_|��B�--X��{غ�S�w�rL�1?�0Ξs̵
ϟ�'�+�ٗcѹ�����J�n��V��$�w�S�-	��k�Fwzh�T'�,��9Sg,�dR��j�e�*��
�`<�B��K����D�A�Id�#�˩Y�\�-7߈�ﾍ�V���Q#q��bX[�p4���8�lFg$"z�t.��jn�TL�1[�}�X<�RMCc�Hl�� ^z����Cڰh�<|��^��/�7k׮ż�s�c���8Y�SA���GX�y��6kt1,pi��֐(A/(7�0�*bÚ�'�yR�ϸ�$�����/�@�`��r�Vv�F�>�1O%��,$�'���_CKc��d}����aڤ�Ȥ�B�en�<.<��38t���r���rL�8�&��V�7֭�O��E�/��Y �&NĐ!C��[o"�v���E�K���N�>]Ү�n��x'�u��q�@"�&���U]vK4Q��'�R7�z��|&���.	ݯ���Bw/]8��u�q�%��:��l�6�HM���MUUi��%��9��*��Y�J�&Vlze���P�gQ�3���1C�`����e����N�q�K6�/�z�8	�Q���4�9��^Ew_�`�kW�"=`�Wҗ����k0���ӽ"����Kq��ix�7O��"�����o��Dv	߼�:�>ў^twtc���?i*�����L�����y\���E��p�VD�z0o�:B
�>؆��VL�2E���+_@��C�ǒϭb�F0ٮ��PɊ�&	p�Y�4�����<.L�"e_���E!8Qv&�d������nZ�ڤ�K�\΅K���d�pˏ�/	i�ߞ��Y�p�����i��"�O�O�M&��z}�v�څ@(�Qc��?�P��1o�9ر{?V�ۀ@C#��xх�G:1��;w�����Yg�þ����z�:\����������6��f���R\��C�r!�l�;�U�Q��o*�#b<�Y��*,$R�*�e��+ZT(m��`��.lzs߹�mk���+L;W_�^M~�f����A�g8�fP��bhkn�s;N�<)��̙��s�.��u;&̘��\�j�<�4lN���5�0j��z�}�)y/������o{�	�>���"����P�XK�����i��]��+x]v$c=���p{Of:t2Y��(.����Z'��W�.f[��%�2�f�袈�b<D�����sf��'��b	7|�ZL܆��	ǣ�����H4*񠳻Ç�����1t�Hqv[�j�8��D�4c�~�/�x��8�/�G���ݏQCa�ԉ�Էmۊ=�����>���vL��O>�����f\l�H�bC"F<��k���[F4-tYq��)%��G֬v%Y*S�������=`_��r�;�R:DVē�e��o_'	��gެX�h
���'�֖����{}ș+�{4�qDz�d)c�I��{�A�������{��{�I�q���.��=�&N���`��^-���,�U�+_}M$��jٲJ���W�c)��I���.!�1����K̢~]P
�6I2ӓ�@͆�,	���E(9���	�;�ǫp��!��o�=�R"����'�5y">޶E�qBM�eS�W�+�7_u] �b<����9|�m'���X��f<��3��9{�B����c,;w	���D���?Q��X-��˯H��1����V9"�*����,\ҍjd#��j'��{g��8Ǳ_B�������\���=������c�fkgB�p٬C��ɺ��f�B��C܅�?�Sg !D��� �V�cD{.��|��x��#W��6^_�=}Q�]�J��������h�!��-{���'n�W�����$���6c� ��c���0c���ǻ����U�����X��Z����0f�Y����
������];v�QG<�����KfM&�C���\<���K���{P�f�L��6K�m]�,� ��Lg`w���{�=�ٿN�C�Ƽ��笝�#���s	$�O�.�E>��ٳ�aƌYؽk76n�(]v}c�����l��a�Zu泱���g:�r�$�2�Gm�&�Joz�����+��ډ'�xK�����c��M�0ffϞ��Gذ��S}1��6_�����"�[���(�,���_�����k7�4�/]�ǃ���{W +�(p������K��R͌|��gW��#�N�ʹ�ݎ<�e6MԨ�(��t��&R���t94��wP
���"�[ ?�e8�6�,5AUH6�f�[�2:�&�R��P�p�V¿��6�7�;7|(����ɣ�@����^��g���O*�>ݵm-�b��c�n��T���fã�=�D:��}��0u�4���;�=�����{���!Trd����*$�Q&������2*$�U�r��ݟ�ZA�a+�B:�xO�b�Ө�_��/�I�d�	�tݺA�U!��8�<I=j��C�G�ѥ�4�L�r�'O��?�����s�����¥0��b�B��:�HȎ�#G�J�N����Oa��i�y��=V��Ł�on��ݘ4c�9o)�y���4˼9���I,_�\>g�/�UkV���`޹����t	�AKF9'�Z�&�M�[�,(\,��K+Y�7��K"��J�J�8�B���.Y��s|�g1J��/�"�I40��r�p��n��7_ú�����c�Eh	����w���tL\�a��/�D"��p�T@wg�$��[?��ՃRɆp�Plٹ/mx_��5�	O��_�(�C�eRGt�����i��_���Z��ǟF��1���rM)=.�l�7s+�\�X6�I`|�=H8�]$��j�J��KNuR��i�vI�(5>���%	��9*��`.��xs�*8MU|��+0�!�]nC0��7��u�/2iCs��Y�M�0y��!̜<�D	۶~��c'�+��)P��>ľ�1d�p<[6o�5W])�`��'������/��ACcԸ�X�z���noBg�N	�2fS�� C�Y䶈�J躯
Y�ʷ�
S�֯�ؘ���^��yv��?�����ے���slueե���}�jS��V�B|�RjA-�����y�f��s��)��'(	�б�x�GE[Jf��4�?n�)Z=ؿ��P�ǃx"���V�X�:y�Y��ۇX2�"�4�]�+H&"���%�4z���u����c�	y��D�=�%c���������KJ隒�Z�a�Y�0t�H�9N��Y�9�/+�Qm�ϯNe�
�7���TJz%x�V${:Q���m"۵�]�x���a��ihk��/��}���Q4�4P�>e���o���X�����{c�����TN6@Q*'���k��(�CT��7^���n�3O>�Esgc��!ؼ�,9g��0�i��T�v딤�������n�z�5�[�Dj����,�1�2��}�x��\AT(��RU�:� �P䜩Qٴ�%��|�8?/����*L�BV�탳ZĈ�F\�����>Սӝ}x���8��O}�DC�F1����^���}*5с��D`�����w�Ɔ���6X�!I�d�"3Wdr�IU��k�AC �������[n�>�򁼯�.Z���6���@�1��S�fYD'(��<����l�;k���@w1�i�z�iTM\����,F��gN��t*��7c�С���䮞��8$ω��j��L.��KY�����լ�O�������'��
2@�C�N]4�DnZ̉.<��J���7C4������"���(��M1ʅfO����������4���X<w&^��JI��F(;Ȯ�Zc"�����}}Q|��GX�d� d&���؂G�z�{B�����F}��G<t��t�#���ގ�׏P�{�ĊU�Q1k�g�B�������r(�"��s(��phK��u��JH�i(����ϗv�ԭ�������eM�1ӹ�KU
\�I�?��l�
�M�5����݅��=�WW��9�f���.���F��hi�G=G�4V1���q��#�:BAU��ڦV��w^Gժ�axq�z���1�u�wpذg�ǘ1c�4
�'O�ɓ�1g�ttt���w�n��	�ї�`Ś��s�ьՎ-�mV��f�TW�Z&�tO7}=R�q�������Dgb鴠�|�%�Dp����`�W��˃��\� �ق��ȝ����N�v��Ez���݈���8��w���L����n�i��Y4�����*n��ر.@>��%<Κ�=;�a�ڷ1j�4��nT�uxu�&��b��I�7gV���H,iX6i�h�q�ÿ��&�ٝ0e*6��re��\c���"��%a&M�a��Z��oP���D��:b�[��$�'߸�����P�z�rBQ
;οK�"KS���b/�L�x���{�0�6��ʋ�`��1H�v`��6kV�?r%hxsӻx���R����~7n��Ԍ��Kgn�0�]��a�u8v�?=�5y�U��@��Y�0o����,����J1�hm
�,���4�g��y�fY��k��i"�����m.!i?ZچH�5��'_@��Y�v��,9�1�7�Ȥ���D�t��%"��
=����YS������	����_�
��|=���eYJ� $��t>��}�HC����:@��lλi�N;	^�C䖋��Jh	���-_y����6JV��$g�vu��I�"���D9�C��G���@��,J�;�5|��?�VB���K�7�gm1�H�"<v��L��\�g��"��'�7Y���oq��7�,��ʥ0�!����]���;n�<x�ٕxn����5����=���|��(���	�DM�Zp׽��o��E�u04�W����U���R��˯��3���/��2f4���BP��&�����L֩��$��m��4�p6b&̙�7����?��l�3 �&�m�蓌ȥ;�x^�_�^"r)������T\�54n����(�=y��b���m;y
�G�Łcǰe���%�	�EgK��%g/�yK �d��$�]$s~�k�����Y5����    IDATQ�iH�*����$�r\��Ĭ���}w��'8v� ���K|�N�Ĳe�D��{�╆����	&�����߂!C#���HW7�L��G�^�O������u�����=h<�C��=;y�Ĩ��&�|�F�8z��9R1l�bh���J�b=G�ÉNΚ3C�>�Ou��n�lH�bB���.fL����&h�<��aVwo:���O�b�J1Rer4S��
)4����/n��WV�����_�Eb�'��߳t�b�<y���Qh.'ʵ� A�ڶ�#ԅ
�a�:`2�P�z���x���=y2Ϟ-�������O��/|C��Ώ��㏶	j���&gu��oa߱�����&/�+���J��L����*�=z�L^�͍���b��݃".��W�@�V���i���mg���XCB�9M�R\��GY'�*�
�)3!�D�_��j�:���/� �]r1��:O⢋.�3z�̈Z{wOw���G����f�9xc��@�jF��+om@_2��'`ᜳ�sǇ��`�;�u0�>]@�Cj6�����;�3AA��KQ�i]�[Y뫚���U� (����s%����R��K�O���������?������6������Іz�� ��]c�$�h�$����]D�"����;�0��9����~ϐ|w���r��q�]&J��{��o����=U�j\m��,��G�o���&�E����1�h^!7p�I�H[c��M�l�����.�ˬ��j���jl�y �����dd
�4n4&��|�M��ٕwAYyo��λX��f�ʠ�����P,�$`"Cy�2�6�.�M��b<B�7�}&��ܹ{���8�_v�xt/�*�5;9ž�]x\�J�w��;��@8k�yQC���g?�lA��:���@��=f�:R1���i�ǌ��1j`�ܱݺwAC+�]е[/�}Q|��W"���0v�p\~�8q�
���2T��}!��ڛh�`�͇JoF����m�d�m�n'n�{-�d�7�"�� ��Pd}F��7��onmǆM� <�p���#Kd$�h~b�Z�TCKE_"��K�b׉�0�r�N���'@8��!�A���s�)�2 �-t6B!��DC�#�T��:�Y�Ŝ��㆙8u���y�;�p��9�t�{�-��+�.���"����uwa���Ҭ��#	�nl�wo�)̹�08s�R���D=Nb0�I��kf�o��ذv⡀8�雯ʠ��U"Cوt���Fr"�0��`1K�u,�1�ƨQc0��)hGq��_,_�xR�XB�"�]�؄�L���?qOdЅ�>�iI�cQ��X�7�"�h� �:�����;~[6mDNA��d��ǅ�::vF��(iT�'_�9W���ӧp�M��(�1��!����CR����A�k�Tٓ��d������&��7_��{�y�����8cF���\R��_D�H&�������$DZ6��>� j:��s�0���'����hECS�Lk�XX�.Th��51�0�4E�\�:�f�Aj��F�b	�Q�]m�c2C5ʋs`R�r�y匫p���x���ص������t��?pvn���*�O�Y��V?���x湗����ww��_L*��4v4���c��K�`�����<��(��C8�cv�^_ȇ@2��)C."~�1��=6h��dJ�XJ�u;�`��Ș�0�4r��aÜL���)F@� h��i6&��&y$�g=�&	�A3R�3nmF�SгC�ü��dMu���^������N�%��6Xq���;f2�� �F�A��Lvv�;���vɿ�ds9�������p��:p��sУ�o���<M���k��P�Ê�sg��w���RK_�����6hZ|�n�N���^��JkQ�g0��J�r�Fx�J��Е#�	����In=}�4�K�P�C������{�0�*-�.l�A��0*5@1��������lXTgA���T���/��>^u���5/���p2-V��C$?�;�4ŧل+�������D>��$��܀P[z�`Ҙ��{�X	#G��8����V,��+�4�	<�I�i5�y�`��i�<0�ho����[PU[����Bg�A�/��n�d�E%l�0�|Z��p��P��?�!qLϩS�����h����O<���8��);O1�/=�3*ax&��D�Mt���v���E��E_w�0�qN'��V4�d����K��{`��0~h�0{:����h?� �CO�ؑ�hljE����]Y,��֛пw�"�p�dJ٩��/�����WQyNj��J1�`�`*	C(�qbh�>p�5�^�A��E��jj�Q�� _�'{�!��k�'6�d�s2 �KK�Wb
�<�&�$�g�vY�i+�-�j�U(�-,)F�I�S���]��$Ȥby�	y�Ť����/ȷp��i�B�8���+~ܳ�-�:�A�����w�?���.t�5H��՛��QԵ'^]��\����`t���
�L�*�N�4I�6nƍ���$b�XYh�I�X�V�n8| �V�چZ���r�Mp;Dä��ͩ6IS��եшo�nÚ��j��8�jP�Gm��PIr#Y2�(�,�L�l�f1��N���dV�ޚs��C�i�<t�h�����������D��'N������R���g���\�o��*�&���p��9�6�x
���@]�e����g����}$�!��᱇�����Pu�4B^�H��H��`�H$�s���ԩ3��wzii�4Q����~`�%�@m�"��-鋯�_,	��*��?dI��zr�j��� ^��4�6;ڼ~!ّ�C�Q��1�D��	o3�wC[�a�s�;p� \:i
�[<����;��6		:��k����^����?�������7��ѓg`�)��Y ��Ɍb���J��5ǆG��vmۈ���˻A~��l�R*Gq�Ymi�Fi�	I3_^\}�;E#	<����lvCmv`��m�v�$2��b��$��8X���b#D����0*��͕�h"��'s+�>�iP'�ȳ���u���r�<t�/0����hʽȦ�	�w �7�6ֺD����6u1��+�d:$v�Q�m{���{����]�`��.:�R@AD�:�?ƌ��yA�s����Bi�"�Y�TaI1Z�aSPd�
��OǱs�4��#������1f�D4z���bɚ�P�R�l[�IǂR���\A��:7ND��#�xb-�F�(��\���'��Y��l����sB'_�z�!�,����hBg �����й�����:qA��:EO��*��);�s:��p6iU�5#���E�>���C��F<DN^�^�.�Z��*�Q)0���x�'��vH�ݾ};���_e78u�5��X�~������Pv��\$�Ń��#�m�*E:�����bV#�LC$%�lq�+��銭lF)J,آ���%��2�Ƶjٛp���i��iG{j�ly.j0��l(���:F��Nھ&C1�n�y.J��d� |�n}�%��(�J��A'�z�������T'��;v������F��<?����J�{�� :3�D#���cԜ9%�#��H�W
�d5����dp/��.�@�'�@o}3T)J�J��x�y��b�� ���[�2jx"ʥk69��ԦD-!�k֎H$��-�_V5Qr�@t:��c��Zn��>�kz�eEb�H�����{Ǘ�V���#�-���w~�ԯе�)zl2���*���%��ї��K�VX
�3푘�	1P�A3Jӗ�%WJn��x.�$Ց	�KG�/�y9B�E��nq���O�\��1�I��o����F�v����Jm@R|��j��z�N�F�A���(��Ҫ��$���HY&!d���'�M��G�M���'����1#Q޳�up��a�}���]EBf�JA�1m*.3F���y.�|~�,μb<��`���p��̑8фZ'�)��"��;���=�K��$Q��|�(Lv#�	%܈H���@m�[[1u�TA4X���0s]���=1X�Ź�&�\�#q��}a�4-5��H�DI"�[Y�ͮ�ƉU�Z#a�w�i�{�	)�Z��fs���݋�3'0q¥��� y�k�m8q�.\(�r[K3zW�㓏>y��fQ2�ټB_("�v�Ћ��"��G��0C߃���G�B7�͘��]
�z����SZ/3 A�#~�>wk�}�`<*Ĭ�'N�����@����
5�uF��ٗ�ph?ܥe��LN��V�����DZ>�͊��-B�j�I�>�˴qh�����7�#�Z��o�����OŨU���ըUhhj�?��(z~N~{�W�c¥cp����i+]�؄�����P��Eq�^��s��hE6����>������5r��^�'z��� w��bA�6:��E0��QX\ ���A:�@��*�3WN�i�~��|��QBŁ��a�y*�Y�M��`�&f'l��������E+C1m���AAW%C�5B
��	C��:�L&����+�9p��o*��b�n\!}��a��	=[�;w�T��;��<lu<�������'���>�`Щ��<d����<#V�Q�9��n�7_/�3���<�����lw��[9�۽�Gg^�F"��HMvA$N�0�O��1|�P�4F��`�%e8z�8֮]+p����`Ҥ��`1�/���j��H@Fk[��;���U���0��+��
�붓��Tu)��@E��)q��"QɒIH���H=��_������ ��ҥ˰i#3��B���]0�~}+�ȃ���ɮ�˯����ѵW%�^=_-_%лŝ'�yFeB���P�ݤ�2�x=�����x��:	ʪ����G8ER�N4�т|W��"���XK8��No��dC0��U+��A��d|�z�0�����otg�V����=��R�_�D]L�o��F�:k����:�̙W��Ջ���x��uDoT���Ч��=cz�nٵz}4�I���>D(��v�\�]�w�6w�Dg�5��i�ωM��-r���sA�݂��f؝N�:���~��1�p.��@����dz0�ܨjjFaE���Q���O�&��S7M{�ν�V-�?5��%~�lJS1hRh��h�����~�������r��������
�������Y�P�~�v���_>,aA$�1q�o�x�ǌǲ5ߡ��'������	aZ̦�b�C�y�ɌL4,�&�5�q��I"�����φ�onA���:ӷ������.�N�F�8$uVDx�4���"_�9�iH�$�Z�ϡ��H,ͦ��Y9��F"_*����ńa�����'�����	E�d�۰}�N������}��ӫ7\7O��Wϔ���V8s�p��)���{�ihA�憺�;f�i�����7j20#��z��n�ʆ&/d}�a�[b\Y�$2	�>_�3�Я� �(��F'�)2�4
r�X�wNZa�x�0�&ڂ!8MN�i$?�x��+��{==.��PT:�0��W�D+l���L�H g����BE�B�8�W����V�덦��a1s~����o���o��*���p��<��J|��d�����g_�|�FwL�<q��l"Aɹ� ��޽z�Hn�*#$a6��` 	"�Z-��;�l�2���	�g��(+/G8�\�1��5z�֥��{�4��? �6��'�|O�u��O,"q��.ө����%1[�f�+�b�b�X�и�� �wN��Oq�?.�0������d�_~����'��Yo�qrB�!��o.;�O�.P������lXu&!��Lȏ����-hS���q�Q�Ђ�B���P�f�$����3L&����ZS2���݋��R!z��N1�syH�x
*T�D4���g
Yi��%�XӫG<mmB 
eR���g�~1G�.���+*{��S�L��U���V��*� �7��Uk'������$��������x��[mɩB��A/|��g�!��!�z������ʇ�l�Ȝ�<���Ņyb�����*D��4�z� �1Hܤ��@���v'�A���C	�ၸ���Q���`�#�n"��LQN3��\��b!�G�n�9�Jt)-E$���gZUuN�K�Pܫ~�|%�5�J�c:��}4MIĎV�I����C�-�8ҡ� *�EY�pJ��V �m���<��Q�!�e�_��AM�+���ߒ�93��Tuj$CA�����|��(*(Dk�3����̑����.��D�J�/����,���RW�uǐ��`e�9�N�|�v� ���:=��ޅ��o���qc� ?'Wdoj/pT1F��`��Ù�&�m��5�?G.>+��x噐_ �v� 2�� �s\!�e��ᄬQN�
�5g�|U�k��5j��Kn]��idE��
�.��y��	�a��!�p�{��8�)3�ƒ��*���Px�:�QFJ�.%U1����6F��5�����
�D���F����Nx�$&>7%N	��N�"�GlJ�)-2z+�5
$���]���^��$�J3�ВLR��������f3�p5H�� �ބ�ݺ���I
�}�݃9��!
�S���#���#�0�@�̊��ޕ��?</iy9�������p��E�8y���bh�{"��JAg���=�c~E�������Z-�eR�D�����r��po�&H��u�,ǝ8et��Rȴ*��������-H��v!����Ԗ|N�4"8�UjiY�.���Fiq�H������7U᯿{�T���8]>��Ө��^?�����w�r��%ԨϘ>M��zW��u�]'R2Wn��`?�l1�o݃PF[Q��$m�y��JFż� �����'-tل�S.��!�8�H� )��()t�q�#ʖ�UU$/�@.4�c��$e]�����N4$��̀"���\��Y��q�,�Y����Y�WbpE�&G������� w���s^�v���c/��L���+��q�ԟ��|�-��ςީ$M)K�Q\n��T��S=I��P$B0�S��:���f1GY�ݝ��V�d%��Nm5:������;2�����y�BJ�M(������`�I�0}�����K�j�d���)�c'�����i���Sg�u�:/�>�}1j�p���a޴䝨�X�|%zUVb�eS���o�U�/B�Y��Ĵw�f�e4v��� �!䥓�I����`kr��Ch�Q����̸>:��R�@�7�O\�D�2����"���h��Ce� �Vˤis�#�Rd4<��I�������#�^�)Ν>���P��������-((��f���{Q[[//m~n�U��M�Q/����݁�f���7X��l;r~�h�Tĸ�lt)e*�����L��M��:��A�!!����æ�C�BKL<$���Ey2h��l?��lݾK�\iOK�+Y�=zb���rAщ��Ⱥ�z4�u��e\������@$Ik�h�9�)�#\w�5� v��#,-�&�h�9��ɨ>q�4�|�L$�̛w-
s���D0���6M/�Z*F�ā�xi��0s�c0F$&�r�hG�%�	Y� 2�%�ia�ݨ�S���J�L$C&}2$�OS�i���������{i��;�_6�Zq����{e�[�A���)��)gr�O��`A�dA��)�E�� ���{w̙~����G�e�����iGL(���o���߿r�U�f�La�S�*�3ɀ�2(چ�UuX�v#23R�b�$q�*)�B��̛����g���.�m���?�&�]���0�C���dv�Q��>}*1d��n)y]��b�u�^V&:\�P{߿_1�♥<���as���c8W� �� w1�Ԓ�t�z���X�.��E���i�5��ӏ���x d �x�f�ja��Qѽ,&�<'��f�Q�e�g��ђ��x{3�n��1�+�D�#��7`s*q�i��řQ���Co�US�ń����cx�rTt-��SG�P{���Il%�T    IDAT���_bm��x�װu�v�wp՘ Ң���0�����p�n�V|��*�k���WwY�I��E>C4,k/~/1�I�/l��Z2���h�Q�*���r����@|��YlVYK�aR�J!������@�;wWR$kg�0e�2��tI�%�Q+�`kS�bC�uq�Tj�� 7@ȿ��`	�e�����N'��NR����^�1����N7�=��N���'tE��y�p���C����e�H��BR�g��;s���LzI�����#F�U��!mF�%��
ÃEe�>p�0\}�,��߸ޡ5ʡ���� ���;oE��X�ŧ��y�$�b��թ0e�d������A���E/4�w~�!9x-M-Lr����EIi7o}�0Zd��HT�Ӊm۶!�a�ȑ�C8{�,���;v���L.���*i<`0�!�FE��E+�!/j����������yO�����d+�^�'���'��X�HXTi`�ؤ�k�V�� [^�9*|�2�?�L�R�T
yN^~�o����z�p���7s��	حc��u8s��H���'�Q�9
�.�H*!ų�KWT�/Œ����o���a��a/(��"���/�P(���B)��xH,ᮞ^�
Y���1Ҳ�Q�2PŃ@�6U��r&#��d�O@G?�
I2��L�Ŧ�]�UZ&����H{����� �����K�ms#A"�I��{�Ba����Ia6�,�55�)�p�998]u�v��a�I�WEO�?��y��d��D�PiMX�i�]=��"����ֳr���b�����VTv�)p4'z���1�����L|�D��y�
�j��5]@I�1_�ڴh[�L(���wK��@���H�[\��XK�Ѥ���21l�P��֠�DBc@�<��f������B��i�|���bD���.dK^�p([۶m+|>?�A?����F K���Y!��B�=��°�#�n�KN!���4��]}#�;�;�4��Q/���?�j�d6�;�`B�@B\�TEv+Zj�ĸ��8N�]�ѐp,,�E*�8,q�!jς�T��Y��	F�߶ �!iP��h�H��Q����a�B��!ߦ�m7�B��\4�UjHc�\��W�=���v���-?� �f��;�IR�
&3LN���K�G�����?x�/@g�AMюϵ��U8M�ԹZ��/Cv:�~Y�"W(�R8-���d���%ׁ��'�o��ݐA��$�ߕ���˕X"w�M͂(�}p����۫�\�^S2��O�CG43Ss��i4����s�c���ӣ��������� �rA��'�a��o���k@yEoL�1C�Z:V�;+�${�K�p�i�� ����%��ѵH:��S!�1n��b����N�픬u�ْ��ЕLy��*xgA�+)'t��w`.m�WY�~��I��UZڞ�f]����^U�1����O7{�N�6)��*�8��VKHN)���AR
�Ԑ�N3��8��C��!]8,�Y�b����/��I��j4HGC�	���iM[K�c�t)����q��Y>yZ"h�"d2.�˥��{�s'�a��~�(ַw��\N��_1�����}�^.���'��c�d���"�kh�__x��\��n�0���(���&\&�^�p��	�ܾ=�Ν���ݻ%���c�B��`��p��J�
�I'��1v`��O��	���a��%d��9՟�7�Ah�I�RzS�&�66������f��� я~��4���f�@!\�|w--�#=���/��jF������P}�͝'���=�u�.&,|�H<b�JC�ᗌ�y�����G���ر� ~���b͖��~�N��艑c�"/� ��Tɤ_֥�|���_���F�}�lv�x�9iq�N�LE&��o���g�a�R	��2N1�/�b�͗Z	? JV5�:��l��*q"��B�#�V'>ϱd�o�I$M_|�m����M����&³O=�h؋o>��ó�յ��v8�c.��+V��M$�f$�b�(*z��-7܈`{݋���kbi-����1a��hAo/�3��v2��@���hA��R���
J�7j����ZJŰ�2<�N����܊.X��ّ
�p��^8�Zh�1���LYnG�ci��<�<ߢH ����b��_)��hy�]p�\���V�<s�/��~}��ɸi�,��?`Đ!�v��b����+����Çb���8p�X�h�UW]%g���믿�Z���>�����o�|*�{���p;lR��T�$Ұ8sq���K;�
O���l1�i�y�&$�c���">�&>[e�P�hH����E�=4�pq���g��,T:�}q-��`R�G����RD���5�ކ�.�x��g���e����q�]�p�Ο���ic�T2�����A �Å��A �����d9EE�|=y���E|�z9��=%}Z�\G�|e>�Z�L"yd�K�������%�_�Cj�����v��iD��0�jN#��:��|o8��9���8���%�>IR����M+R�m�Ml�܈9 ��b*���}b#=v�plZ�~O+�\N!�c��B��.��6l��*-��ӥk�&�\���͕�h�D�]�Q����C�'"l����V:?2�:��i�(�g��BT�TB�u�E��.wV`U�����G)��$��b��V�C�DD0�.��]�����G���zmm����/;��}:�5�8�KA%�$��nR�^Y�E��s�⁧�<�Ci�=[Џ#h����l�j�%Vx�E4�W���P�"9�i2�R� �N1�a*T<��~�K�<{����͕'<�y�P�>o�����R�Y�\y'��ѽ+z������e��Q�S��	���N���|B��|N�>���H�KŐ�X��pv)���S����1t����%�����f��ѣ����~�U�f׻c�N>zD�mZ�r/����Tf���p�$���QdFzIQi$eBW|���0_�aGyI�sM���h�"q�H�������[޷�L��/_(����$�%~�Kq!n��z������El(�ΟW����¾}������9sѳ��?���^���
L�:Y�#j���_��7��k�}?��/�џ	<7�y�@�AQI)���q�-�J�VAq	��Z�?m�-'G�,�٥����#F�f2��������5˰s�zX����jB.^�z^����L��&,��s*��@�����E�6O �K/��n��\�����V��x���Ɏ��w�u2�c`ʤ	��Z���g���zSbSo��N|�h��.��2�۳O>�k��i���_~�����qխ�"j���_.��������z�j�7�Ϟ��s�"q������
!�>ٜ��b�G��V���&�R	���9=�/�mZ�߯�!wN�C���w&c�<PzDf:����ِQ��7������o�s�a�v$�9iu�#Ϧ���
7̙��|�)�]�>y
�a��U�4i2������A��}��iP�}B
i<�i�&>���^yUt�F_�,�	�%e=1z�h�2�[����W_����]!�8�a��"
:#*"���w��JνU�B{S-�m�"F�x��� ���=$+{U���I+�-~ʊ��8��&;����a�*��Cw=i�h����$/����v%�ڏ{�@�;��/�?�������U��@*o�ʰ82�+a�[��1t��9]�W�~�������uX��&����9cC��Ϩ�%DC��T��Η��4���q�Lۋ&��g?��"~��-HE|h8
Eyv�?hq��f�n}��I��r��<!\"�4�1U녴��񋳥���	-�0�r B���w�0p�ܹ��^����QÇ
1��qt��X�1b��f���p���Ί�dа���,�P[-���S`��7mEA�J�s	�~�є6��F��ɉ�������q����(���Jq��.����l�E�޹BS�M�b�ϱ�1���������_�m��-:w�,�ʄΝ��KB�]m��$ĹlA�`��".K�gO �?Z~q�i2��-Ck:���&\d�w��t��K�)ߴ�L&q��a�}8r�<�J䰐DĨSa��Q�Z�x�Z>ù�'$q��w�EII��t��NO����޻�����MH�����^��ӯ����,E��A�:y*��&F!�o-S9����2iX.���xZ�۰m�vq2� 7#ł��ઉP{�oߊ�]���)-[eQY$f���K�b��ժ����#C	�^�D�Kz|A�8y
>��3	 ۝���h� '7̛�M�	����

�
��"����k���K.��z��P؏cGa��s1��?v�4��qd�Q47�����º�[�n�v<��#rY�ܴi�$h0T�ݻ�����}�Q�֢a*�6W�6�d�M�Ìۮ��>�g@�ˎD�f5I�gAWg-d�Ϧ�r-���$��1�!��K�]6'�@,	�Ŋ�~\<�����$���q7m��q��W�"�c�a��hm�C��EA^��'�)�:�pX���k%��o�N=&0���Aر� ���{̹�N�F����%�Mx�w���8w�,Z�pݬ���0:l�n�v|�z9�
r��F.����4ױa�}~�-&�v�l�Z��÷ˑ�P�"�뀚je�u��Ia��@$��������<r��,p��׎4�",�3f�Ûޕ�2���[��Ť��}1l@�ݵ}+*�TS��}�"�������]�����^xA���GK�	/��gQQV��k֯GY���0�����g�(̹�&�[���yH�{��x��8{E]���ߐU@��i�;6XDM�3}8ճ��0z&��=?m���Eq_��S�����}6�</��9l��vª�E�Ϗk�W9��2qƓ@ EnaZAdt���4��$���w�H��g�哦H�ơ�q�k�į���vZ�=��������~��*��.t��O�`٪o��3������A\6�J��66�]�C5���ޣ>Y�9�N�!V�[w쁚{sr!xn�F,��S�H��sc�Q��5:yx/~�~��p�]�O+����f�/4�)��DL��gW��Y��9���VFt��C�(!��&�"�����ǀ�}�ڋ/`Đ��6�r!ű�x�伽����k�]��݋Ғ"�2q\9}�L�DF
��I����c�E�q�d�J����@� �+;�DG$�� �#��
����H�U�TH�!���%�1��/���N��UM��� ���/tm�׻8��F�ygxeq���lm���p���|����2�Gɐ��]�])��c�2����� �$2!�h9;z"������� %E�~����b�y0�@Hז��^�#5�`4����cO������G`�e$MS��qL&�sg��e���_� ׉��j8�6T���#/_/[.E�fw�����R��c���|�eX�`�@�cǎEQq)^~�5L�b�{t���_J��̫f�������#G�o�^\;{�|f�OS#ZS[+{�#'�� �;b�H¢7#"಑��p�4��܆��dD��5�NT��=�$�lƃ&�ov�Z���9��TQK������F���2\2a>��S��T�<O�tޜh�%�f�r١����k���?^~A�O?�;�{����%�}Рؿw�ͯѽ�?�p�1�FT����C'�ؓ����k���}������;��kQ��-����ܳ�c��زu'J�wGms�t�g��ђ�CO�K���z6�[��;w"I>���TYB����t��C�4�X�S	x�!�q�&$P�,2O��r㖻����;�e�n�k��h9��`&�Ɠ�����iƏ%�gNJ���w݉����%����Q�-���5(.,�#�=��{�#�WIΜ�Ŗ�1��������>G�~����w+C{K ߭^�I�N��o��K&^u���Yc6dC�eAo����	q�s�o����!��Q���;x�{5v.e	��,��#�N�9�Q����v�¨1"�Ⱥlب��ٻ?-�F���������b��1#ѭK!���	�����&��5�M��k�q�f�X�R�'�E��TWW����� u���1n���(,-Ä����G�����?�uuuX��+a�O�0��}�6X�x��̇�Q̩��	ӱ42�4҉�L��V�K}찡1�>������T�I�jf"�Qtj86��{���=��k&�vlB�,��u�@�H,��6/z��@*)�K�5CCw�H\!	_�s�Mصe#��E&G��0ѭ����Ÿ��g���I���z��z�Q��zx�~��Z|�h1���q�]�cզM8T_�֎ �=sgL��u[�uۏ���C[�V�_}���7=6�OdMJ&]���3t��07Ν���e��oj�I[�ՄL�C��+%��4��'�cygek�Nn	�,�\��N.�m9�����ɡ�i3��Í��_���ޕ����SЫ��^�9.�������>u��A� �墶�<��z9�͸J@:.���ŧ_.����W��}�� (�&\�qCFaŒ��i���@S(���l߱oXH�\u�;����V(��DN2��_�*����R���9��̈́�?*��<ǫ��mu����tٳe���	�1�� �����=��p��0���6�+]~a}+�$t�=v3�C����]j!�5�/ #^�x!{��6?~���q��I�>x=���rI��B!�q�M(�s����$I&{����n�{	���0{:�v2���(+�ƅ�޽S.6`\1�J,��	h7�
���h�P޵;

D�u��)ģQ	H!k�ě^����b�r��Q��苯��]Tv2�4zZ.����ېk��~��,�L],���!�����#�A
��V���9���c6b4&�#�4'�_�Ae������B�J���'�~�J�?���.x{�d��1��Z8~��}�'�� +���e=1}�Ԟ�ǡ��1�۰��u����ї�y�k�"���y7���j�K�,EU]����%_j�%ğ K\jע<q<�a�
�8�_t�Z�J
:��|7Md�f���CZ!�*�hLvpD/�GM��藥�<���e�v��X�v6��] w�悐q����w�=��ׇ�V-GYa��GD��
�q�/����Бð8��ۭ�ި����O?��˾�0f�(上�q�})B?��}�l�����.\:v����Ũ�7��
���ش�E�x�%zؙK�XB�Mi�jḬ(\�46��AGk��_���NߒH��ٕ��
�2�[O���\	ˈI1��q���貺����9v��/��^��(�����b4�\����1w������У{��v=v��x�׿�IvժU�ޭ�4ݻ��i��R�����r�*��_A�w6�CF��+�}GQ\w�8t� N<$��G��/�m^̾�|�d	��;fx
$5��`�J��,��׃q#��[�}�L<"�Y$�G��ʘh�$�%L��!w�8�u$�Є�����RRZ&�Vm}��޷E#&I��)��)���A��o�	�V/G*CNA����A2�ğ��{حV)�����ڰn�4[�{���NZ��ft+����;q�l�\w3��;���E�C1y�$l\��6��[o�}�V�Zc���ذe+6m�	��"�/���t�����xs$#�f���q�w8�w/�F���B>
r\B6d��0��x�˜�E�`l��5�P�լ5�$ћvט���#��!�!�2�A'��UӦ
9u��(�q��0_TTCm��˰h�"i��h0�io͢CC1i�d�|gO�Fmc�4�e}�T\���7���CqAz�������CAY	I^8t�4֬]�3>D�-�����pSv❶Y$�fW�����y����qB�ܡ�?+�::�~��V�/�:��sB�=[�%	F�T4k��LARl3I�X�#��d+    IDAT~���N�=���t��mST�𔢮�?����2��E{�T� ��E�Ŏ8��鎻���1?S%��$4pw�/����cG�kQ.>��p[�Ъ�h�P�݂P2"����/���.Y�d^r�baf�DYVn^��܁[o�ye����BX]ntx<���!�U,�%���������bwH�M)\9y�����($�T4��fNCs�Yٱn�U��Ւ��V��IA���tHa�)����n1��:w�),V.�7a���b�t�_�O�����N�P����|<�����`4iPVZ�M��#��I�1��=�����K���lt����V�U������t��ȅ)cFuUz���웥�q��yn!��cΤ�l�3y�h�k�T1��h�&tp� ԮS#��\��ԯv-�����²/>��8���yj��Cf񕵎��ҍ�x
A��Ԡ��:��I�c��='so��n�[~y$9|7;w�=p�����\w�l�7�a��-pڬ�^���uسw/�y9��|�B:h F���{�"�����1f�x,[�F]6M��m�$�>=�	���J�-5�C�D,���o�Es{��OcJ �LJ�Έ��M��P��z#.�=�M�WC��àM�sbJ��h�����e�*�>!oE��)��;aS��� Ğ3�Ha��1�/(�'��h�|�$dQ�M_�9�f�4������#�H���C���p��7J��7QZZ&�n4�����'�}��Bt�Zl���V���Ëo-���ygϜAqN�pfR��\2U���'������Jť)�CA[(7�J�J2�'����+��G��aA'��j�J�6��p��g��F"��3sa/�j��ђ��{E�7�����<4��s2O� R���i1����Wއ}������"AknkG(��)���{��S��r�y8{�J� ����O
���G���[LDQ�w ~ڼǣ�=��[~§+W���?á}�g�8@�x�|����ġc����=0��d�u.�g �zMB�N!��lT�7܀��6�ľ�H���Hţ�$(�h�̹6S��O�#�"b��:B��tBV,�Lu����H�5�4��ٰ����V	c�e��˥��#!|��Z�E�S�N`��m��Y�]�va��W� �rŷ�w�u4t���DͅYM�tP>hT��X��Fx�!8c��0z��ػz�]z�c������["פ��j&B�⢚u�FId����RI�w�[A��=��p���S��V��2g�� r?����{��j:���3"������HqRG��&�.{�0m���	��a�X�I��<D�rqgR�F�`6�t0R)�֒{b�vP
�R:=��.����p�wc���8z���P�N���hģ�z�T���˾��P��]�JD���т8';���-B��ٔ\o��3q:ep/J���y�=�cxu�8sr䂧	��r\.�+/A��;�dJI#�4�C^���f!/Gt���q�<Ԝ<�û�#��]��&���_܍R4���򼲄�{*�-_$�vJP�І���c��1��%˛)�)'t���~/��g�7Ԉ�_,VL3t:�G�_s�nx�~��i)�<��T��\�`�!�"䉠��+���KX�чX�a��_� bZ�2,#�$��i�w8rd�$���!���N���L��EYV�����7oām�䢵�I0�"��K��v�"*�B��qd��u&�x���2c�ß��f�I����a#���#͘3��|5"��<�D<��] ����:��V�YOQi1|� Z�[�;�G�rxJ�7�䥘AeIOh�:�5�c��7�=���>��j�)�����z�qL6���tÊ'��XJ-�;�)H�3�ho��w�
U<���V!��5X�cH�v�/NּF�����D���y�|>���R��+���>L�2.w>�b1�᤼_�3��GC�:�Qx��Wq��Qٳ���9+|��5���z}��	[ݝ+��������3((*��iW����DC�]�E�V	a��l�^�|�9w.�}���f���CuK3�>�MZ!t��c�aW��_MԦ��]2ZdvK�Xtѣ��<=�u�4
�s����Kh�V/M$Q+�{�09�p�@Rw��0�rQ_� ���^?�*5�q6@&R���*�w_�>�@$��G������*9�ӯ��ŋ�����\Ķ6����9s��o��ފ�}��av�BMn��v�Z�G��Pѯƍ�`�Ok��܉��'���bǪ5���Q������0X̅�GWPn�UI\9y26~�-��j���M4�Ly#V����N'7�j �y�w�f��Vև�xD�3�-х��&�7z|H�Y���L8�T4�_�|��c��o�[q�~?�vXMF�t��8r��0�{���8�Ft��KrA��L�0^d�z�^xH��6�=+��O?�ݑ�C�bܰ�ؽu+F������]\��F�e���hq�� Jn�~(7���]%�!��^�0��JBsv��d~'�nd,a:�΂>m����*j��v�/x]���o����d"T+���2�b'�+I2�����(	P�0tZ�A����~Vw���?҉��م1�N��(޼2�g셹-�8,�m�\\��xɛMV$Tj���}�1l۵���D~YW�H�(V�߇�S���K�"�ᕎ��Wa_ 9ynx�Y6�$�o�������+���/���K��6�3�<>���V�Y��p�/놌\z����ģ1�FE���[�0a�H\���C2�T$��ӯ���?nX��M#�d(�PP
�++D<j'$���BBP*��$�V#��gr��Ջ��N�%�.���'PZ8�c������w�u;�j��ܙ3H'��R��:�э,(�w�B]c��

$��p,���|"ᄰ�[�Z���q�ͷ�O?�4ى����3
7���\��@��G�(!Q������W��i�RR��'~�vo݆�[B���V��)UZ�]�]O�,����g���NΆD�*{4-I$30Y��`��ҵ�uQ�m��!����=%;��^yU��B�ɾ�,D�MͲw������(��zi���-��]�W���Dm�����j/��W^�-�%��@�'�ӳg^��V���8�)�I�^B��x&��,	����P#���|���5b颏`R'��B�Q䝲�˚�t�EٗR[�5B��H��Y��&;ⱴ�b�3%e�0���Q�~�;d��wx�0��ј7k����#���:��ݢ)�����P#���T"q����h�{�w��hoi���*̾�:T�?��e�t�/�=p�th�	y2@�h�0�h%���]�6� �	y��8l$�:0k�i@ޟ�&T|�� �p0�$N��[�,~n6�l@�N��9$���1u��O ���p)�e�m�|��)N�ii���9�F����x�[��>��#GbӖ��,��Z�����V^H�����Ƽw����a�F@G���3����æq��	���8�Ҥ~�E/��<��&+�g'>!�d�Ă�u�"�wݜ�ذ�[�:z�N�XG~	#b �!K�N٥�W�5���H�Y��?R|n���:�x0NU�&<���봚���1�M7݈=��)��5�4�n� �ٌ����!�2�����u5"o�-(ô�WJ���%K�$}�w`��P[�B��|�Ji�#F��3'�!�a�=�[ڱ��~�s���̴g��!d-V�?�RC9s�P�$� &#�r:�i2ЙHB���Oz��<k��w�cRܱZ�{��%�����%�&������B�EȂ.�xJ���R��� .�!/Js�0$���&����7#�&<&�RH�N���W8�M���	cd�Ǥ�(�bkX����w�pl�sYs+V;B����!��!]�<�S܀r�.�W��5��0Z�Tȏ�B`h�*��dG;?�"���D��d�g�af�9's�E!���,��s&t���F#�m���!�����Ps�7���P<F:�����4ZaW�uٕ�6�]<_�b���G.�\�� ��S*���gΖ\ߥ+�"L�6�E�g��c���F��\�L�,ZL[�Ϡ�u�H(��Ǐ�Б#���;v���t��/%4D%�NJ�::|��o�x�`��(�W�Z�BA������Q�B2yD$���JƐ�pߙFQa.fϸ��_�#�wB�I��%���#���LǧEzGR�3 �.�I��02��x0�$�QAQX�so�����G�{�YY^]���ާCz�i��bA�=��I�O~Ӌ&��h��H�"(]��0�������9�xss��y|�1��ʻ�^{�����c��2R��EO�(�g�/f/�4�p�DB��\��Q���;����x�]w��Im���B�z��`6�nE��}���]x��PZ�x[�]as�`�Z8"*��"���9��è�P,�g��i�N�Ξ���栵�V}�:-�J�,H(��rMr�v�犹�rd��T���Kc*8���'�ce7���"%�T�e�jH�2h �|��������+�Mͭ��}���f�-�ar�	Э[7y�(�̻���Mi�޽q��S��OJ��.*�ч�-M����D�&��H�`Z<ƍf��8N	���m�=kƌ������AP���PZ�w�s���k7cZ�d���k+I�K&�5Ԃ��<g�'7�1��a���V�%sߪ�(��DR�~���a�����'+�7�����f'���C��Z�vD	���2�E�����a_746�z�W���������.V��v�@�v�liv9��5әx��o�����*5�@%<p�=�lç8~p
�N!Fs-V\T$g`"ͦQ9������W+煬9�HJ���	�U�*C��@m�"M#�c�0�YX�v��Jvw�/��O(-)B"F�ŋ��1+!	�y�������!�Wa)J��P_S-�8��&_��g�ѱg?��v�\�F�m��Kڒs0��`����,�"��L�#W�͜���]~z�;�`Y��pU(���\A�#(�Qu�j�J�}=���=��P�O^
x^yٳu�؃)�ј/�r��NV�*艐.)�u'�A��"��HA��C�l�\�����+:�DƐ��2���D��3hFL����Ȝ�$�Y��b��}4Sy�g1k5B��o2��&���698x������@L4�����0��,NlX؝n���8});kE����C���Y��	N9,����%Cq��dbD�~̚>ϝ���[PR�h����%*����"�οO%)���4�h~B��F�h4�¸	S0`�p��P���7*����*9��Y����j��nU��*i�Y	h���%L��q6`�DgBW�.iq��n�y�eÐ�䒐�8�Q�o�(��P,����6P��w=��H\�H{��}�|�rN���V�O�*p�UV	<t����{�гD7���m��i�����^��0�.�8_>�-�w��sWq��aL�/�KA�GP&6elLi�9��l�1�$p�@f34h� X-!�jufi>ɄNƒ/�"���E�&c���<�y`'OgUB�z�Q�#���^�Հ���d������/s�ti��k���/6�
EM'B6
��<�BZ����|r�9|�P�(�V5�:�e��MG�n��x�j�9�e�}��iq�2��>X�'��/�H)�����!7cɒ%�p�]�馛D��B&�Ma�sM��V�Sg�������N?���=F��89|���ֺ���J��ڡ�y�ݩ�776઱�лG%-|W�FN�D@X��Ï�BNB%��ey��bH�5���Gɹ	0AY�x~;=Eh	G��fS��wj��1���?O=���.|K�(��<xu��٭+��ݍ��Yq�A%�=��ό�%��Ͳ(�0��k���Ğ�����=��Y�<�X��:G�>�[B��$�?�f�����@�s�lq�̗���Gi���w2D�].�¸���%����M#� �0wea�����}9�f�6���V�x}��z��1k�L:�����C�#��f��Z��iko�<1��0�фΕ]��TٱB���3J�ր[����!.�̟��R�B�d�QJ�E	ha�Ƶ3�W�y#u�(��i��9����J�.t�&!�G��Os��~�;O�g��/���/�j��ʂ�VS�����Y�y0�������[A���~�΂N�>H��2N�Oa����I����Ce74�b�a���)�<u�N�@B)��(�Q�K���bWj���Bkԋ{��=��0��qd"`�#Im��4)�����Cx��_�b!�$E�n`qv�F����	j�Z+�dX��K�b0JA��B�}�l�]8�/�m��i��j+Lџ�����R�m��(bZ*��p>�5=�U�Ȟ�b/Ĥ)�q��)T՞G<�Q��N6,h�5A"!��s)���-���$��K@�v��쨕��(?�D�jX�u��\�X�8y�J�e��ޑf9�]b>��Th������w��*Q�#h�e?�r��G�K���Ga�i�:���mF�i���U��d�+�󼺂��p0"���YH���҈e3���;�(*ņ/��C� ��"I�"ۘkR^��p��.�7�H��A{H&�/���RLNA�mme/�͐�t��]T�]UJA�Ӕ�Ł�W8D�� /^�ըG6D6�Q�F��x��G���(�g.�5#K���m���Z���uЩi/������r��t�m�59�JEB��Qe��g�z"��`�Ѱ{��a�v$T��6!�)�N�U���)8�V)P�t������d[~f^C�K�B�Y4�ɤR��M��=#�!I��tJ�R����L��^8�D4��&�pehL�I%`�S9W2�ip�I�����k+�B�.� ���z��F�yo2�`6
����4�q�V#��[�S�����#�ɩp���V!�R#��2�q�A��S����6\�'�|�(�J�is"��bϗ;��� �/�:aw6'���gU�N��[�}8v�,v�ދΕ]��$�Q
u�>p���Z�j%E)�1d�4�").��zn�~-V��gN����HD&t��\��kk�k�/�r�jXx�9��=�Mʀ��>N��4�H�V�R2�2�1�Ǎ�R�X_۬V�[���X/��G����7ZZ|�B.�q��P�ȟ�H�@�ن�N�p��+�oB���2�%���(�i����M4�莑��tF�5	��H��/I6��VA)Ā�L�Z�Bk2�S夎�i��{�{��=t�߹�n�����5��w&�����Ν��9?���Ǆ8�	�Nqʄ~B �|A�C�fڴ��/s�B�/�KTLٿ�R�)��"s���K�~��p�d��>�r,&[Q��X�믽=;wDCm-�
�n$�1��R!X�6ѻ.�x�0�y�Ϳm��L*"˖9Il<�	��~r�g��r�
a��/�/2Y�|y�lv� +��Nt:e?���b��o�8��ۈt4�l<����b�)|�{'�6�R�6��(N�ҕ����C0��
+��2�Q%�K�/��Y�s5u�g�3�L�S�f�p~�rҎ�������`K{��F!�����Rى�^���[���#HFB�r�$i���>�Q��k�19�����u7�T؟�ρ����h�aD4VB:2)�}�AH��p���y��7Ҟ�D�hiS���X��Bԝ:#;Sj���4���U
������Q�#�w�-�S�	�#ӊ)�[M=�d�'�j�u�]�x0)R�(�(?�-�ҹ�6��m,DgϞ��/��Æ�}b�y$d�s�%��S"Mf�eq�#Z\ʢ4j��n����(�L6.�$�p:,Hƣx஻��X��b �B(Y�M�>���j�r�������f�tT�I>�4�6��`�,>w�Ҷ8?u���s'�Q��������_BZm�����2�)M�F4�,���C���]�}�J�dr� �y�w"!�]�`*�$�,�fY&���Np�Hɔ����f�S
�%9X�Y͂�A	�\�l�S
���a}՘���    IDAT�PZ�u�>��l��Đ�Л��犀
����Wȼy�b��$���d<�^	$aZWeh�f�ͩ� ��.�5�4>*��ء�(--F��/��qm��*@{k�\�dZA,��-#zӒb'�I�ۻ�ZLV�H/��Eȍ"Nƕ<pj�5���f�ː@�1�{�T'�r��l0�4IeA������������ J@����7/���ܕ�T�H`B�R��4�C2	������f�\H�b��R�Y⪀�-�W~QsN�M�[lɋbs�a���y�_cY�zlv�)�p�,�wl�:c������%(�5��3��8��:�ЦT���c�B�� ˹�.�C��s|'��������!�NC�g�C��5a�?����Ѧ��W�\���Hꎄڠ��+脙x��:�?�.�N�\��̲��$s�;�/�l�	��abVC��\N6��h�I �FVg������1���ĮDn��"�g<a��έ>[��tF����Č��)v�]����F�T��y��1�>}�L��Ӎ�?\$>��,]���ehjm� �_px�s2ƐE�樳hJ]����d6J�f"�ì�SQu�(���3�BL"�QQ�k>`<0x��|��H&o˃��
\�BBlX�;u�s5�b��BdsX�|%�	!K"S��7?�0>۴�tj���p�Z��إ��(V�Z���F�Lt�삉&H��I
�_2N^ �=zbȰ�ٳ��\M���ȮO|�٤)ŐS���Hjr�y��e��	��s5	�z�^/zt���ޅw�zg��0���^HL54����:9y$�D�
EA�)[�-�(��8�Q�ŵ�5�3�;��Xp�|L�:�_D8�G��P�5�$%y<�رk;֭[�4��|�IT�w@Kk�V&��e�g�7Xĩn�K�f�Z��"Ƣ�����|Q�`�����d3"	�a�����F��x�I��C�{��B�t�U�&+�^^Z��hyՉ�*�O�_���MQ2}��P�VU�G�ŒHd���UВ��ŕ�^<�M���E��y�3�/"aܟ�ܹ���p��"O�4i�|���-E2Ō`���p��1��6�C1��cA�LQ����$���<��N5�1u�T�0��ECl[�"]�v�dq���w��f2�����H~��"] d^��܏��b�� i�����Sg�6Ẑ�iVԵ���=C�NKk���7��Tt�-�3�f�\�� �����{%i��r�9�r�����-Z1Zٻ�d��.�^g6�,�r��ڂ��Ƹ���L� ��4T����Ŷ-�p��1��*�"Qٱ��� U���y"��t�:��[�p@��Ndè7Ʉ���� ĝ���$�*�6�p!x��|�k`�¢7
r�ՇsFGn���R�l��U���G�!t���eeB�Kѧ�ꀹ� M��u{�z	0�V�r��_=��DYÀ�D*�VxF�m7�k�}9������
�YgFZE�9^�('t_���?�8a�w/���7�����?6GS�#��w�WYЕ(L>���td��ѱ�	}2
���/7�,�b_zEAgg�7�ZE 	�u�<�9Y���Łfo�xR���%`��_�X:*y[q����m�F�9��k���]�ƈ�c��;oq��2�+�ԩS1f�Xl߾S&�	�'A��੟�,�Nk��/�&�M�� yxHn,+/������:)�|@�,$ƀ~�QP�`Tk�cڄq8u� Ξ8��R��t͢(ȑӺNR�U��Z�����1��b'Š7Y��7�x6��,k�`:�J :v�$i�2��6/����I�Ɏ���Z>���W_���H,�N��ݺc�a�sǫ7b����-Y���T�����˖cۮ](,)C	~0+�vꅹ���I��)@��8''"?F���Չ�L��@ ݺt���7�D�ٳR�Ut�S��:G�[sP�f���c�:A��B'w|�t��AA�X��Nq��4*�Y��f��ɨ��p?|�f��d-Ə���"|��KD#\u�X\�T/���>�{�ZZЩ��((�v���B� ��K�8}�<��~9tｳ�����`�T���� #Gl0�T����<��?U"#�<`�����8 ��5`�����WC�(?mC�$�1,	���z����E���V��[���=���8�4#TE@�K����O�z�֯�6��]�nspl�Y7l� ���fA���F�����<��Ν���cas��O���I!vҜâ'7 �h�H��4��j�4n�e���AdC�%��n�1Cd����gd1�0��A
�a6���-S��*��<��w���i�4�Qi`w9E2�H�@a�Y��V���3.t�p�-s1x@?񌯾x��jT��\����ߒe�p��q.�u?�|A׈pR"IN Y�<�������}��7����DD")q�w�6�Tΰl⨐�H���Z��,⑄�9��|����p����dV��#rX�h�h������D��|����l��(�%���'����˦�`� ���"��ɻ�g�������(N�>#�O�ݻuE��4$d�����ę�p��-��V/<e�Ҥr'���\yxO���*$��c���8�J��(��ot1IeA'\�_&t�����^�o6���\h)��{+�k�en�A��o;�J!�\Y�I���NE.)��+��l�y�DYL4b��}kr'|,��ܮ�Za�x����Q�������a��r�:�<f����Xd1�2�&q{�:q��^=��Hӯ�CF��SO��ƍ"צ����C���~�#|�a�X�q�w����f�X�V���g�w�_�ԩW��j�'�V�����8t���}�Ķ�1r��;p�j��G�)�B��p�U�q��~T�<,�aL��R�)�,aX���e��!�If吐���D�D:��}�7��YamO���_حF�Q:�x���������]�v�%;�|u�6_ܻ�~�i�^&c]c��A��?���D�m*�./�|��窱��{��k�@}s�����%���'�J����SQJg�`H����셫���B��:'��H(�
3�&�(*��$�c��o���9�"gF�f�����+DR�o��C�����	9�r�+F)�|�Z�B�Ӱ:���-3�R�)uF$�A����}	���Ǿ�(
]n9�kΟ�kAm�[/+��Я_?ABV�X�z�<� �����w�ǃ<��Kx���a�Q�L�
�	���.Z}^t�; 1��H)��r���"
]D}AD�ðHE"�e�LmX��#�p�	Q+�׃ӝL�9~���r�3���_�b/�/�	�%���j���՚DZĉ��2�Ns�]{���'~�(��.��G�5jq͔)��>q�8��E�ǵw�]�
[����cGлo���;����7�v7~�g�Q6�Z2��V���).;2�5�p�:�IM�yZrr��F����W��.˱dѻ���9�@��.ş�,|�i����'EO�WB�4D��b,�
�âNR�9LF;.Ե#�QKЎ٩��h�\������vmیS'�a�����ը�T+�R<I~۱k�Ğ����6c�u�9A�xBP/z�3X��R<�~�ܟ�i�v��h�ښ`s���ʜ��A� GZ��*,w�����K��l�":�]ʋ%�(�mCQA�V����M�D��~����ZY�i�y��s&�g�X��Y����Z��"�m�͘u#M����s�
�����qXm�� B�,�PB��ǏÔ��!���T�h`s�%f7�գ��k6n����B4 .��J���Zd8aE[k�~y�q��=:��<�0���I<��m���Nȝzrw���^<�3l�?�|W�ު��7>\�Bs$9;�3k|�LM�Si�@��P�	]E蒓Y��8: ��s��xXX�$}q���{M(���7��B΃����M*;��$�;/(;�
�
שw_L�~�LX��AHk�e,$����h�p-u�q��qĢ��5v^�t��nW�������wP�^��DFjcs3N�9�����lt�v�ڋp$*0��cGq��a��47g�<lݺ��w�w����z}�p�R�KEba��(�(J��)L3��ޅ��g`1jD���vΙ��H�A�b��J+�;JXNj��i 0
�ބ���;~
�f�]������1��JQ��`H|��菹�fbӺ5�XV����|�����c"����Ĵi�0p�`�?t��t��)��ɓ'l���Q�8{Vصo���--���G�r����'^{�U̽qƏ����ט;�f�u���������"���BsU���ƂΟ=K����*�(��5�ń$�&%���"�̄ͅQ
ʚ��E�_U�l�\�.={K�:t�4T+��� Ij����g.�V|�1zv�_k+��,+..�_���Ȇ��u���ի*;uD�^o����c������
w�}/.5�w��fL��fΔ0��;�܍��Gb�GK�o�p���ڍ��d�1�(�x��t�ѐ3�'$��7�F�ۈ͛�J�+s���9F���s�q>w�_�O��X!�ѳ�� z���I�I���-6!Tq2�ޜ����N����7��f\3ER��h��m�#=$�W_���;�yUZ�43���3OK��9W��cFˁ����(*�C��~�G���Й�BX#9ҨS���Y݅(���,P�ښ��TAO(Zij�s�O'"�:y"�Z��H��!o�x1�/<��j%a�ɒ��0Bsr?��ͱ����Ki��R*�V�����$���Bͦ�<�v�{�Ox��?���	����8s��՜CsC&��/��%g��8a���W�I���[�ϝ<}N����~���7q�L�pX��� 
�S\���t�p�%a������l��1슈��:���`��)��n�r�;u\�p��`���@	�p-��ym8q*�02�E��K�6�p2��{�}L����HHrŨb�j�v��4b��סw��x��1�Oo�����G��E���p��I��iEd�MW0<�t�Ut��k���/�F�a#P\�KW�Ak��pXjDSc�DiG#䂘�7Y%'�"�p�:�WX�94+נ��{�%㲇#*e�\yȳC-���AMt��Fb��{��_�yԘ׿sA?P]���E�^l�gf���]:�o����W��t�!��5�G�B4���.�NUI�Q�����cp��X�)�K��	ه�|�.Xѡsǣ1��'q�ÏI�vCs��7��+P~�n&����F��X��/]DKS���c8t�_��@��r;��\�h�LPS�N��@�}Ί����KrC١�Y��%eR�X<�w���P���[�r�'2l�����w �'^-V�l�nU"I�C��ޓǌ���w���s�0T���(9ْ̗�4�ˡ<,�w�V������:Ƀ���A{�̛D��ޢw��Y⩢�A��ʡKw��#�c��-�׫�ߋ�Ǐ�;��= ګ���Q��,ڷ� ��mڰ7�x��V,G�N]d�%t^Us�����5�P�Ԋy���� ��,B,���sS'O��~��˯�wy��]�G,;-[=��bdԓ��A���zu���`��o	�Nltje�]��\Ag�/����G��d�J2��#��m4���a�lޱ��Za�;�~џ�k���9o|͗P{��H��1�-�F�n���ॗ^i��G�����������@C[*�T�бc�� �꛰nͧx�������zL�v*v�څ	S&�K�م��a��;`���%.��n��W6����^�̝	K��ܓ� �<v�����6g��sk$��_b����t�(��E��BX�1�΢bi��}Y��� Ə��C����o�n�$�P_'��O>%�>��3�������Ç�{���f�;v�@s��*�����x���Ψau{p��<t�0�4h��(V�ۿ܃�3�ûK�5��ff�����y���Ƀ9؆y7̈́�f���¤�"���i5 	�*v���8�or�n�y5������9����hA AE�QN��O2:T+W{�?��֭E$�Ť��q��9�"!)�?z�q����F]c��Fc��H.)g㯏=�=!�N�4�k����D�?���_��M^a�-7�=Z�vLfr�xo�x���p��G�W��pɻ�3-�AW$��k�"�����ضe#Ο9~YmB���b�|��TЕ�L)��<����.�2���j��`��:B��Z/�8�_9���̝y������c�`̨a��xm-Mr��F=>��#)�T����l&,g�w܎�����V�=���ko�Wq	�3p��?/�keE�Hn�$�����O�Ҩ�()�B�ȰF�pn-���B�LB�X9cr�����*�z��rAϑ��=�\/�0����v+i��;��S���ﮮ�pњ��#��:��:�K��Q��L*a&r�/�K����	�KI���傮# $�6���}E�H"��+�9g�LB��eT+��q��9��O<�ӟa��m8|�ϸo%˘0X<���ߋh��=�w�4��
֟��)x}����� @��)�D$�x�	t�����ѱsd�*��6��p����Oᓵ�1�$OX�����^:�w�-D;�ld�����~�x�8�9�J��S��4�$t���%�bu�z&��eL�N�U�*��Uc���U �*��ku��Tbʩ��G����!#F�g��X����b$'�%���.����a��U()p�ı�8y�0,��u���
��Xˎ;�����"8��[���O^���=�()+�Ac�=��G�֠��"�y�A�a|�u�X4��w��ұ'����Y�����������Nx��av���7K�a�n�7c��tN��XP&t�ɀ��U&#�6���$�J���c1��Ϯp(8Yj�h�%/��w�u����Eɕ�Vy�}p��Z�m�}�2�t�R�ǿ����T�@�ջ�����C���y≧���Q{��P�	�O��T.�anٴ�ĬY��N��`�<��}��ޯ0������y,Y�
��!U�U��V��&��<��$��$�s��c��DQ�[$�=�+�bZ��a��C�xy�rS��	=X&h�f4�y1e���X�X��&���ŸH�5x�'#�<~,:w,ŗ۶��eG���6�`�'�	���[R�X���g޵k�\�Y7�(�U����}��eŕ�����G+᧮�jø��ѯG,��]�4cF���l��Sg��_Dqǎh��V�a��X�p@&r�F-ҾI�GK��ʥ���Ҙ*�6��RԘ���I&�9�B�9�j9�s�(�N^��r���p��HC�X�cT��-�f�(u�p�m�aŒ��ǈ�`�+1�}����׏~�8T�,Ǝ���Z[ŕ��0�O�<)�����r���3�s�|�޳{���a�§Z&�7b�ܹ8p䨼�{���DG� ��쨃�b��#���a��sf��k��8r�!� z��\w}{BW�;��O�t���l/�Fh�6�COs����,�?�#���(.t��J�NC�;5��ڵ��Ͱ�殝I�[�|��c����
����	'�*���[�:v�q�'��}w!ƍ��#GIC�ɊU��k j�#4��X����RR��	�I���(h�¯�s�}"����X�9�;i�R��7��?�=�j���t�_Zb��SZ��ۤ�otE��ܴ+!wN�,�H@������yLq��C�|�Ť�(e��7(a�����KЉ�`�C��#�TXl���G�sח8|�$lN�**!1$:�������ւ�֋��o������ΨÖ-����RN����@�8s&���W^{�:����޻~��?��g������HA�8q"�-��ZyiF�+�"��?Q���:!�e��FJoV$"�4�4��aA߅ڪS���Ć��D��s�b����5�ϐ���Yйs$�^g0#�j�p�w���Ͽ�<%h�U��    IDAT`���a��O����!���oP�a԰�رs��~�gϒC����Ңw��a�����޴�3aj�3���칷����{4���O������a�+y	�̻ӧMûo-č4s���E%D�X�f�HF��},�Υ̟9�>|g�)�;tq��N<�3 -��\��CV����b�7-m��NRY"z<�ď�|�Z|�s7
i�HB Zy�J~����u�&4�7�CI1.�;/r��.21���K��RE����6~���8|��(���BC�V_�53�Ñc�$��'~$��k׮ƵӦ����߿/^|�ϸ����ȹ��o�jw�C�
�+Gh���Ю�.c&�7�B{]v��D6�NP�$����,-��ݓ�ϙ�\&����mZJ�p2�kn��x�e�ۜ0�\�I��~¸Qܯ>ߴ�.N?�T$&L�_�����QVV�s����&��믿Ɯ9s0z�HT����C����W^��#�**ǻ+�����
n�YU�C^���b�U��\�ޯ?~���%�J�dJ��*C�Ai���g�0�i(q۱a�
dRQ��A�3�˵I�Is�H���+'�+�,��T~%�*�,u��������ڜb~ԥ��q'���4^��V)�l����}������t��߀�غe����q)<6lBqQ���j�p�̹�l�Vlݾ7͙��]+�Le��~�8�KT{��J:��%˰��q8<%��h��ltz�,����a���ǆOW���q�x���m(t{��U
:�xBΊ�K��R�u���r�	�L#׆�'Z�Y�UL_�r���-���qӌPg��r�碃g2�%%�BV�@��s��A�0t�0�<v\�	'v6�7�4K�Պ`4�O7n��n�U�{.B���F\�d�Hۚ�[��1�W4��Bc����-DT�A��D�MR̶��]�1�q�(gz��{A�ϝs�9\r��i��~�,�|Ӹ�^UY���&��gj+.^�zk,;5��#U�d.��)�U���)./[�NF�J w���	).B�%�+-�8�1P�qń΂�	=_йCWأ�4(Lo��	{�Ek.(��ٷ`Ǘ_���N`Q�)B��I*�{�Z���F�Z�1fL�&.%W��en�\!:P:UW� �W��-�j����M2���ޣO_|�~�?�����X�I��Z�T"%S>�Ԧ�����hH���z
\� J"T�DC{�TB
��o�¥�S�Jv�Z�)I�}�s�Gqz�MŮQq$�n��C=�|~htf�]%"�>n<���%˗*A`����FBP�n]���o~�s�5cG���U˱���PVV"IX���yńAGX��@���� :�)j舑�;oV�Y��Kux�W���;Ե�J�B����C������܀�C�ʋ����8p��p���9�-�Bv�ZI�U\�h�ؽsn�>k�.B��Ӱ1��o:��N#��Y90�Y�5���%I��
�G�=^����ъ��9�⓵�}�W��܊�5w;�b����⛯va���?v��>�TW�v��k�I�R�<��`6]++1t�0l��s�.̽�61ܡ��3?�%���ॿ��AÆc	�����+,~���W��>��<�O�nG$�ЗRy����dL�2���0���u.|��{�dc)�dP�X$���|A���.g@"��Ӧ��FJ Ы���XV���[��� �˥x�gSh�P�y��������O�@ߞ=$�#N�$v6i���]�r�mm�Ҝ���?äcǎcҤ��ѣ'�y�i�4s:v뎧~��ħ��ڋ��_�@3���̻�z��r����i�q����)FcK@�#�*�Q�q��W_B���4Q���7���P���v�P�x,,)��ٓ���Z��k��rn�Z���1e����s�`�����~v�@D,dm�{Qdq��?��6"#���1��e%%���?�c�<�M�eE2q�0�&1�a��O~�SlٲE2�uF�8�Y�n�4�nڂ���92�Mҝ`���v9dűt�ǘ��X�~6~���O�&�OY������dN�zU3�����6���YX��Hd��@%��]١+��l�9���&��{�
h�C�9��$H�V
����X�T�&MBY��?��+ʠ;u=�qո1��_{�58HP�����ݸq��v�}��Л�D2��T�}�#��H�ҊO>A�N]q���8�VO����k�[@'QWi)����h��йg/x�QX.�	��s�J�<��[�{���w�/��C�t�.�U��ˬ��_��}��]��x�mIL�A� %$���S\��K8!&vaB�WHq�p �;KA�p�t-�r]���(&j11�<��!w���e���b��	��qd-*��������hhj��j��S/	n�wοgO��;o�!�(�v�t��uu��n4�!v��yd(3���D,^뛛�����8Yu��n��D�Z�����T/����sh���o���tB���
�bP ���1L3G��A}�Y��q+��/9L�ѵ��a�la�>]�7dA'�%M �H���+�����
=���K	�O��"�V�ڀh���}q�u��󧟂ը�pMm5@�GJY�
J��m~&N<�� ��s�{D��&5M�m((��O~�����`h�`0�QSS�`��Z����T��HD�\�$.f�~/�M��L�NeŘ�t��h	.�<)r6���+Z��� A�Z	z�嫳�-k�ɔ��~�t����w�ͷ߅u7K����F��Ɗ2o�]nE�عuF*Ń�K����WZ�#����b�¤7H�4�?�)Y�ojF�Ε=f,V�~�����,_�Z�I���@�Qo .�}��������U4\�G��DY(�.�b�0T���f���}�Zd"!x��E��+��bU�+�����W����	r����Q�v�웑P���w?��;G�N���+��4�L��IcF᏿�f^w������+1��ޜ�&|��Rk��7�����M%�j�,�o���
��0�Z<��/a+*ǜ[�{["�Ǧ���0�1w�l� �������N���Э_�#!�|>!�:m�kT�2~4
�6�Z�v�^ȵt���g4g0 R5ҹ�l��,��"/�w.���.ޛ#Fbǁ8����)�*m��*����g��ﾃ���Q٥B
�?�&L�[�݌��Vcߞ]p���:�ns����7ߢ���p�=hk���ƽ~�\������fb�5�\�n�j̜1�M�.�ˎ����V,�d-V�6L6�X�Fi��bM�f0�V�3�`���|�I�j$�R��v�B����+�t
��ʂ� ����F�n�jI�Qh�iL�/Z�gRbk<�O��б��I���&�gϞX�~=��:�W��͋�ΝQu����:�~�]ر{7���8r�*{�@i�r���/�SP�^=zcذ(�"�W��[eػzڵx�o����$����e�'����� ��'1c�w�.��
R:���ݪMz���zӸ������U���h�[�I��hV+]��ik�O�s��)��҉Kn-B1��Y�{u*�*�	=Ń��:H*�"j�+�����.�$0B-L�I*,Q�3'+Zv����a..��waݧd�iwJ���L2��}:�����%)Z�,��J�%��С#X�z��=�&^5�*�Hw�N'8jV����-�j�|�s�tl�`D��T4	_����n1K�֜g�ENk1&���r�UPz��#����{PW}N�Щ ș���0� )
<sEAg�ć��;'`r��\Eh�1n�u(���+`�9��@�,f$�`X���͞��W���
���_e�Z[��nlly ���x�2��P3�/�%�(t�V�����xG$:�
�X��P�tX���4�Z�FC���f1
a�!��E�D�d�n�q�ঙX��c)���L\
:W:,�|��A�+Ӏ��؀�m5�ܟ+�bի��k��w���b��O%���É�4YŔu��������Sx��7D�,rK�t��(��D]�%���S�8�E��5��uZ��y�|����D}k;}��: T�eFJ�|A�;y���@$Eܪ��Ѕ@�ꡧC��!� "�J%KFZ���y�4�5�HA/'�>G8R��s�e�9SR��we�'ZD3NQԟϚ7Y�,[�����(/U�)\63���~ݻ��?��zt��ۂx"��v"�j�9R�P����C��Ƒ$Lv��#G�b�%�:#����<�Gh�n!�1�7hG[S,F��N]�A�5���fq����l��0:��ۣZ�ꐎ��kmӧ���`�k�Q����.t9e���7��JAϧE�hI9�K^K)`9W=��$�C�.�KCc1#)�E�^N�?y�1,y��3q�?}��h F�CBmM���6���Pޱj�FVEE%8q�XdO�>�D'�T�?�%�|{!6o݅n}z�d7bϾ�����"B�e咖Hfw ��#�D/�,.��e�/@,������0c�d�[���j�ioH�R��T��!�a9dLX߹�Q����M�4zA�x_9�'�z�U4���CgGڛp�-��W�.���~�a��Cy	�'g��������UP;��D\���Ge��6����O�7�Diy̸�z<���(((ļy���](��޽��Pe1h�(pz#x�����r���`u��N�4
J�r<(��g���CCA�Hq����C�z6z�2�+����]��������_�x�۾���(�֕+�m^�b���E�'ɲ")N��N�N���%�P�C�=qɰ�l�����`F90X���#���:�����a ;֋-m��t��<�%˖����0I"d�ӡ��p���P�Pf��A⾎A!�[,K�e���&'��]a���g���;.:3y~������j)0�����L����4���=N���a� DJ^/]����F��Ҳ�0%��)c������p������F
�@9l��T �!��G��T�|6	q��P�(�z:�9���a�5�EW�e�
��YJ��f��f�𼹳D����A*�m'��6$n\�I���4z��3f��!k,Q��B��7[���;gF7yL���Qj1��ڤzt��i���6J�B�O����l1�Q`�"�a?�w�YӦ`Êe�!o�3.��N1��b,��K�Կ
�Iyn��0��$}1<�7G b?�..��{�[���Rk;4&��[r!b��G�=�vűC��'�^�Z�i�6���;";a��M`d��y��&�@�٤
5/�[Ͼ�=pv|�5�رS����6;|�m���:�Dk]�3ܕ��qG��#�)���^�@y������u�-�6�cê��Х�\���3��&��|aOq�bb��˄��
f��U�7��Ye�X�r-�%H����+|Y��[fވ7_{�U���j3 ������I,�gX1P�qⳤ�	*G�U�����Y0}�l5�/[���8F&S	h9E�B�y��R�4��:JB],��bñS'Ӥ$ӡ��m���
���D�Ũ��+W��L��&���Tii:�[�d��4 T>�'9�OP��Ͱ��?>��dJ���;h��4&I���Z�f#}�>���������Ѥz���,�IqA����l�[�ő��/5����7*�fj-<�%�.��6��?�w?@0��7B ��m�����)�.�K~܅���M���چ��"	���OwB摗`��)X�v��ka֩��HX	}|��l�*�;���q�i��>�5,k�:��M6�|��4�"O*MdO���zL�8������W��#
W��X&�I�^�sg�亘f��qO�j��F9/y��y�ر�KTt�1���/�;2*
��҄+�x8)�_�ˌ����oll��o ��V/�"Tt��#W�4:��=:SJ���3���d��ј5Lg����OT
z�R��挟��w.������'k�ecC	��F0�F�)k�(V���{�0A ��4�HEѽ��g�@"��êG<D��ՁX��#����S)�| ��L%L�-*�9�ɔhT/56�b��^T��~#0l�$,[��>t�@C!�0=�B&��zW���,����b����b៭��{��t
:#��H��zR��D�4�BY  �w:oE#(+,FkK�L2!t���Ƽ��3��@�OBCĮ�h��aC�ȁ��X}%n��hN ,�T��Ie�U���K�#3��B�z'lC��H<�X6�� �� ��86O16n�B@�\!Pi ���p�N�FBAWi��D?K�����R��	%�6hIX��%`f�C#�&1��"Qz�G�1،Zh��(��7���5��/-)Gqi�h�i�ASk��y<%EBhj�ѵ['\7uV-� ��F�I�;��B�u��d�c�H�6A4��9�r��4z8�nD�	Ixjl����{�X��rD�Y�p�M�A�4Z2D�+��F/h"@��J{�1N�9���A�x��VY)�a�Z�J�(��/^Į������n�ܛ��+B�I<���m�݀��"�pp��mj>Ks}<.�+:���I\�n�e.ڛ.b���
��G�
)�|�hJt94WL���z۔�rf�s%a�*��|��F��Yi����A�`���ka��-��b���]���{�E�)�>�H�F��(�f�4l������r�~�7\�~�:�*(Yh�C�8}�o|�A*6z�ل}(d�P8�@�W�o�д��a|r\l�[��R�63lFq2�'���n�fz�%(v9�XS�Z�Y%�n�ɘ�&�k�G(�`#����{�9�310��"ItZ���F]{�XV,D��Ks��W�J<����j��=u�xD,s�3MS_o馆fi�� fF\)�kf�܉�0aĘq����q��
�	)��Ρ�iE<�C�(�$b�as�$�ͨ������sv���K�0��bw܅w�y���f�A"���)+?�V+y|�t򣿿^+��4sb����gi-�2��*DFg���B8�AJmDF��ˬ����'��������1FB4�2O+��N�����J��hf�*�r^�Iq��*I�����gc���X��3\��`��a��M�j��3��� W�K�5���ɄK�u�S_S[+�eDN4D�#9�������R��(���>Կ
:>��ThM\Q�`ӥ����O}ˡs=�[���PV?:W����t�QNg	ŧs�;�WgSRЩ��P�B4Њ��М$ ���������F���U��"�Z.6���ʋ�d�e��R�t�ܳ?�M��M^l޾M:!_&�Y�zXxٝ���1F��I��x-G�p9\��Lbeh�
�`',����E9xN���Z&-e֦F[�J����!E��xB e~��Upzܰ�,�AB��K5��G�vy�S�J����o^_CH�~��}�? ��	U�z��a��CM�Y�](3�M3&K	c\64y��?d�e8t��CX�j��E2*)�DLd��&Z�.YYu����/�E)�B<�@VK�0��2�Zz�)�l�8���
3�]��"�r��.�/�0�B�g2H$���HgThii�{֧wO�"A�#!�77�dGLS��h����O�;����Tz������A�g����S|�r�:�\�VV"�Z�PVR�@(��� ��i���/o�2-�$f�3��F��A�h����$������{�$�	�$�1I���i�}��� ��i0���IP���D�a+6�=}Z`ߒ�2)�t#�f͙3�&I�Ub�b�90��9�7b˧+�6f�I�e��p�"��y'3��fJ=��(`�xCs�<$-rb֨4�����0�U��Ps��t�Z�β����� ٺzA�:w�����"��(�>���ʄ���5�I��H�+�&H��Nij���#C�x�ANT�Ǚ��<nA�x��y��(�Z�
�E��<����"��Af�`q�:D@�N    IDATњ�7ͼzu�,]*��H{�D0�H�%v��+�3����Wa����R�����D+R*�X�j�.�85M��i) ���M��1`�Q�קR�`��ƀ]��f�Fm�=��Ϸ�̙��q2�M.��D��&�qyf%�M�p��h�JA�F�l��Q�j湅x�����%%� �N+����8�x��LD�קD�>�����-��$���hN���)Qr�ѐ
*�7��T�$㊽+'VI )@ֿH�=TJ��b3�v��N7�Uz'��fӖ�
�mذ!8s�"W�F�5�x�C�z9��۷O�w�`ф���(��eC B�C�A�a+.Ż�W��� c��Z1k2��H�²�av	�maYL<��Q�%-mJv=����R�LF��1��M�Wi���4ʢ��_��"�V
:��(�w��o������<�q�Tυ+6-�8*�傮X���]�o]����SS��Gm�U�BK�4Ԝ�^�D<�'^@�ޱ�K!a|�kW�`�p��PC�I��\����&�U�hJ��ƆP��dw"���ki�F��7�V�i�P!_%����(L�&�&�!H��;|���`b����=yV��9�7�6�f֣Ki)��틸��Rb�AG��GKt�]5b�d��=�����S(�#NçO�:D��*�L�˪u�Bk���a�(�j$pCR��s?Ǉ����n�����F�!#P^�&{1�}8t�4�*��K��M�s���Ծ�縙bŘ�8�%�2K����}/�b:B�Z#�� w�S���2�nV$�Yes�rCD����,�ڠSkj�O�����d�PP����W&d�������qv�W��u��w\㮄8A4�H)PZ�V��Է�mw[�P�^(P�H 	b�]'>�3����s~7��y��}7��'M73���9�9�`TK��f�~�o8u�0&�4 �߇x",.R��i��F�(�<���{.�U̩�(�HoE��D~R���GEEC3~��k���3<����Z��r�J"�J}�pC���gx-����u�F�����J,��W���� ��b^���~�z���a|K���PH|���Cr��GP뫐���𰬾������c_{�x �n�'~�;/>Օ�6Æ��(	���H��T�t��6&{eI 4!A���CE�y�878�w�o{NoM#"1N��/�6��2T�8keu%I��tN�B&&�����0�7y�h��~`*��w��32E�4�u��]� �!�Q�5`,n�~�
�mf��kD!N�d��p[�p��P_S�7^~u�^�wv�ɔB�$��JɩҨ5!�+}�pӍP�L�y��̵WCoq
\̂�4iN�M���M���'�����`���D�0��F�-Q�Pr�$���#�~�b��b@�'y"�\�rhJ�2H1��(+Û�,|��Qb�!}E�i�w ��˳��DƦV鐎'�hZM9�J٤L�=�1n9�$�,��0;Ki�(q�Q6TF�D��4'��}�il��r��W2H�ek�E�)�A�k\Gѳ���t`�;��\�M��I�b�����ݻw��7a���EF.u�����[����Ƒ3�q��9-FBKC�/�c��@�l��!��m1��K�0<2(�	�)���V�K$x<o9��)� u�]Y_�-(G�}^�u&-J�8,�~��%/�n�(�����l:qn��_�״�4�"�~�	˂Β�	��I�����D�)�{jB���
�p��Hgr�0�+��"I�R��Ov�݊@0,/��D9�J^X~��')�iD�GP�,���޳�����"�����S�'L�m~MFqTc�ȇ�LX
�A#P���|	�����à�*���>!!�&	O�8����҅x8�g��~��pT�Ƹ�K��օ��#8 �������O0y�x��9�����%C?������g��8��p��b(ݛi"�Vԩ�e���F[\�r���AXY��SI�=�؈,���U�8}��}Л��̎Q�mxu�rzT��H�i9Җ{0y��#���4a1��p��g��#��?W	)�K"X$�
$��P�����wݼ&�)�kMd糴�������-��Es���@$��`d/����K�P[U�|&�Հ�Sg�~��k*��tQ�'�B2+"��H�Zy���IFE=�dq��t{��څ�<O�lW7,�D�J:�Yг��A���-��>q���H��
GY](F���� O2aw�GA%aaqF.���Ǣ�ʋ��0LZ�*�q��q�:#�����^s��D�~��(z�>�>���!P��Kf���ض�}�P�t ���{��t z n`*�'�WX�dѓ����O����F�,��n�3�u��Vj��_�੗�����4�PD��^rr4�Q��PȦG�SA�4���@f"6�q2����M��%w��d!c>�N�4Z���/( ����d1aP+�+�N�w��)6��]���G��v�t�a��mpXL����t�"dԳ�/�f�Is$���)azWjL�c�bI+A1FWZ��FW8��H�b�C	�x�3��4��<�_^"B\;��Z��_NH �T¸�G��Q�E��";&Q�͢��6��l"�Q��A��,xz������.k<��,F�����hC�D�M�R�ظ�����#�A]@�?(�S��g�=��������!-��iN�by*�	C9S O�,#�F�f4
'R��ufi t���)	�h�s0A$h��<˴vV��6<�N}�t��J͘g6\�^���Am���%�Ƭ�3ס�B_Fd�B���G�%��ߩS'�s��f
E$7�duY���tV�rO���j6�
W��bJ��,��MA_w�u�+�{5���N��ݣ"m��:z����fW%�Ir4�)f��������%S&bɢK��F�����2�F�%�%�����=X���k�Lx��W�~�'Xp��2w8��F\��:L'Lz�iʔ8��M�eҤY�iI���?e7$��ߗS=��}F$^�:��I�lF$�73���k��G1��_�e�5�"�N�9>�`֯]'��J��~�\{��n�@,�o�����Ne1f�d��=y�0�B.�,������b<�g�~>zH�㉘����5%�N�,�O�g�����[�%�ؿ�J�$Z���J$sj2�H-=C'G�,6�I�i��
�<ti�[&uC%B����l>$Y�({�"���ɾ�)i�Xu5�H��#�{�]���%�:�/��zB�E�O�Z�C:BC������q��U���i����Ahx ��a��@6��jT�p���u9h6����4�d�y�Դ���a�(THf�oD�/�َ�� ��)S���]7�}
E����{\ٶR"=i�Akbj��z/'�q#�T��H�c#Zv�cP�Ѡ���a�/~�C�z�8w��^/�����O6#�J��o�y
�����&ڌ}��`՚u�3pV��A���'E*8�Ho��n��4�B�?�s~&�x 3N��\.���v�����0�atzਪE^g�^Bb��Qs,�:�J64S�K�X�oq1'�` ����pe�d�"���"�H�=2�s�(p�B©�,�bw{͙���&ìR����ttv�=t$��93gHDꩣ'!����1�D�jj�0��V�	mgOc��K,_�̣�S��� J!�ʈ��4%l��YF�2s��q0��tA�4�x+�0i��%��nҠ�6%F0+	h�e�y��0R~'��4>b��xN�!&&R[���'S6�b�R���d\)^Z@�K����DV��r^=�á�N�9'�HCm�B��J�cz;���)SkUm#��j)�kk�޺q-��
)1��˳F�j��dr),F"� ��ZA��pa�+��21�h(3��F�67�-P�<���֚�/�R�ٕ��Et�b�ϵ��i�j�B���?�'���@d2M_��|�h4FAK���΋�U`)�u1��l�Yk A�}ج����8mVe�ֈ��N�\d�p��5Y��%$�uT&�R�s'��::7B��������������Z��dA�t�'Y۠C�L�$�a�H-�y Yԋ9��at�C_�����n�~��#,N����o���W�:o:
,���?��)S���fJ�o����nC��4�����09��[���HFA�]�M�N	�\���9s<TI�*��B�O,w����Q��e T\*ʞ���L����G �J��Z�p��at�]�C@�����#r�i��ȃ���7�l�)9~D�RGO�A(���Z�TV&�zo�̚��K����I�l�c��C���l:�!��@�|��<��_J�"B�� ,�������ko�U�]�,�Fo��SM����d���d/tE6	�>'�@#�vA�h�y�u��D��H�$wB]�ި���t*./����7�,k�������������@G��_�k���ϊ^;���=�e������݅�b��V��(�I�_MQX�TR��t��z=?q�ܷ2�,q�ܜy�s�:n���b	%=�vt�w�u�,��e4�V;���#�,��`��z��$G)*� �r-�Sg�X+:o5��	YӯA��&�H9ir�1�1���n���F�υ�z 6�(��D�\��<x�}}R,oY~������։T"��;w��HFyzT�7 8<�Q��P�͚*A�~�����`�V�Bp$(HQ���Ji��O��K.�T*�׋�6�����	�ਮ���F"hM2@d��YUQ��fE��S�1�%�������mї�I����."�yQ~�ȡ�e��n��XЏ'��n�z"Z���,�{�B;^x�w�bٽc'���*��W�Bog'r�<V~�{�dD������q�������!�WR������\V't�U�$��X\6�U�>i��k���Q���Վ��K�hD��-izTGp_��D�5���K!�q�C���-��>БӢ1�Y#�ˢ�4���R�X&�l��	�5��� &6��w��لT<"����X�a��zг�����:�X��r>�'ZOb0��[)�;��Hv,f��ǂ���)\%���r5�d�qY��Qy������EU����3)Ogs�i�h�>D�@F͂����:I@4����Q��kݴ�`�iF������.׬��ә�$K!y�u�dA��0�J����P�D|X����&���@<��d�̩S�s����78��m��@���QpTT!�/"���\�yR+��I��e��Y��85���}-��̈sB�X���Eq�R��즩�V�B��ߑ��u2�a�si�s�rܼl)����"�LIg�)`wx���7ߐ��Jkȹ�^"Nonڹ�(ْ˯�b�g�~���􆢰��������`8��v��ʃ��QD��Η�hp �0{�puZ����Y�|)Y�����
�F#|���iI���r��?���vlG_OF��d�V�)>�7^{��a���^8��'N"M�����.��`_/
�8~�L5J�qL��������w�vl۾]���0�y�
I:"�DOj�������/�|�����-P��2;1�⭐ɜ{��o]PC_PCé�'�^����v�P�Z0L��~N�|A�T����-�b�����Ĕ	���}���B?���H��wx�K��v�^�L������X��&��\2c._4�]�7�g���g ��悚/r:�H`XvǏ>�%��;�U��]��ف�{�ݽ�C�?8��-\�H&Hv�}�w��tz1�H2}W��tf$r$A:�L�� ��H��4���/� je5!��GgQ�����yN\
�*}��C�@K&	Ij����c5��)��{�´1���m��z��q6m�@0�=ʿ=�\�x�R��tИ�B��p��U��e��d�XpK��O�]9���4�ɐ?���si
�*��/���_V�?��e]�gl��8x씸6:뚐.j�ߢ6ZP�	�Z1֐wL��Ə��4��r��N�I�2��랋���!�6<W�ʆ5�I⺥K�<��ӏC{�#:2�k��K����NE7͜����˻�c�vL=O��_Q�q�BG;>ټ;����p@�A��c�(��}��➂ZMS�(�����0���v��݈��n�/�m2M΍�3��w�=H3�#�m{`8��n�.X���$���S�AԈ�#��3���%�
ڞj%�,"����U�b�!I������\�����2�&�4�*��� ZU�� F�4���o��R�;;�%:�w/>�9ӧb�������p��y��lF�U�W,��jKX��(m�e*��C���۷o���V� �e�^~F��'N(ˇ38{���U��֚�0a
4�JĊjd5f	K�0���˳��g���kR:�p6�Kj�p����I�͉�J[N7�2r���U	�!�O�aJ�N��ˮBh�[�SfNG�`B�m�#���
_~� 'Y�f6[w�ƪ�7"�)�ꮂ��}�	�2�K'�:%��k��JAg�Q���ڃ����ݵ�e����FHq�VŦ�?t��偺XЕIDx�~�Y%�Dg;�&�Y��ܶ�}�t����۔40gz����ٝ���Q�U�hG���S���c$Uj��}���e�0;�0�}�fBg�4`���yx�4�Ɣ�&s���5��+���H	)Ca�}~aKE鮩�d��OŴ�5�1�߃*�W/Y�����Y�%b��uk>ׅ�#��M�ȇ��3�;��ƛP���EuW� ����U'�^q3��03��aB� L�e?u�H:3��"�F#�͝-�9��f)yL�<�.���}���6������	%k%�1���-�ڂFL����l���^��:��9 Uv�Z��h�XU%$I�)�3�؂h0 �+�XRv��t_��n�Ԅ�X8w6~�DK��ı��k���`1;ffN��'�z��!ES�44�h����3ȥ�:a�������8~���
�(H/�}`����je���55�^������̝�u?�[﭂���N���Ȗ`��0�q%[�RB'č�T�{!+��tG�%��g��8!�r�P�FC&�W�59Q��n^�V�F�v��O��
;*6hr9L;���7n=�\Q���.L�>w�ur��/�`ͦ-P�(hH<BllV������.Ǉ�>��-[୬RLu�����a#��MPuU�X�Z���
�>o��Ŗm;�������S׌4��N$2482ʂ���l�d �ӛp��H�!aE�%��Y:�|N�!<S����$aId�7��zz:J�Ë/ <8��3&��z�!?z�:�z�:�Ofp��	�v�����۸v�"l۱m�=X��I�ղ��4�E�hL���/��~�7|�[�U&6B�V�����z�}�lv�j�T��y���1��IHkn{��6m��]{᧲��C�>�Z ���7���JH��^Y3�hh��N�:��� �k�LJ�)�k�0i�h^���pP��U^�T���������X@�+�ذy36lމLA-���`/�_w{�A��$�I���J����S=��6݅��ni"&�jD�ӂ��������QY׈@4,k՟��Op���fP�#hh6'��#_��XKsJno�u,Me�9��8*�[�s��I �SQR,����sCD��OPW��.��Wb*C��Z+)����}��1>��5��+<�P��1FD�~ە�c�5�c���@��F�I�������
a�'O<!�)6x�
֬߃7�[��� ��:T6�H�	�
��5 e��-��)\��
���)��O�N�`��%�4�p��.F,��q�]a��t.bx%N��$ �x�N�Q?���
7�-�[֯C,���E�C����x��Ԁ�d�"���O���}R�����Ҍ`8��h2]2͌y2[�i��F�Y�����N2�XX �x4�Ńx<)]����}���9    IDATȄ@��@mCX8w�L�,��ZR�fN�!Zl(��y��@L�p@c�Y�$;�pW*Zg�/��Dq�cPC�?�TQWUL�d��x�q�F����l�XL1��L,�?���I��Le��k���%x����V��#��c�,F����䪬��S��6�	CY�&،ɷ��g��l@��G��"Ȓ�$`���HG��=2�X4o�b>X�>�L� ��HHZt�gO�_x*j=V��\���P��"�N�̩������a�ͽ��Q����(�����Q�&��'�	cF�_���ضq=��+�Bޔ�Q��s�^фrgq��)ddWI(��g�ĉ�����3u2�٨�[�%r�%��GM�[��w��*�7���̸.@�(_��8}2��E�zh��` F�s4:��1�7���d�[XFb!ͺZ�+��0g�d�kl�O�K.����'`sy$ ��l�5WBU�aۖ͒��98g%J*�����}��8��ކ��N��6�/��Y�!|"J�PdΜ�2���!YY�0�K��./���Ϡm`1}T� �ѣ�7#O�F��v���d�˺�ɘjdɹ((.},�
��v��@�29WX�2 ��>�.�5^'�47�����'�s�,�p�X|�d?�Z�
[�mE����@ۅN�ttbҘ�X�h�X'2i�w�\[7�C2��6 ����C���i:|R+�[�
�s�`v�ȡc8}�����c̘Q���J*�}z�9̾t�<G?�տ#F��E:��i��k�$�6
9��.�l:�^��buB���Bx���y���{\�@,�I�V�0��)22�|:���j��I4�k����`�XΞj��næ��p�TG����;�'��n�a�?�X8�uk���\;��:���ظ�t�?��̟�G~u���;%���-��}�OX��475 
�9..��O&�"6!��c��������fh�d�dU�1qH��0	���:Τ3R�S,�Ez�Sf\V ��s�H��ff��wS���a�ˆ��N�����O>����Q����I�
X�Í��ge�b��Cd��}�a��IB��;��:�?��:�°V5@gqCc�![�I�Q�_�7Q4�D/j-vo$&`1#�}ϯX���m���[�M[�y�k1�~j2���.�'�$���+�$��,��Ka�X����_��*�E:B:�A�B`�-���C�� �јs�^�M��H� ���>���Ã�V}��Wp��]���&�S���d��d=@��~4�pUT �L �nf��9��l5YP����"J.�F�\L�[��@L�8�V�ƂK� 	K<&���t���ȁ����G$��R
Bм�ͦ�ǝD	��d	��I�l�]a�I�*�����$���P]S#�3gNbh�Od(�Nd|��L�0W\�XaF���#��H,��3�ą���+Z�5����� �_�!�̔�l��E��H-x2p�M��uk	��"˔h� �O6+��u�L��i�ƌ���Zy�C� V�\)�|���F�8��ܯ�mc��F�y�I�Z����hI��-�K�
2$���[]����[�xK��J;�*�ܕR�$Sr:��s硩�IҼr"�3��|W_?��44&*�k%3�8�$_)Nq\�p�a���L�D�F��e:iq��B���7��f\�Rf޻V�J���/Dww7Ο?��j��x���:�q�*�u��HJ�Y������@4��@{F1�ˆP�yy�l\��$�Y./��<�r�8+݂��<�Q_�/,�q�'�� 7� ��w��8������/�ԧ���H���N��
Y���Ű����6�c��.���z�X�^2!/�"�!�Pٴش;%A���B��S�'e-a�q��<̈�mB��=i,��CsC%�͝���|6�W��x�pDP�p(��S&`�9ذi;1� �P@�Y����p�e�GĻo���Q�ر{���h�)B��aV�>�O�xܸ�[��ӭB���Q������3Y���ǅ�>4O�����g�ޘ+T��.Yg=392$�r?,�4��]N�gA �b1KS�g��X���BC�h��3���%��ɺФV��[-���`R1���>�x=TF�4�;w�B00��Z��.̛u���>�p#R���t�+@TH���٧1���wlI-M��E%"����`�4��,��<V�|��m�o�^�?����_z���5ɒ%�V��D��9�5��'G�.y��s��\��WT(*i,�oPy�բh�9�5�y��u�Ѣ�-W^!�j��m878$�إ�����P@}]zBl۵G��W?z� �j5�_�&�ӦMù�lݽ�z�)�a��Ac��Z�x|���qBR�I&oq���щ���<�P��غ�����P�$r*��ٍ=�t�sWI�ϒ&aă��@�92�S	��Ã�����|��H7�-�HRIw�i�Ġi&HAw�b��g�^Tx�B[�BN4�z�'iw�]sI���f���XI�e	����[-&	^��$�*����*�0S��`E���s1��Y�]�x\�X�w�Ŵ�d����u��L��"��+�x���$ӓjfUs}���bG ��?����	Z�ٜ�j�j��J��(��T��2��+ΖL��g1�ӅK���KJ����w���;v��'��{*+��Գd"'v�L�Ӫ42�ID"Y�&=bT1�4b|B���Ȅ-,PdDi��e����(P6���z�51��?oƎn�ɤG_**�x��W�	�O�Q������h�))̤/j�I����'�i������Y��1��,��j���-"ea8
N��w��N�`�:�wǍǘ�c��(X"4�D>u�H|�D���Ս������F4/"�Ay -o�V��#I���ԋ.4�\����b�ݨǊ[�����e˖��;o�؏� N���_�h���p�ş�+��'�|,F)�I��� 㖶��%�*�[d8,R�DH�PW��n�bOe�7�ń������%q��.��r�V]=ݰ;�BȪ��p��I�p��!� "z
v'U��f6/]�f��I/0;�4y��b���;"���ϝ{>wlr�x���I��{�q�4
����J��a9t�>�*�O;9�9Fh&v�ъ'`�M�"Il|���P'o��?C �%����D��&Sng{≨�׹�6��'���3��F;�b��>lٶY�.��@D�x>��Q���:<(��H���}��sC�5�bZ��4���$(���(`~�Q�	��i����`�g�?�M��61"���rB�)I�v��)�
yT����q����o���!?�t<�����.�h""J�OoD�E�nj���FBu�p�+`V��vn76o�����e�d2�@*�@�	��,n�en��f<��ou ��Β�ݴO����G�/94;D��t?�&
���x>��DH_g�H���;ׇs	�v�}��,��"�6#b�$J�<,�F��(Fp;�A����]},��@._0{O�i��8$����Q�K�]�|A,����p2�HAo�D�]U��;w!��š���F�I�Nx�em!:�������^�oO�om?0c��ݯ&5�)�RЕ]=�RiXC�le��2��b��uN>�<��CAd�Ja`�hw�D��]�Yv����r���T*�Wz�[<�L	�"lB�2=�Z���T4Z ��EQ!�h00@cC�����Bc]���K��.��%����u�d��᫪����ť�/��];v
,z��W�W^��ko@oW7����N��@��3��f�O$�����%���-�C����gJP�0&�G�+� �3�$b1�fA��hG���a��D&�*�MvE�� B�!47ԡ��D��MwW��N�[�Z�DU5�B<I�2ШM�G�ttob���T5�#�.	얈Ea��`T�a�1�!�@(,���f	\#0�5��?~�[�	O�@<�0��{v`�ޝ���[�p �T�1	���N��(Uy����m2I�J&at���dFR%�f�C�p�[�yO&�Щ�ª�����<�1�Q��$??G	z��G�R�̜,nh��Y�	�q�	����]!�a�2�����)����T�*a��QH�e'�Md`�X�3�x}�]Qp���$f_2�<�p�>����y�FL�2��~����mp���)�Ҙ�W��XJq���'���&�Sdu�N	���\�� ��NQ���i�������{r=T�P��.�i���P��"�N���������������"�N�d����g�K�p���@�D����4�t���9�G��<�B�$�E�C�Ų|���I$-͙l&#�\<u�5صg/&��_��ߠ��aP%���.e��<��>+D��D���U��<���d��8�#B�����S���4a��($�rơ��lO�w�J���J�@��U���A>;9�9�?zkk+F��+���]��Γ �$�TV3���)W�ÀRdZ��+,�2�h���98�Z+g0"?��aFV�|�;o�#�����5��CW�_~�-�l@ׅ3(%c��2h%?�$��XV��h.��d
.�U�"8䕤�A ��_U���l���h�񠷳]��� ��ۏQ����}tblSn��.�^���N������B	�D*�����7�%�L,��	�!�����kE�2։�/�좥i,*i�D���Q�'�a]���cڄ&��PaP
s^��֣�q��y�9�t/j��aB���48�&�@5U5�(�q����Zh-�.D*�`DE�8�6�`>��L��]�a+���]oe��I�g8��,���7j���2�d��C'��_
���}n*���.��(J1_a���y� ���*��j��!.�fL�tǸL�^����A�Mf��T{܈�B���p��IT"8��sfJ�4��&�Y`=�LK(���ӝ���Ì)S���0�7(���qc��X�ɧ᭤��JP�H")�4w�{�ƬK��ʫ�a���2I54�a�ⅲ��n�����V�ń][6a����t�]R���b�C*��!=�L��	�L	��f��fq&e&L��$���E٥�m�w�w�Ȝ��N�â3�5c�\���lhJ�|}C�LrDT�Ö��}��%m����ڄW�؀����4W�B�%�^����#��J��WءJ�F����Z�{mu�'Lf=�;�c���S���t8��pPЗޑA +FCAT�]����h��'D�^�'Tj6 z��V<�)�#�()}Y�P��ILm����j�IcB�Fr|��j���s�_�|�1LY��N��;=��1�$�~�ؑ��Q[S�Zo%���Ct\��/���Q�C�9y��±0f\z	����hlnQX�C~̚=?���n�`�{�u�<NI�b����xT���!�Di8�S��Ʃ}����F�`CZmFQHW�:@� H��i6�,:�Y`��%!�U��dL�k&���G�,ݴ�������������S��R�8�����VS_'�4����т�`P��lz=RY¡Jä<�ji8�{���ʗ�*���A�?�'��m)�� n��6<��S��4p���m?��(E�DF���������$�BU��H����:��u;�dh	I�+���`X��
4�ʦQ�����/O�ND�j�Ϝ���fA�h=�w�.9?8�gUy��`��	��,��������g�cl0W�4Gbv<�w|��3n�9g`�oB�]���Q&˕���o�� %�.ĢE�ahxXxG���[q�-7a��w膏�DV�}�aTT�d���Y��J���BH��0�}� Q�p9b��Ø�Z���ZN���������^Qc}���e1�w�`T�Xa�W�<�� �p�T+δ_@"���n����dj#QI6@�����Q��޾>9���//"d��kV�E�S�����'aӀ�X1UU͕�q��8��c,�:E?Z��[���/��֎:�	���\�BFL5:���r��N�����v�Fw���##,�:d�J��!��	]V��D����+�;u:�`��������[���`��W�:ˤDI�t���B*भ��	��JJ�R�h��Vf�B���Mf���L�5q�)�8�ӟ"���V�A"AhhP|�k��pP>���.<;Җ�:��ø���n�R9�_v��
���������[�����X "���'Na�)Xz�u�s�m&��5��Վ���������0c��\&t����2�{�vd�b�iطu3�;�Q�$�p��:�@�ܠ�-=U�֎@<GU=r^���.;�����-�?��	���2���Ƒ\����v!���v����D�E0�BoO����LR���|��ZO���c�1g�t̛1�v�ƅ�gq��!�А��j,�;F75�i�(��>=� v�8�K]�Յ��/���D,��M7��Ѧ�eECh�ps�� �����уhinBp��%�].�E���>O"��AE�Q��x��ېU`��@�{m�4H���0�P�I�֤f3�A�zz''S�V�B	��=,zar��b��#�f,h^�sfNG.���F4�0����8,����PP�K�յ����B8���N�{O��'ϟ��o~����<��KbaI؝�
S>\��8E���$ch��!��K5�|��-6�u6��D����P�:duv$�F4zaM�*8MZdQI�'1&�щ�dV�k�ģ�l"!�P/9Iibـ[�6i$��G{SNҜ���'o�њ,�XR{�9���QY�Տ�V���n�� G�2����7���ĕ#۵����_~��^��L�ƍ�ر�q������u7\���z&=`A�x�&�Ǣ),f%��gL��d�uU����:!^e�F��tF���F�PW#�	�|��0�TԈ>9���^X��-*�?N��M ���T[/�\�#2���:"�]ND�q���d��J��J13��I�lVBWI��IԱr6pՖ��k=6AD5��؜r7�`����oE}�ҥ�TV�^�W{T֗�>ـ��_��`�y)�D����~1Ꮊ��˿)��d:W"��0�����&W�|f�wc#C���g��󂆃KNt�Dfy6��N�7_B_O?�N���c��='����3��bHd�bR�����H�%��6I�49�˯wy<����nA� g)������]�d3B�Y�-PYux���qt�z,�9]֩�=}�4�Śu#����M|VC	�dL��*�%�B�P�� *���1�D�t./�%3�v/R*#r%��*B/1�D��:K�*>��y1mMcQ�PLª+��ջ��e�e�}���Ov]������iKH�Q�,碬��.t!��5���]:�tRD�,~��� ��c4�bȡL�$�%�q��|�0��A�_��ͳX�G4�td7.�
K�ö�1B�����G��������J��b*#��V�Q<���
TTסqt�����e��e�������Ł�,nL�!��$���I�%K��&���_{'���֍�u����'M��y�bˎ�h=}
�&�����n��Y�Ov��$�+!�+�~�b6+�L|�Os*��Cr'�"�����,�
�CC=B�8���r�r �F4U�"��ͯ�j1��W������~�k�{�VL�,F"55�p�L�B�0fBd�PL�h�7��̸����u�<����G���]�p�d��:�(s���I�q��kP�sb�ʷ��"W��l8ŝw�-/�-�f�XQ�4
��\��'ΊG8#w���j5rH��q%ޒ�zV��^W���d%��,�d�HRȚ��D+�i%́k
�{d�bЫ�z<������iĢ#����[A��Μ9��s}���^4��¢W�t'-��j\y�?y�G���׋��&L�>U	�]���ȫ��Y�0��!!T6DU(��p�U"=�`x�W�@�ؘy    IDATgP?	�0jt��w����3�$�n��08=�$)j�A���s��+��a�OQٿ�`oi��]�U�%����&��=.ӥh����-Y�ٴ46�^����ա��Y�:zT�&ꪪ᭪đ���98��H5MM�5��T8�5k�j�p����-G�xg�BD����ҹ�<�ze/��J�)�ܿ�6m��iA&8���������_��\����cY�d&s�3I*���3|��ń`�/�k��Q 7@ȿc��:�!��֢��� :b0�3�=��8���XW'9�L1c.<���|,��-{zp�f�F�d�����dV�s���`� �e��YӦ�<4�`Ҋæ��ʬ���~\{�X��:l߱5���B7i*=&D�?Z������eW`�o 9��Ya�ۼu�`�F��LbXR5ij� ������ b����/�+]6��1dS�0���F�@Y�A
���Ʌ0����\��LU��Q�B$��Ȑ���i�B`�Bd�hO\�qp!ǂN9$:��ƌ+	�pP�M�]$6�칉��e����	ԌOC�}9.ڃ�3�c׎�8�z
s�,�u\>B����tEŐ�%��(�y�U)�B/�2�i����Fd�"��euϒ�G�{:1�QVL�/��3��Ê����l�bll�����8��r���?�������=��޺�Y�u<�O�;�F2B�D���{�rh7�W�X,���Н�6�E�<��/v~�x'���c�}#3�c1qú����p�Ԁ�{�������nG��#8qh�_{ƍn{$����ش~-lf|n��Z�Z�%���,�Bc��ЅL6\��z������������_�X�wW�GN�xE��n��L'"!�/PuN��:�_{�a�_�>Z����P_-/";�-�n��<Bʌ���üyK��5�o������J�x�`C�d��p��f�t�,�$���-5�d�C���v镸���زi�<���z,��j���`�ڏ�T���}[,1?^�!����عm3���g��ag��V+�Q6���n��i��ՈF?�M��-����6���l���܉%W_�o}�8p���:qUSi�<!`���4���+V܌k�,�sO�C���y�Q�e�)�]� CH�2���2w}�!��n>=x�:� �Q�XN(:d8�ӿN�Պ�DKJ�D��C�n[ 08���qcG�G�����1x$#���RK\���/����@�F��L����g�Һ���Lf�&��B�o@�E�4=�َ�P 5c[p�wb��m���k1}�<��o�z�&�
4�1��"�­`XM!�DuՕ���qx�n�߽�dZ2r&n��z�X}罕"�,�������?�����+o"or ^4 M�2����%�2W��5��:ѧ�fs O��!��@�#'�3����f�?�O��L[�bA|8������s���/��Sǎ����<�44t�S�DP?�V��1
E�WU���`��	�W�p��E���� �?�����B���hu��/���<� ɶ&zz;p٢��d8�g���p����Z(`��ْ"���^��i��� �	��zSyh�^�w����n��i�A
-o�Ɇt��P�l}ڭ����@� ɜ\�Q�b��GKs����;��T��Ok�`��|ᦛ����b�$���ta�}صo���8�zaߎ����1��9��wVڐ.d�t����oo��5�����e�_���t�`׾}��p�ǌ��5k?F���};��|��6An�S�W�F'����ń�,N�y52j'��)4L��9��/���J��i��irJ�:�1�N��FW�BNLXؠ�b�B>�������$�0lV"�\2{�O�$י,y��k�����Lq"��G�Ȅ��(��)�����I��0Q3"Zá�G�p�6@m��K_�"�?�{�0~�X�C'2�d�FbadbCH�{�4������K������3"�Z%K���j-�[��ஒ�!ew��%�_�Ue��t���'t��Y��[	8��z��7�����l��a���3j�8��N�+_q�aV-� ���h(�_�r.vTe(^~/�����p1p��'f�o29�UU�����Y�JHVL?"[��W�s���X���s�M������H�V��ZO���-8s�FUWb��W!
��d��;�t
:�gj�n�]��ڇ�D���Oćw�?�
��R|�i��	Y<�����E���y���9��.�=u
��s���:�d.%��_~Ed^�'L�܅�!�࣏?.�'yJ���+9��P	 ��]�IN���Dor�	�X�x���tw���ʇD,���G���ݸt�t�;y�����<���N9v S/��S�'�u�FԺ�8u� �:��_��N:������j���
[���+nB���ƝǱd�r̿j�|�/�q�0J&R�*52�*'X>���˄�p0��/�/��g��2�E����.ÌiӰ{�.�a�9Y��C��N�,����K��އ�ᬮ�@�C��ƒ�'WD$k��g�Y�����(cִiB"Q�ҳ�3�c��Y���y�V��w�w׭�1y,^���h�̻t����$b����� ���jءF��	g^��4*�.|z��������5k����sl�u������DNŀ�ro-�JZI2�8�A�/�Ϣ���K/
��qWCekbj���f��	I����/�VU�W�[��ڈ0�S?Wh�P�b�d�|+�[:iQ�Q�����d,��jjjd¤Eosm-,���dz�|&����uUX��=��w��`d���o�ɕ���-�h���)��1��.����X~u	�Q��n@��	�&���/��N�F�l�
ҁ���X��n�dbMDXq�uXq�R|��/K|)�(D)q���[���){�s:`2:����G���{���_\�H��@�/�+�э�h|%B�V�&=��fH��Y�X��*郪F��8��Ev��:�N�on��<�"�*2)��,F��@E����ʹ	5ۥQ��]X�ч��͜>{����s୭Ƭ�3��x�s/�"��˔{R�C�����e��\��r�����O�w�FhK98�8��u�c܄����+�q���w�̔e�o�H<��m]0x*�U餑T洲6�����)�J|�ȦZ1�)�g�7�0�u�=�oj������2m�K�B���è.��ѣ�<n�0����"dď-[>��I�C+�Jyi$�;L���%�%6 �X�CQ���?�d[�$����:)��!	c�	S�E��vZ��c�&9�s��4	�5}�,QE;q
]]=�,�R;y:*j�����	��"Hl��R����K�3Lyꔀ:��|IK{�,�bl������4mt��kB��7�m�KVm�JR��Rܭĭ�	t�LEC�����)��?�_�,8�
U3��,�"�L2�A<�sr�bQ�����)�q鬙������{E���c¸1�2a,6�Y�/?�I��� ��V�_�|2�|"�&����`B}=t��Lݢۗ�Q�	g�Ķ�{a�zp�-7a��F���x��a0������B�,��M�ė_wƷ�E"��c�ٸl�B�0J/���{���0[p�eȕ�ذm7N�<���3W[�<r�Q܎��n��IB�T���A�����B�͏<�tz5֮Y�	�`�q���p�{��?~gOCW~��w�u�<�}���q��|�e+J�
�8�4�FSE%T�4��6��j$0g�#�c!,Xv
z�j;n��^�d�_�6���Ţ���Δ�x�e[�e���ٳq�5W!�׉�3�p��Q��g?'�O�oò+���CGN`�Y�i�I���/o��O����B�Nl|�ʵP���������sgLi��F��@@�s������
�{O|�֭��%3�a�;o����������ǜKf`��f���_��O#00�B8�E�fb����f�h290��.��j7�w`D[�]��u�پ��1�b�8z�/���"y�^���$�-�d�KFa7��_�P_/��ك��_�V��[طc*�v̞9O|�	��Ӆ\�cg��ӿ{i��ŋ��N�d��S�ب�x����)oe8�b�`��g�,���V����f`��c����02؍?�]T�l����q��1�p�n�5ȹ��q`�>�N1�z��ВȚɣ��F��p�>����c��͸i��xg�'�v�(����\2�0<2Y�ºf���l,���g�%���sO
�[0m�d\�dv�؎����8x��������'~��?ڄc�DC�+j��@"�yB,E<D6�����+������XƷ4ɞ�����[�#@~��lD_���Mjn�}������C�{@�y����e��+0��ޫ��&��DG�lo��lv�M�����v�DRL)�%YV�V�V�H�Pb/bE! �����^ֿ����s�9� 	L����ק���؈Rٔ�z�P^ַ��-]�m�~���j������Ju��)���7k��������_�ˮ�Z��m}�����=�b��=`G&���/Q�џ�hD��;}����~�C=��i�7+��jEk���t�E�u��)U��z#ڵ���?�7�b|��U$7�F'p��S�|���vD[p�H��D��h��j]��>ǝǎ�4>>�>+����_�VB�]�Ho������JSǎ��oM{D}(��� xU��z�ݺ����~.`hb�qR�m�@�M�c�)�|�R���9u�'c@��v%+�VC�\�UW]u�>z�G�ۓ5d?8��y��� �:�z����l����xZ��A���HW�#�S�Y]��Cү�z�IH�G{?������_;������?_��7��(��N'M��~m� $c�\�{M��ڄ�.�˙� X�7ې���9�kE�&eth�٭�7i��5:��^=|Dw����c���k���}J��{t����~�G���z�aӬ�$�z]������K'������f��η���K��;~CϽ��U�������6�?����/V"�7�2 ��V�r����j��:Ԫ4Ԯ�@�ҕ�]�+Ƶ�0���k�Է��]��6oݦT���zTsK���l�_)V�6��_6p1�x!<`�4�ue#mg�܁��t�e��g
��RqQ����{�z���f,V�?��:��~�����T*�-�G\đ|�Fr<���Xi`�0ɞ�^�:�Z<b`\�؄&7�����_�O�Kz�gԏ��R1�LDY��CU�iB�n���e^���4u���N�4-p��M���4B�s���n���h���k�+�飏kTf"cI�$�Ng��AbGA�K�rq^=)|�v{�[����MW]�Q���?�n��_���=Y��mo�?�y����.�h�����G�� ���?��gϨ���ɞ������/��l�U_�G:��@A�۩j.��S��u��o�^�����_�:Vl�j�'7�v���}y������Ȉf��Ѓ�oܩ�|H�+&�zr�>��Ѧ��u�wj�X֞������X�H�	�]���;�q�vÜk�x�����BH	������7n�Y�/����^g �_|����;��'?TqvF�o����z���i�3Oj�p�v>�����/��N$j5�M�W����X"��h�g�RH�x��M7���o���u����������j}9E��Y-L-i�oH�ڲ*�EE[u�q�-zÍ�����ƹg�����?�������$�/?�)��c�)����;ޥ�}��:tj֊���xz��]��v.��ܼ��RȈ:�7Ǥ�^V�����>�\s�U��W��7���ڳg������������s����m�efg�~�:�0|Y_��t��:��1�=xX�����'�z\��'����gzr�.���[��d>�_<�W_�ڷ����w�ٞ�W}�1�Z�vj�e��eu��ߪ_���������Et����QO!��V�O�R,�ԓ�������?��N�/�s_���'֩�0�]���iG,��ܫJƲ+��+�m��i6590�/��w�m�؇}D^�ݬ�cG^ѣ�<�t���|J{�}R���
�����7_��}�I�\S���h0����z��̽��?t��e�{�'t�5׫�N�^gn���Y}����ν/iWQ��q�͂(�zAN��������7�A�����U�����^]�^�G��ޯ�ۡ����m�@o��}�{���}q37?�t�6��Y���nx��K��|@f�����i-����{�W����?{���գٍ��`��hɉ��ڥVP�
O��¯��?L��<��e���V�*�����zDF�N���W�l���ܪ��1��--�ꁟާw���z��ߪ���/������#�v���Z����А^ڹS��c/-k��Ԋ����kr�:M/���ܴ~���S]t����>�g�ݥ,�H�%T�RXq("�{'��,8�ח����]..i��A=��C-p}_9vT�V����B��*h�z�������8����zص�J���Zղ��zmͺjr��m�b:��l��];t�y���?�_�^z�z��:v���?�?�n�*�q�{Q�3~���<d��|*�!�c)��L[ c�mZ�e�^>~D'g��S�X�F����R�����#����e���&�t�-S�T����^켻:�&�pӍ%�=��G{���q�1�H�X�;���{DMQ�~���^�#Al-�U�HP������Q+��������.rAq�����}��_��箻��}�z��w�w�C_������3F����_����(�՚;�ឬ6�ݨ|4�LE�&t���je��q�7���q����koԝo}�����k߿OS��E�wC��Db?�VR�g�h��r�uZm:��ߪu�6��HkW���w�����k�*�k�ˇ<j'�#��@E궽&���A8�^�N�ؔEO���'�*o��׿Nw�q����޷������U6�ӧ>�W��?�#=���:s�������V���_<�o��W�83�t"���T1K���-N+�lh��\1��j%-����[ubaYW^y��o�H�����5ik��qI�+M��*������8��ccz�^��#�ٳ�E��o��܌�~E��{�דO>��~t����wk�R��W�u�f�A��΅'w�#��Mz�a���J��#o�Ī��6�t͕W�=�K�����.����]���'�}�y���+��/Io����曕j��jسw������<��=���]�V�����ɸY�U]=�g�^�����J[���wޥv����G>�����z+j���ܼWY�F������O~�}Z58��{�衟�LW_~�~��[O��q�'V����kv|�-�k���zf�K����d~Xu:t�I�v���#q�ޤ^��~b=
<0 [�#��n�����ӑ�jV�%ǚ��7���~Ww��=��c:�o�V�i��a���U�^����~�0�*����b�&���� �QA�vS��N{]sۻ�֯���e׽N�0����;��X;^:��R�w�{a{ ���P�+{R�u�y�������j���m�u�e��]oy��Ɔ���s/����R*��Ukt��W��ٯ���;�%�#p6y�*�'
�l7������D��	��a��o���O�ڠ����~~�g��,����F��	�*�o��
;��1���n����~�w<砅f��#sgg�p��%c*�I๋�B!�sR�
�Ƃ�����;u�������GT257��˟߳{�;�k��J��o���C�448�;�~��}����II<��o�]�k��G?����8�d"cp�S k���tqЛ��*FF����޼��~V�Q�c��?0�Nc�ٲH௮6���c(M�R��o��RD�[MM�����`p	�r��CfP�@C�sb�
ڼ���H��_���Ɔ��{��ܱc��Z�q����:�1K�    IDAT�����~�k_Sy��\&�b���z����J}����O���`#�+����_�ȉ3������7��������"�n��}����N�L���Fms��0���H&5<��jq���"�j�kڐлX�.n^'�� �
ZX�"�r���m�ݬ?�����rQw�q��������}H���M^e����ڿ����5=;������z�=�rm��U�v�a���]�f.�ǟ�`ǡ��펷�7ߡ/�o�����Y�i�t��@��t�V1S��� DQ �k�n���Uk֚DD���+:==��'Nht�"���1�yR\�:�R!%��D[NL@([|~4	���	a�xB06�'}Dׯ�(#�o|���������o}S�<������X鋟����|��w� c����=Af��0 �7@P'_9�d���⒢����\���e�\��.�F�|�3:p┊�fx�i�Yb��L�<�C�a#����ԕ��1�v����͟Ս7^o�ڽ?��|�<��d��,���j�Z7�Ӱ�zd7��~��5���0ivw��ؘ��}�!=�-�{������G�z�
��ͷ�/?�	]��<}���{�Y�ݻG�g����Ȗ�4Wm�P['Wk������@��{�C�"5=�J��z�F��Kt�;ީ�ZK?��>��/���)e�GlJ����P\k<7�iC7����1l_za�����v�|�cҖ�[��/|�l�K�y���:p���:�X2$�׬B�������\�48sAB�\��c'��s����;��z�n������������с/������ȧ�fbD�=��Nς�X�`*��\V�_s����-4���1p��z�gu�V�Mo���ц�.Qax�7�3���^سǀK�5���'����EϪZ�~����jP_~q��<�+��]wi|`H?���z�-�j���_����;�������}��t���̔�A��}RxV]��С��ɳ��И��1�*���7\��_[).$���GS�JKU����=j�ǃ%�p�����]�.��<��]~���x�3�^(J/9�TF�&1��}i��d,��@u�����J��1�?���i�鑚�Yqqa������z�a\�C���3�	ųF@qA6�=����"�R��2�5�#q�C�نNE��!:ڶ���ҢU�@��X�&_��Җ�B.�� �Fi�gh�2�~�zND�8�3�N�\������N�,Hl�y�@%W�%����������~z�M�U^\� I�N?�v����n:��L�3�<����C=z����:et9�P�p�~�y��Yp��dFD�L̱�G-i	���Ϭ���!\�{a��Pho����1�ך���bH�V�]�=�_Mꡨl�1ѨV]a�u�0���\ ��u����_���GGL �p��|@��r�n}������v�|ޅ��Ƞ^��48�g��UW]e݂�/U>�׮�vi��M��;��K{���1�x��U���ku������}WO�ܩ�R��Й��/ܗ��8��l�A�Ĝhw��!������L�f%��S	�M��ѩ3�b��#��u�
�.�@E��i������#�����~���Y9���~����oi`hȜn���?�>~�G���{wk���������x�|�=���+�4�R�Y觐���M[�̵���r긊�N�-����:����\/�;`�`/VP���5�2I�'�x~�6 �81 �����i kA��ȉ#Z�n�Z��V���?ʕ	ډ+���v���B�,y��x-��օ/��JD�����?�}Q]z����O~�+.�T/������m�������ܾM���}=�Ѓ��..��|��P�dB�x\7_s�F�=Z>uF󧦤HC�VU�fE/MS#�W�ʕZ�v��z�oj��m��'>�G�١��E͕kj���r�#E��(;��_�-�V�<��fqYÅ^�.��+�a?�bŤ�Kz��]��cx�:-Ԛ*�X;�5l=
�$�v�#dάG��2��,6���v�Dh�~���M'�T���������k����c��7���6�^�����瞵�#؜H�����L��m6Փ&��Lݣ)��7m��k��+s���Ϳ���	;��/|�oL+-�.�[�v꾆��OOO'�����ܮ5U:;�����-6j�Ν��K�~�����nf�]���E��e{�^]Z(zʄ`Xw�n�7��Cn�`��F��F'�/���˻n���/[3|�M3�������pӣ�_�\+�^W.֜�%� �P�(\���^r���ht��&/��B�zu�N
�t� "�����܌_I+�ꇑ���c��پ��I��9���Z�ұP@����F�Y,�]uos>�Qsz������/�y�	!�d*���N�W���N�&+���Q���B��#�F�R��=;��HZ��-3��j��_!�=l5;�]#Ϗw�el�=UP���e7&�l�Y�9�0� ��OŃ4.�h��z�ra�P�(���ј>u��+�N���>�񩓧Փ���' ����N���h݆-���'�aV:b�E�Ie3����֖�XA�B�ϕ1cJ�k�T�m3�8��Z�E���K��vq��|�NP�P��)�����O�:���5�,��9B�:"ו�c6_��-8���U-���J9x���yˡ�eP)�5�;�=��iI[��KEN:Z��c&&W�壇u��i�bz�N6�G�bvP�T���oc�i`!����$��&R�(�-�\���8����b�G��?.xB��@k���]��E�Yr�ĄBg��1.�Z�b6s3���VD�e��(�Vq����o}�;etϙa�388d��#G�{�r�[���[t���zO��7k������sgT!�fҺ�o���
=�ȓ:~bʨ�V;j�(V�\b��ړ>`s &��@�\�1e�u!P��)�+�u��jE�i�q��Z�|��=0��=y�z�kǏ�R��J(�1��nڴI�_~���D������*�<�:yT�����ګu�W���~_�y�{�ן��?~�Q��<����>mZ9�L[VΌF[�Y�Uz����*'RZ�~�r}�����Лn�S�����{�\k�Tk*��%�c4�Ų�v�iG=h�L�j5����Q+��X��Ԍ�Ku��i��N��z�XDY�X=���am��L����6,*��Joiv� bk�xo}˝f����wiy�M�w��M=��c�B�>~ؾ�FM���M���˞m�u�%W����R�b��r����׬�y�_�}'�뚛n�tvq��?��0��Z��W�&
WrN�_��))���o
0�Y�r�R=9�����������invi!�4'��v����c�IeĎ"f�*�EӠϦz3��5���u�����N���;?z�#�^�\#�Y[���$a�(U	�0V��Ԯ��kp\7 u�]���tnz�i��\��M[+�|�H�$x��r�`���X(�F.�LB���'&0;!ƓV�*���бߵrՙi��2x�$ul���$p@_�WP�����`�qӟ�����Zu�,�'/�	���σ�#�����>�r��7oYZ���%�txx��`b�I��7�&�\-��y3�+L788�B�3�/�fM	dl�ߗS:�PqnI�$.u�r���3��{*IF��~���������
W��cNx��gĸ����<B��@e!��s���BW[�_i��Jy�z���q���_�(|O���%ꌃ_=Y�Y���Mk�\:i���gRh��N;��\�ˤ�M��D��8��f3��\�,-�Y���HR��A��Ғ*5w�UԢ
�jU��a��wQ�Z�@�U�����x���k�+=rG�!��&hV����$�}�Jc��P��4*.B*��U�p�cO"w4�{���$t{-�"��4�]0����'L��� (�v��F�RV;�R���,�4x�+'V8��9;�ɕ��s�dsδ�+����D@d`�_��9��e��;�-,+K)��>�f9_����6�Kx|��t3Ʀ
c�bD�F�Џ]���3�tf�zs��I�4�XT6��D|�:���9a��vm�ZIk�k<K�hL�E�2����������V����&ƴeդ���/�ƛ^o�VX���O;�������^�TZ;�{֚K��W���i���r��+��V+'תpL���/��g޶ҕ��!��ҼPoA���4ծ6=��ݕ�@�0�v�e"4;=o��v4�����d��z�l�R=��e��q�H�	���!.z�V[�3j�.����{LRJŢפh����a+r�Ӫ��tۭo�����W_6cJpO.mUɹ�3*��m�fڽ���4X��E5�R�7�E���.��*���R���G>|���UO q��!1��4<�E�mm�q�;�+b6з:ĸ�F;`P�'������53��d6��hi�Z-`�j���!�{�a�jNOΜбRuB/�������o�m>�ku������]?�LdW5�XT�����bT��F�\V*V���E;P�bW\*Y:��B�'��x/�C�8�˽C�O���aپ�(��n���X�jZM#�}*d�*�M�=���C,fԖҙkE7[P�!)i���ғ$hy�YW2����J�����/-�+E���ĩT�AM�@��?��n5�v���Ξ���9�Ӑ�D>��)BLQ�>����RAE/��a��qw�y�s�ĉNgB��K���4����<cܶ�2�ܠp���ƶk���xA��_7��{����0�k�� ��U�Ɣ��MYo��τ�%:�r0�`�a:D��g�û�k�{W��L�`Г�p�8�Z$I���g���A9	V���@χ$d�J�x�Y2I�����pɘn�������q�JuED��2!��@�b���R�<��	�8
��2�%�)�NY�pi�+:iVY��T�R{�Ҳ*��b��6�^֏���" ���N�o�����kc�B1Et����-�l��l�)	ۖ��P<��V=g�{�~1��l�}�<��<-A(�↿0Ao�3�J끮�*����+s�9�$Y��Oΰ-U�(Fl������y�fEu~��)]�9p&��O�ծ��%�j`�۬��������\��P �(��is�9�ϜTŷx^�
�WHw����3��=k	�<��b4�V�Y��Ч�((��Y��Ɩ,��[���i�`*���K��l^�\q����_�R�hE�D*�͛7��>;s�]b�IYM����^�5��{�V��Z���4��F�B�eP��&�d+L�"A�)ןwB��>{�%���*o6�*��F�c�곆�x��:�g_����aR .��AW$�r���h�xwƆ7M�2�4� Ī�Y-��j���j�1Qm+I�7��z��QQ�>d�N���}��r��щn~�񔦧Nk�X���#-����<�!~uX"fk�E�F�"���'f,P���A�>��ܢ��&��	ɸ�-��x,�t2�8�ڢg�!�8�Y�жG��XS�Dki�H���r�e��͓'~����y��O�9��f<��m��Z������x���\�h9l�'^*��Z���6�&�w�0��Q��j��d�*��^�����n����ț��Z��P�zq��eͤ�I��E�{��C�H9-O�NgB噌�G <h\��qZ\֞����̬R��N�[g��t~��o�x�����Z!�R>�$b�.qp�	$xZ�-�F��펌���G2eS����E_��1`��wQ.���Ǩ|"������'ب�V]Y ������d"�+�E����\�0?���(��hg�D� ��tlzZs媲CÚ^\��j`x�E�"�R�NTA90�;f�|�X�B�������^��r,ڴ	�58�q���=1
�4"�z+ ��E��%��g�M��:8Y"��l�Ht�
5��AC<�J�����f�O��s�؊E�faT �r���b��N&ѸA��^�&쯾@�N�3Pv+���}�	�u"�ix������պ��W*6��[ӻ�L=��	�Hxu���j�N}�^9�w�����`���l�#��{��7I8�pI��vTlԭ�X+���݆Q*l�Ag3�m��蒉����X�_�aw+u�HF�JǲJ�s��-U[���|�����{�>P���a��]L���b�^v��:8���sG�ǅ�x@��_&v�wA�E�A>��J��ê��.��ɤ�^��@�m��Vrq/z�}Z��S���d�V?|����^�-]�e{�/���91p�`K�Yr~>�
��(�4��*ͅ�N"t�ݩ��@�㬃��HU�d�?$��ꪩ��`�FGG]О96�v��vUQv�񄛮z�� =VLK؝3��p��&�5[���� O�?����r�l�<��p�d�<,"'���<T��{6!5*��/@]�12�w�e[v>D'�K3�QyD��T���o*��YB4��E�k�� G��ܚ�	"�������	�m�y�si��W2�����&Ec*˞��
9�R	�k�|��Ϟ��E���;L����{\"�T4^W_J��Ɔ?����į=r�����[��{诚�̪F5,�٭�q���/�Î�/�� ��
�V��WW�n+t�T�\Ƌ%�t�G��si����ٛ�;wP�� ���\RV�:o�:]p�fmXݯL �:��P��R:a��7���O�Y�*�#�=�=82��~�����~�{zՊ�<1�í�T|p�!:x���T�`��X�jj����U�0�|*	Ϗ�Ex�����^%�DՓ�9 ��x�r�0N�.�9�GH�w�U'��V���C��צ5k�y�*m\;�`JGK�P3��3e0M�5��4��N�kH�;���o���:�ei<�}U��u�n�̻�vht�q�FRJ��hp`�I�t���E\JŅ��X�`�Ze͑��N}L�3z>�_��	�]��*4?���>���H:&�Z9�|�f�v�tN�6�^��+�;�*�0��Z�.`��� ��Ɖ/F�$`�y����v;��G��od$�S
�}��=��"�������p*LV3r�uQ�e�'���'�y�L��g�c�<��.+� �Y�9�g�����wA��ȹ�U��ja:f�09�r|h@j��nǗ��й� e��9��	h`�����Z(��]Pkƣ*R�$�j� ..��J�MYo=�ϪQ^R��Q�t�
��Uh�	-񥯯�σ�Dǵj�ɠ��v�.�;ŧ�	�"09���w4Tl>��5r���̒G�q$� 9[��Ҽ��Z�t14(���E(N��Z�?`Y_�W��G<�S�iK+��d"�SI��x���С`2�w�̭�[V�L�.���ug��{�h#`6�H����m��(�a�|��؉�ot���8�֒p�t�����W-�l5K+�XB�=������,UUo��^�?��S����4?$f0���z��dK��G��k���GH�S>�8��~&�TV�fD}9�b55�H-���!e�Ǵ�Ņ�Ј�I�.,�j#f��dOB�#��a\,���'M.kAŽ�s�
E��n3AcJ�� k
��0r��R�y���=s�oi�'6�ur���r�uu�X��S���7~x���z,�
ak�W�F��%Wڑ&�~mݲ�*SP� �T�5'v�7�RH~r:v�!�lg��ś7c�Ȼ��� �	��/�+;;Z͆z{ԛMi���Z�r��Z$(F4"�E���!�����QS_n����`o@��2��lF{��?���-��wc\,��1��h�R�d�F�݄�e���|�ctvۨM�L����ic��9H��G�t�@���w�p;��:����uPco�D+�=���jE�n?_kV���7\�u���$�Y"c]�`����^��s͎�Ƅ��;`Ҭ_(-7�����_�[ڵ�Z��r�^�R:S�5�c8�yW�۩�@Mz�8��>??���RqW[�L҅F�De�P<�>^�pN4�<: g/�,��f��C0    IDAT���mg�`�=�,��"MEaj䎬��ѳ/dҺ���u��t��5қ�"�'�}���*-���o��t�aM�&�p���9W�y~�~���zn�^t�� 	>�л���;n��P,��ϳ�.�k��t�%�()�=�S������Z���Ḥh�ɼ�xR�L�6��f�T�~6�ݡ�Lw�Ic8����%���J6�R�����&��_���i����#�����#S�g��T�+*�%~&F�����9���ν�Xn+���MQ�hםTu�U�M�V�SV��f�Ng�� /@п3�S^0v%&U�QLS8����@�lu��7d��sc�?�#��ƙL 6�)��{i��F��l:��(��O�yr��媖��hrtܠ�,L�����0&u�3{ЌƄB�fc�V��E�ת�W�T,W\\�&��ʚQ;�b[ip?�䬳�.nM����|X�9(j�݇�]����V�17:.�	�&-���Vhv�y�������=v���+;�M6r��*�(C�a�%���E0�)��I�@<�>&?����&�L��`��Zk�w�B���f��F|�^�D:S�:�(�z;<;���\�h~��x&����
ۡ^�x��.1Ź�"���V�)'�^��?���'/<ޭ�1�aJ�D��4TH�_�z��p�埽rea��j-���r�����W���L#�^٨�}^�Z
��z���՛�q���>*媖KE'w����נ@Ƹ+�+�R�~��K���$>_�X���0��4� ���զ�+ '|���8H��)�\T��*5�f�V�#(��1bK�5��C��q����ei)Tp�O"�@�c��ȩh�?q�;���E2���V���uWߨF��l���yFPܠk�)�A�h@��~F�\ P���žn��m_��j+�qE�2���y������U��q���`��\`�z�\h ��aҒ+�Oh���Z�7��T��*�M����g4�;Xl`=�@���B��N�5N��GhvnJ=��ѮO�5>�Z�֜�nȓp<�w���4u�\l΁�G��P\�y�3G�>ߌ�Q��e�Z�r\׭�$��h8c��Y!�Q2����
F������;M�9F\�hڗ��lM��٣�?��Y���Q�ZƠ��t����I���_my��,_���ME��?:��.����q,C��#����;O E���0��+H�azH�g�t��dT�^�U7^}���?�<u�9e���z��~:J��$Cq̠���?�~Ҳ��/}^���A8zR�M�Z�+0e��9M��Pe��	��n��3��XS����ڛ�U:Ōq>oM�c]|��V��c�v�����D��D0����3'�nՔJ"�$m߼^�_���߬��+�43��\�w{�Sv�m7!$u�y��6#��x�\����hi��#�ծ:p⤊՚���y
Ua�kBV;�R�M�+A&pT�B�&V�����SN���K����(�u�+�U���-rB:�	�A�Ŋ�I��j�s��=C:B5�|��L}ym߸A�Hۀ�2S�c#��Y��/�\�O���w6�S���̔`Z�Ϋ�pX+jo �e����y�bʔd�%?_;�h"g��H2���A%3Lq����3��P,y�ɋ|��{�s	�k�@@ָ��F ��+�¶5������겉B@��������׿wǳG�|�M��UA7L��A�x�����K���g]�w�������3:u� �0�Z�=L�
�o^"��@���(��*F¯2ꧻ
H�0~XC W�R�X&��q`&XS�$B 
����)��@7�b��1�eN�s�EE�)̀Ofl�B�uw�|������Hn$t �*�U��N�<�'�v:�0�`�Ԭ5�e�6���"͜�?7��e�J�i�� +���dRC#����\y&�d�L�K��)��DA+�%`��	gM��÷��l���rE��tw�I�d�t:��#s��X+��BA0n��x��2�̄u݁G�@����5-����M�I
��Q���=���h�h\�}c�X��/���k7��G@�s���ôb�A�fCו�u�E��6ݘ�����X!Fm��W�Z`52��4�$u�,G�@�m���Ixa��!�=m� � OY��Xc�$�N�cY�Ƙ�ǘ1$� ��Q�`���:(�����֑Çl*A��ؽF�5�����70��r��i�qzw=�}j���
�z蜬�P�]N0�b��8TM�.3ɘ�KV�Z1:����Jax���U�ݸ`4���v���h �L6�����<����]����fg�¾�:~zZ�vB�:S����U��nP��-�-6�
[
g�rX�F"�/.'HO�b���E8~���;j�[\j��e��#��@�h?���1
�)�Ru��W�ٙ�ŷ���>�t͕z�[�ä9�0X�E��d�-\D6]!W�tz��:��R-K�(��,i�$��B=��v�t��N���{m7VHF|v�x�<�Ri�O*�9�Z��	���}2c��œ�S`� �1}A�'��G)�T)�]耆����?�9�띜Ac�fm7V�:lVi�XO,LM��o�M�\{�֎�(֨���{�ȸ����in�!��(o�N
w$��Q�];��KKz`�za��g��`Jf{�&�0E��4*�����cRmzA�xD������j��C!FB��:?#�V�	�$���a
�ҝ�ᮄ{�FJ��{.��mb��[���S׎���,������3��D�+*e�*|ӕ���CѺ�K�/h��LOt�l~���ȝ�}��1�|$�x��l���્�+~:uƁ���E�F�*h9�S�A��U$��}�EhP�cl�!c�ɞV��5̡l�h(ۓ��;된��%Q� /
#�͹fO��b�m_�Jg4��KuF1�#��Z�8y�F� ZM����k||�������l������,/Ag�wuv��Q��3�@:���	�.F��/("x>�Ғ�=I����DA�<U����pxy�Ʌg8 
�}	ٍE�HK�e����y��,��Q���ւ�~߻�N�����O*�ـ�
9U+����u��Kڱ�9S��_�J-�q]xѕ��._�N��y5���$�1uح�􆎄����m�����i� ��咘'�8�F(J۾��"v��f�����H'Ҧ'��j��۩����P��%��V�@Р��:!h\,x��p�� �D�#L��@].����zq׎бw�!
h7��MʱV��? VO\�v�z0n�"�j(�˹�(..�=#�hL�eP�ժ�h�7�_��`o@r3�6>��]�t�� �L)Iy�C�~�خ��(�z�J���g���0�$�`Xd�6�&�m٩�Ϗ�bة#Al`>&��$�X](}��}}ށ>�裚���
��g�bz۶m�HFɐ�{e��o��ڇ����2�L�`11A�h�UJ��6�b�=�ۧ�\��F3��zz|&Xg2��$�n��]�^8��jf����K��#�t��I-,/�)����A|_ڊ�"~�1�3�#
k�t�5����ݳ��˄x�i��`~���8�e����q�}:"6F���9GG�D��8��5�8bC\GCT)/iÚ�ھq�~�]wj2+-��5�M�;�5B�ׂ�	�w�Ͷr�Ġfj�R;%����_=�C����i�9��<+�H"iV��%&��
��4�}v�d�0�����ryV������<����x`�0P��V2Tm����I���6���ѩ��_K��hq�������⦵#S�V������-;���d%�^Qa��Z����o7#ںi���љg����yYНN�>(i����]t.c+#�;��kG[�L��C���}���1�*�b�ƕA؀o�Y #����@��\�`Fǖ�x��Qx*)��h��Τ���hM��ۘ�#�qh�rxG�0�jB�����I9r@�j�����Ͽ�T҆M[5>�V�%KY��,��Tq��3g� �W542fkE��FۦX0be�dlM�0"��؝Cqk�S,-./Y��/^ʽ������~�p����+~��9X�̥��`#��A�\^�3sA��Q���DU��-_��]~ ��Eg�:�1{:��SGu��+ЬJ던
�m�r�2���N��6��x����S7m��9�X.���T]�tDD�xڡC���ZS�TU/�:<Z�����Ōh�cCx�\��X��������)��B1@��}D����h�Ր���J�]�K���t �3�3�&J�"h�2���A������}���KO��l���U��9�S��E���}S�St.�/wV.�4D<���e��_�{/�E@@qᄆ$NPu����bi	$��3X\�tB�$���a1K���y������X4c��
�hХ��?��<=�e���2Lnx��>X�0A�I�L���>��U=��c���q���ܤ`H�m���{��qk
D�~��9�����E�(��Ңi��=��LyPDC`��4�|*�u>� Ͱe��z�`|H7�օ1%C��u&�n̚r}j�"����{ݔ�)��h���lXǵToU�xݡ�Htɀo6��������ʝ�J�n04���N=����Uiv���xO!�d.�Ig2�C�5�� �IZ��Q0[p^
rT���c�,�ff��P.k��skU����.vh��{P�Fb����
	M�^P,�R-��R����}A/8��bM��� am`ݫ8��״�0�@��l�Tk&v��Cf���%�3\@w�#磋G���{����\5�^0!�{�T2�?HK��Xi�����r���\�jկ�C�ÿ��]��?�܎L���7z�͂���m��)�Ψ�X��0��e6���,*`��ʤ�Oa�'�t܋�;�nr�R��J� $��`I?��Պ��-'Q3
r���	y�#�H\A�^).{w�Tkhxl�t#�;E��R+'� (iz���0��
ϣR\�T`IY���l��@�ة{��6t��a{�:|�\�������\��{s)�u�͠j5�&�[�T֝b8���|�/���Ɲ�g=���5'!�4௳G#�x:�c�6���x*� �"P{J���k�}yDU��T�����nS9W���n��.��w�z �0	�?T� �����(�"�����޴�y�1͜>e�։t���Ƶ��M�L"����e�촅}L��޽�."�öڤ�$�\�P����Uݡ&t��Ǯ$x~��r2�F����E�(s�����+z&��{k�5yƞU&Q����,��#x��0*a��Hkq~�@+��
~ #	P�R��qf��ђM-p����� ��'ۯ��q�Z������][�
kꁶF%�(��9S�`Z�Jf��a��y#"$i���&�^,f��a��Te�+`Oa@4V.������fc�J �=�21�ٝ���e[�WfҔ����GI�+�&���;�
�ѹ�~?�z���[�.9u���s�L��g"�b�ʵmG�|!WP.�P��;���<�
�(^���H|�>���NBc�1��L�6��N�T@����{ ���Hx���5(�0��P�Ìh�(��Ҙ�s�n:�+�x(�cI�k5�&�O�:��]�\-g�W��He|�FG�ur�zz���r��93�x}�CJ��k|�Z�Y���>�� ����-0�s�e@/eE�
��`Q#�V�)M"n�?�/��#�b�`)MB���Ϟ�ɩ��8XE���x-�R�qv&���ye�;������ !f��(h��r/��L�p��c(��`ʽD2�-��ǻx~^�*b:����A��M���.&��cj�M�Co�?+m�ܛ���7m\y�����՗���g�?V�D��'����g��X��B�mڦz��p�2���A�N��+�͚Zez�d��6�^.>sǯ- Ż��J��؁2
J^4F��I�T�>���^��/)��7
�:<L]:�4���/���v��й����� ��h���M:|=T��ޙ0p�ЙϤb��$�����u��[l��
�*�Ֆ����m����+���[ޡ���}y�[���^}_��4�nb" sh��y�V�:�{�oѣ�׀�����\:c4�����;$i�:è�L�g��9��LR'��#��F 6=iY�(�k͞�M<���ES�̅bɀG�#�]�r��"�Aq�6;^�M�Ui��f�U���Y��������z���]���5�L;b<}zJKs^=�rY���0���g~�O�D���g��5�i�p��#�̄&}�{Z+48����z{{�Q�:P�#���>�K%%r}�Ǹûۚ���6�Q���2�</D[��O^B,	�E,
�>P�ZA���2v��|!L8�h7$u��!|�%�[��-�].W58�B��am�t�.� �Jyy�#f����05�&''�����F�°�;3x��>��� (�|BR0'Z�����	=�h*M�<0I.j���b�	(W(�ʦ�m�����z�����lZ�gN��P"���"�"�����B���"K� �r��)�ɸ��Zo��˳z��*��ڇ�?S3�D:���.��b�j%�x��V���D�=���왟�$���aQ�j��7��:�)]�D�3q�Gu�lIh�ag�A��2�W13R�J�~�덮�נ얛���FI�H�Vej�3j�)F?�p����r�4�^��kOn-�k��SNR��v�xF�V�TE,v������F'V��0
Db(��.
>�ȂP�@q䙍���N���1ϖ;GC�j�O=�d�W(���D֤f�t�{�G�w
8p[�1H��M FL1�9~��#��?��3�;��+H��썽JRx�9���c#]6��m8�j0�2�رc.
��>XX���4;;�^x!���I-����I�lj(]^?�����Wz��K�D���Q�j�o��u�V�Q���T��$�䊕���98&�7��F<��d&�b�
g:�B�\?�d\Y��"�Rh���Z���P��O�/}k��T:�c li��'g��C�_��������򡃖5�NG\cv~A۷o�Q /��wE��&V��K���uld�	�Q ���rM�d��!�'��Q�Ssyɂ��~�=�F�W�:�� )���v����.��jcj���š��[d��8��*�.��Qj �;]�ħH]Ǐ���*fh `�,����&����j��N����j�Y'M~�i��W*���1f���e߾}���_}��?Lrz47����pPK�y�O3�2ɶ�l\��^إo�I��e}�K_ե��dЈQ�u�ɃX�W!��]�;�����'G���)�`Sg4�cL��t�AD�i�{9�fR$,��(��h�?g����J#�GNu��dZ�8iD�����Ӫ�MN�����N��׫�����.=y���S'�nƆG�=:x�������	=�����W���`�:������������K�{���ګ���:��ӊ�M�a��s� `YX������l`$Ӟ�A/���c'�z��t앻�Į;����h}��O'�&�18[����I=�!/C�J�v�(oZD�ӦzK�t��I I褧#M���Nܧ�Ų�\�<�MF��x�KQ����s'�k��]Ъ5�tz��f��)����a-��ilh�b��ٸU����]ȓ���KnVo�Y	SV)##c��,����{���g�ǹ�Z�r���"\`���3�X���d��2��wŝ#�t�8��U���)�]  �4+�<L��v����T3�����܎x
 �ެ�#�N������C��/k��W�3�j�㊥{�e�J$�^Op����}��4.�cnbܧj`Y$bA�k��7l�PL�'wGM��a`a�C�y���`"�E���+�zi4��B��f�V�Z��G������@���ȍ�jtb\'�FD�    IDAT��P �Nk�r����4��$x�n�}�HҢ�I��U�&44<���S�r�����Ǒ��4��,o��­�_��_�C�����{^�Y�X5#q�6��%�Cg;I�^�0v��r�:uJ������=�I2i6=�dW]"�����#T�Xm�����EE���$^�y[6��I����:o��/���Ċ�L�9��iF8׮����������ץ�_���viמ�f�]p�Ez��gu��1݌Wq*e�$���E�ګ�����ƋY=���Y�ZS{^ڧ��l�O�Iŵ�cZ:{\c���|I�lt��lZ�6mW�w�`*.�z����D��g��a'80.������/C���n2�>�.H��ե�Pd���(�A�cV7nR,��c�?i9k����a�AQX7��~�J#�gNM������;��P���ˮ��O>��6:>������:~���
��[�j�K{4}fF�''�fr���>����L\���s���m^�~�mܰYW^u���_�y�\����:}�8��N��@ÝW�^*�+z�t�hZ[��:	�#BB��S���f��L�㣎�\����hݚ	͜���[#aqV;v��R���	Ɏr��J����K5P��SO>��l�.<�~�Yw�8����hǎ�����Z�ݻ��^mۺ�v���Li���V�ۼy�=�O��Ҏ���9^P��s�u��7��﷛�M7�Ng��T�F��{542�R�j�+�n�!��,�Ύ�"����9Ǌ7��	+P�b�\��J����-���T��T�}�F�ǿ�1�T��K)��
�T��sM���@�4�*θ�(���Q��%4�{����L/8$n���e��؄DT�RE�\��m�To,�˷k��=����߯�z���t�
��#��(�M:b�Ͻ���&��0����n��3�5J��}���UN�<��9 !u����1�f���Ȥ �8���i�@�4f�
�C���o'��*��re<�&��Eۚ����ϩ;j?�� 8�n7Cw���₋�x��-�'�<^�O(G1���nتB���>&L�(,�x��i V�fgq]{m��Y;�y�2*/̅�R-�vR�XV۫$���|�V����m�"� &$t�05f���\ß���o@��D09�T+�������%u���ۜ
������'��	n�d�;�׺���w�>��:�
�O�Z��ГѺ���҆�/�v��qÊc� y�y��v;������-}�����d�v��}syCB߾y������0F�耊QRw�@0d\^��$v�٠�6(�e�k:�.���ڂ餫2^U��J��B6����hphL/�?��v�������$��K/֮�3& ��Uk�httX;w��ƍ��:6����oՑ#G�w�^w��^}�v�����'�"7l�e���nW�KE0u-Ͻ���<�H���^�'c�ӑ�E��x�F'-��e'���1��g��;�0�s9h�s����O��5�w��LM?�D\�~�ͪ�漃���t���Ǖ���2�38;}Z�&�t��Ͷɬ-����%>���|�y�>��CA�V�UW]����;tn��F��s�>��e�X֪��u�eW���#ڽ�E�hU��N?�ᾜN>��w����ĳ��r��Z�z�f�.yO�u vd �}�ɋ ȑ�F|A�;��Bw�͏��U�s �;2�`1ZU�Y5��[7�7����x&&W�_�B�ʵ�z�F̓oיf�������q=��cbo	���k��9}��gt�u�ꩧ��VA�:�ַ�M�>��N�<�[n�������gm
=
�ի�j��-ڳ�%�XT'�ҙ�ǵjŰ�cY��g:l;���ç4�z���u��MM�9׍@/E_�eB��ߏ?̒z�+�؀!���68�"hD �%��㨫��ஒ�������,�dzꔖˌ�s^Y)�1�ծ+�hk| �v���Ц��k`x���|ȸ�L:���+�ʡ�j6�ڶ���[֡��Փ+x����Փz��u��)]~���?g�Nx��k���飪�f�q��zu߽���7ݢ��y��Y%�������Y��#�2#T
o&[LT��:tȝ�E]�8�.�Έ������~�A9���l��O�O��s\�z�}b����� lFNw�,�A����iI������L)����8����z�Y�s��l٣��Ii����df0*�U�֫�Z1֯�S�Luf�?�P��BM}��\�d��ZZ\6��&��������2rB�fϭ]4b�ݥ�u
P��� ��; 0&N�4 Rq��Kֆ�]�Ž�0K~���O�ï�*�l���k�A&/�;�?q���]��\��f�1;?#
���<.�6���dz�ڽw���@��0^K�bJE��-�]��_�Co�����˿���3���H�:	�~�Ahr��.�r�z���ג_�������C��t�`ai�㢆p��
_>�μ{�I�f �R�V����#�i��u:u�~T�.�X/�yI;^ܣ���0*v�Ht�UWh��O�� w���.����cOj���n�:=��3��H�Xc��klڰQ�ׯ�/��Pe3"�:e���׽Η���R)��%�M����fOTq�������R�/i��d��_���s�};�8�ݓs� .��e*��G=����b]ei�rQ&�2���.��lZ��K.��� f0�{b�L�o}���X�Kp�V�v1n�������	.628s�:{�P%��j�$Fȉ7�ώ�=�r#c�ZՄ��p2��m�l�|�C��"卓6����\恞2�cţ�N`iy�)�L��E�=���Ɔ0=1�g���>=;���~|��Ǌ<�T����<�_���pN���'ѯ��;[ے .N�S�y��l�N
��5x�,-<F�����|�]��iL�����ŉ���1k)K�͂���������߃��8%�$���ڍ��b.��Ő�P�L���\V���#T����/>G(ҍb݄R����P4t~bC����ސձ;�����/>1���s�X]�A����~�s�A�̜ѽ��7�y��sf������3u�Z�x�8I#tae�Ԯ�c�˥O*�;>���i!	�^ѷZ6�d�K_�	ܘ��ÂrO+��ǂ��'���e��R]K�9T���;�}(�)ctbrlT����I��O�<���*B�J3NJuM����~7Ν�����q�#L�����]<~�W.\@,�����	wrf.O��x�����>L���q�ŋz�'g�z���=d3T
�%�ez��pjb��8��Ý����n._�P�i��?G���DP�H�F�Ln�!�'D?�S3+�G��O;��[y��d�`���s�?��ŭk��!��Q���,Vװsp`Z��i�� ��Ƶk8:��7��ƻ�+�#J�g��tk^]^�����ȸ�/���Y�بi��\������=��I�,��͌�I��-v�P+�������G���7�)��6~G��K�b����A�p5cuc]���Ŷb��@��1��$a��c��<�8�z`��lz���V<��X;,H�1���4�e�d�Cmx��H����~)�/�<f��9�o���9�ŸkgXy]mO�*�$|;��芠\�c�ټ�}Z�2��^�tSa<���\��P���/��b2�u��Øп-�
���詳8I3x�����Sb����G�Y��1S���C���<�[d#ڐ\����'iNBx��QC���X'���P�$���clm��d�#�!�M~��r�ʤ�87=��g�p�HkH����e$��䍏O"��it�V��	����X�O�7��/���K�u�A�a{gO_<׋ew2K����X}�nS]ݤ�H�ۇY���.N]���#J}�����ƥ��A���d��H���5�J���z���v��}�N͐���x_X�|.���V�&Og���l`�ɠ%L	��������b�S��{�E"�966�������~��G*4l@~��baaAr)�Ft��M����5+�:���`y�*�7������W���Y�>�˔
�2�pH�4�A|5K>B�z'�$)t����ʗ�˄o?��m�u�����hR�h����Sc����ß=��a�(�t����%�q��v;��4b^;f�FE�"����!�6�4��y>5=��!M�<T_�|��pn=}�����x�zKO�k~��Lc}m���1?!�ugA�;[�Q�028��]j68<Q�M	
%S�FE���a;m�cWn�Y��!
&�̆��;-kT�y�ZREB�<�h�C[9,~NM�#��8y�t�DM!����-�$�9�����YEGď��|��_hB$�r�λ�:<��˯�����ocwgC�2��⇿��XY����Ο?+t�������x��(._����5$��^�g����=\8;�'��*`���ѯV�zG� z�r"If�Ţ�[>��0�0l��s8�Ε	C:�Z5C�I��n��-[Z���Pww,�k�`ce}]jP��>W�-��ͻ�S����o�@�� �{�1�G|OWV�pt���kW������rh��{�|Ag3��N��9������#��ӧ��۟���'�KG�*�#�1�|�X����ۉH� \��Nw��nMDj|F��O{�P�͆��-�Zoo�~���o���&�������G�����U0��b�D��h(1�9����P�!VKea��ljP����o���ɦ��o�{
E�r�����k￲.r'z���Y��UL��<�*���\+�o��j��^���e��O_���)?��W/�:'��O���\I�������-�N����&��RF%;xNJ��ܭ�E9�m�����~h�4���ً*R+/��N���| �pE��ՀS���8��C��54�f�
���
ֶ�d�J�I%��܌i%���(Cb� �n;A?��VDʢ��B.^Dgg7^/�`[D"C[ʗrrl\�<w3���ƹ����6��#	�%�v����[KO`.����v��c��m�FN�X3�6�����"�\�#Si,�F�ԊmCʭ��wV�ͥo�k,�\U�>�3=5��.?��#؝���6���	�/���Kx�)s�F'�4��ǔeLt�����}�;�!����k��ؠ|��t�.�����1�BN{X~7��-v��{߈���0����rr���e���qz�	u������u��TV�[[:Y2m��Ug*��%�{Ng��k'��2Ku�ʻ������z}ƙ����|zS3t��z9� �N��B��c�V���/?E��D��E�Y>���!:�v�3Diܘ9sF�?��_?0�L`f��-j�W���
�b ]=F��k����� �J�FM+��Yk�g��gP*ftP'Ѵ��7|
]}���eg�Cz{��t_�7�x2�f��oH�F�9J�h:�.�bMӜGV�TV���*�i�ݪ���Cwַ����'2�X��ӹ� 29C;�8>č�gq�����Z�ޓŁ.hl�/��řS�x��c ���i<�{�Ã8N�>���^<���t*)5��Q��}����x4���K�q���f5�Z!+�q�M��X?|�(6".Ur0��"ֆdu1�����S�w$"R���Z�Ri�[����Y��kxI���v��YM��#�`�=�I�(n�\	���٨����H'���<:"a�?�^�|����b�J�u���MO�
-�����۷�s����_�*����7޺�����s�����za�M�V�oo(��	�7���i��n�A�\)!1��񾑱��,�R�}�vD�o7��dn�I$��B�����8`#����#� %�+��q�B�x���\���o�F!5h`vfZ�ܣ����i�z�������K��ӳ3jLH�	�d�B��8�<Z�S=����w�>J9C5P����׉B����j���p����(�5���'�_,���o�:x�H��y�\̬ԝ��w:pv���:r'F���t~T��mE�	=Fg%�G���J�P9�
>7��6�K,�2�ܒ8�q�r	~���n��(��v����`NЀ�Z� ��VSv�0=1/��lf��	ary���,A2/K
��u����<��!�R�HKUB(�1+�\�U�a^/3�	�V������R*�^�!���������{�,2Ŗ�H�0�[�$�,%����T�Zz\iˍ�^�*-�@�W�?z�%�0�sM;�Q�P����=t�����^.���0y�����b6�j���F:L��CWwL2����z�(�yB���;��zoo_ ��P ���a�Ãu��BeJ�QJEC� +J�X|���
ɸ��'�Rӊ+�� Vg@iG$j�d�J�sjjO�d�K]�4?Z
[�W�!��T@!E�3��u�E���X�<�V3�"�bL��鴡imh�?8����s���]9QmrK׸���}v�9=*��H�����Gs�f
��o߾�L��/^�!!A�(���ҊlD�hUE��Ή���+F�&=�SN!��!R�[��Z��\Ewg�'�!�L��G�n�d�wT�X���Ъ�l����̆��fG�Gߏ�<�GN���V��	M� ���j� U��>tvD���E�ؑ�5M�P��Գ�0��kQͣ'�õ�gP����@�i��'��͌��n��t�s����sI�Nrl<lx��[j*�VWtVPC~W/���s�5,±��._<��YD�H�+����4���;C��'�fO���q���=��H�S*�����EI��VL(��v�mPP�sQ����h9���f�Gz�wؑˤ�0+�+�L���<IzY���(�G����.ɣ25L&<~�����5�~�g'x����Q�y����I���b�e�� n�|_=|�cB��4+X}���6\(�xW�@�aF�g�Sg�u^�;~�6W�}^	ml96��r��1���l��0�vke�O;��j�p�[$�3�"ܸ~�r^�qks�=}X�9����u��̗�J�Fǆ��ۃ��~���/�xGGƄ:�d�:�׌����������ʿg1�����T*�X�C$d6^s��Aux�E���X]_QDh����T̲�b�׬�';"���޺��n��<�f��?����������P�M�_�����IA���y��dҹV&�a�t+�<��J�sj�q��g���&#&���o���e��))�jtN4W����nC�l�B�w�H�I��X����s��|�7ܺz�lB/*����(r��N�9�ٯ�l���-;�Hn�� N����khdP/,�uh��Pr�*� �X]���s0Ӡ��C(���Pw�����A�d�;"����m��3ӝ�j+��-�QT EW�A8�NQ�z�u混���!�~���N�˕Q�6�H籵w�kg�$	"نR��LZ�w~�!*��|Q�6ܻW2�4O`C4���آ|9nݺ-	;~�z�d�S�E����X�d��0vU��5�MXL%,?����&
�#�X�D����w>��Tu�=o�^�i�J��ei���Ǭ�������ª���:#��V~��D+>���Y����EP�Q�\4*�ug��'���"��KY�<
ýH�UL���w�p뺍�#�I�C@�{��7o�o��cCcL�R�JV4!� $������0���p$�|���K��`�5l��`��\	fW�����i��ly�;�i^�!RV=Fz�S��/�{{�F3�I�S ���ìz�ȓň�/]�dLزR��唜�B�M+���Rl�ߪ��I�W7�wL��#���
̵�>�X��H�h�Vװ��Ղ}!�1���b�����%`��p�͠�'���Qtv��sPjiu8q��C�����K���8���4�7�yI�z{F��F00y&�9��0�T���~���PCK�[����Z���o@�<A��n��T�1Q:IG���{�^��� :�!��no�bim��ݯ    IDAT�&����}:Mje�j%L���3��>ϝ�}$R�I���zE���g'��DRZ�?�+׮k��I�SW,�ۅ��=�^�E�M$ɐ�"V^=Fr�f	��E�j@�}���nm#,^�g"amΏ�y�s�i�JS(��j��p5#)��<�*��7�I�
C]��0�R(�'��� ��}�i����ڣWEm�Yᮊp$���Aeq����̬P\*�8��z��~N2��_�)����
Q�=sF*u�ŉ^�,�t�� >��]��ˊpԏ�b�˯�Aϖ
pѰ���z����E��ߺ��� .@ѿWA_n6?��?��k���k �Hȝp�lf�
��aǹً*詤A�o?��	[��Ҡ��m9��Ii�AAo(>4��܃v�{����5x��:"!I���L����v����jz�!N�!¦��8=>3��.'��V�wp(x��T_� ��)�c�l����'����'48c�b�������g�Uh,�Nv��9X8M�sG|(Tj(4��p����)���W�p�j��ѵ��q{��!,�0C3��~�/]�� �e�IH�jZP6����J���5���H��p�Ú���̥V�����(�^�vÄ��޻�N�5�MN��7�͒�X�$"ѣ@(����]�)���/����&�
:P�Q�Cj��Xzv��m��D�+���ޅ�Gw���m�� ��mm4�m��6D�.��>�Q#ɩ����g@x~�[;hI�l(��K�bK�e���A�Vݤ�5���� 8�ǂ	d�-N�u�embO/�fv�uHR;��?��Dx�+M4�ɯ>7,a����R(��~�p ���ȍ�?��n���"v�[��RG$Bo�:���Ff�	�k���	��Kr33&�o[[�C����4�D1(��XI6�b�xW��ZSS��9í�Q-)2t���HXS'�>�+���o������@er[qvbPzt*b�=���oT����0}z�A/v67O�=���k�p�ƺ�̀�V�F &ē	��[w9�����G��xt�W@5�2ar:���0u�,n?j��G:�1���gS�i�l4��������n4=�H�`Y���3�����N�4��جp;,���E�'B��g@d�0u�L���H�Nt\�WTЋ�$Fz������\^dAQZ�����Dh�	t����95�����abtB?#��Ã�)�ml!����$ӛZ���`k	�jɣ}�Gl^C�c����`g�Є6z�{/��<5_xc�h��8j���Cw���G�Aə�Z��΁V~y��G��AO4��hX��n������Q�)�|l��=�&=A�:5)t������e6"S�B*Iv�57�r�~�+�;b�����=��'��1�^W��f�Y�*�!_Y,����u#��b�&�ULw��������ܹ��U��6����������k"�.�|@�Z�v^�M=���)��C�(����c�Y��i<��l���w#�F��S5�i(`�R���c�x�v��F������~_8*�P�nF06X�*Ο�D1�@�x��(��N�!-..#��W��px׃�ɓ���iD!o@༙�Pϝ3:0t=�����P��`��}��K��*�Ŧo��}��,����L��f�/@[On/H&a��mAW
�c�>�t"N�x#U�����x��9}��/V�����k��TuH����A?�[���ȕ��0��'�~��Hvq{�o�	~��ߗ����̃����������MK�)��io�YMc��Hn����2���\{v_�BM��f����;�H6F�6&G����=	�:[�RN�l�H�!��`��)o�猝�F	��T8�JX�(�jx0�[{i�LNɮ�-P)��,���Sp[ G���� �z{�w@H�����d��=��I�]i��tx%G��f�I���ŋ��\_^�u�T�f�?c$����֗#��V#��S��C��x"�r6B|�r{wh<o���*B��`!W�-�6̌�k�v��ƨ�=�jW0��)t��yJD�8��b�V�j�p{�� 6����J�4:�N���[��*��G;c��G�HJņ���$r�#�nm��+�����\���&��r��Ш(�9`��9�^Z���1�� �5��Y�n|��_�e��V<�iS$ڇ�1L_��x���T�G&K\����Y�a���M����C穬�������V�;/����T�B�ac���ų��E�(�2BD��"��^E�ʠLvw 0�0�KRV����6��bBV�<�jT��a�f�t��I���_~%q*#r�2���03&�RP���O�x��P
Kmy[�/���1L�rٸ���r��1��^F �+U?�kֶ�n{D&�КxX,��^|N��`v�,,�D˗�=���.Y;^��2��!�t���h6U�;<���M�m�1R��t��a��W#z��r%�w�g0����E�'���������Hk^��ilΉ�q-æ������sUɷ-�:ba��������F:2�Nzf�ݬ�'b�?��ε���� ���������r��*�4�]9�2��^��cu�¹�8ɕ�NQ�mڕ����`����.���c����n��UH[�c�P�c���aGgG�}��'�z�5B3v��n<y�
�/`rz�4;5	��Ts�qi�4������8�I�uQjF]���Y�䄥X���eG�}Y�gj3��13��3�.�u���r	l/ϫ�[�w^�!�#_��7.����5)�I��7�]�D�(����·�}�ߐ	�8��N��(��H��v| ��:���N�����7y��V��^�ӗKh�p�E�#щ*u�7/�G�������G
 Q�i�� ����ǝ�]���k�6�h���j�1����_���^��:�T�ql�|����)�%i�|��:p��mtB�ljި%Zp�b[\���d�q���hIq%����Z�IJC�/;caM�\Ӹ(c��)�=�S+�B��WK��;ʡܴ�Դ���6d���@�딿 #]�v��L�Z�,�nt�t)p�S:�%9E�"��55�w	�m��>Ie��G���;�6_a{�9
�m8�5�[H5�;08y��!0��-�1��F�?d���F��H-#�R����d�(�+[�2D<���q=�R'�I���|�Z�S�@_��p0*v���:v��ȔDB�IiW�^[A����w����I��֖�p��9vw �<BG$�"�)��?��T��d���ƕ�����X_ߔ��iD�R��>�Ń����YԄK����{p��H���N���q ���a�o��:�j9�����g��H�x��u8��}0�
>#,(Z�СSo,�5��Vd��p�������Z�L�2��[]�IvsA7n\>��� N����;��nŭ�7��L%�vۅ�M�����+�,:A���F��"!?FG�t�T@��]��jI���+x���*�����(T�P��f.��чMfê��s� �F,�^��>�P�"�ÜG9�v��Na�s���N"k	A���1�P�3<.�
���!�Z����{�g�P>�1�����a�n��נBga�zz���Xd.����P����,T�ߓ�6#:x�y��3B~u�̣ !��0��+��I�+(��>�5O��&t��F%7���o�}��WA�N���?����~���`��M�p���Muc���q��t���:�6��S�:}+�$��&j�m��_MI���S!J�
xog����|��e���&.�����6�b�+D�Ꮅ���`�;,8��D4�D��ĝ;�����_I�/�D�Ϳ���8���#'�����=�XF�$���A�%Ə4�Z��xObg��1,�"�J�|*��W��!�=c(�����y��(̗F>u��P"�	������O��ѼՊQ5�zC�H}=1���!f��H^�Ϸ�T��bB*S�'���.��^��֚��4,����Z-��M���ɴ�s�ړ�#9��7N9Z;�t������d���N�j�3�@���E� ܃[�U�J	�<���޺�_�-�B�;1u��
z�L�ծnY1�*:��Ŏ��Um#�� R0��A�����+4-���P�&�4��(O�^+������\(W4��?}�̓�Hq������
|�*��4\V��Qf�]@"]��GsrBd1��,�uǴ�#�����jJ"�ag�H+�U��<N���6w���U���߅��%l,�#�����
����w���ju� �I�6��pŽ(&�Q5$����;L�;u�ĬF��F	k�id&������¡�]yV�Q�[,2`Ȏ��KX�9@�p{�*�	�.N6�{��qp|����8fsm׮\��?�E&����G�P�A2�f�\Cd��&0�V��^2�DF�	n�G:	S43z�p��1P)p��Ï��)���ǨX�8�!J>*r��Y�5I�S��2q6Z\�6��N�j#IB&H�bSDo�V*_
���z�jcg��	�����P�ӗ+"�R�Q7��K�즆�xm�����ry��<y�[�{�}���rȳCԍ:�?�G"�����{�驩1����O?j9���O���׆���x|�3X�9���P�YT�G�/"�9���-yY�i׋6��}�8��k��,��7��ƪ�MA��j�+)q�Nm�oG�W�Bn�	�œ4
��5$���Ϥ-*�qйx��� (���$K��G�d�İ���?t�$g�Y|�����֒�{'�)E����H:�[��ܬaa��ڊ�G�!ɷ�bA���߾v�'��X���I����������/�,.��{Y)�����نK���0����8S/}k�N�e�Z@Y���=���m�r�wX���,H�2�Μ©�Q����VʣYe��!3jt���dӤ���.>}��խ�n�z���q�y���`r�^�<�7�D�!)�ӵ?�����Ә����!L��z�V:=u��qloo�`D�	�^��.�E���JUT->\��t��j2�v�����nc�R�Ӛ���y���5���!f1�D�&��Nc��K0'& Z�AD���BJ{u��� ���p�jV�a8��k�`�[+�ij`|�!F��]�=[�;�Ǔ���k����0"�y;�?��ˇ�R6C�c���E�pO+����9�m���f�T����£/��Y��R0��QX����ސ|ܙ���h�vi'�����]ħ���Ҫ�ԅ&$����Ѥc��/�EOw����P"����}�9�ސ�/�AÊO�����l?�sj�2I����c�}�:]r���I����vhJS�D���Q��yuu�>�t��{� W>m��+�X$"�{sO]�O��@�pKϿA1e@�|��v/̞�N_����g�ϒ�z�Z��	#<GM�M�J2Hnt��N�j"�j��g����p @ii,*�t$��mG�ZD�����lV�W,�g/_��W(��+�˫�^���Zc�1D�=���\�����N�%�v�pz|D6�$I�����jZ���C"��A�L"5Q�χ���*ܡ����B�.�0k�7�������fs#[m�G!s�9Y��}WK��8�z
��k���ӍU��G��D=Hh6�bH�y�v:�y���<p�V�A�q�&3%|3���
53�N��C�_O#�ވ_z1���rkkW��뻇H�9c_��ę�@d�ɜ�=�����V�X8D#~<�H�b��C��j�(߃��O���'p5H.ʅ�=@R��E�{G`uzu_h�Ky{���1o��:�x���F3ujգ0�7��<�l��bԛkU8��MD�X�w$��\��U]�(&���뤧��}]���b��Ǐ%��{984���^�˭�ߋg��{����t����!��w~�w�'"�����a�����c��_|�P��ɉ��VA�8-p�+���ȟ������
��q����O��D���e��Qo2ЀTגA�P�-�4Yq��UďNT��v�<�f't�ktIoZ�����"�8+q̝%LF1bQo�$��95�<侮��m��[b�nolJ�p��#d�V���1�_��D�U�d�O8��L���{[��r��N��%ϒ�r,����SII���a�-_�tV)#��z�2:���\��8{���u�,�KZ���a�Z~$�;Iq���A/r��
���~�@簠2�����"E42�x;C^Ik�lAu����R�LJ���:���`j|Dp'�����eӂ!�=�G����	�QA��V����s8}!Л��
N�ǭi���n�Q�#~��t"	ꓳ$����S�%�'f*Y����2�mլ�L��E����C��K�_�;�)�@ H���^<�����e5U�p̾(����'����++��}[���m����Fa�r5d�2� �C�Q���N�ܺ�:h�I����6R�$�v�Ս�C��$��c�0��Q�h�(���a��9��%��px���~�SS���W��Zu��K�ˊۥ�͚D�kyNsb��I�9�_|��B_D>u���^y���⛂N�#�7���k*�ټ1q{�����vtg䯱a�)���/�ր�A�\C
�w",��J��	���	�|���N`1�9"YT)����]M��VQ�It|o��F��/#�j��=7+�]����3,,,� vF�pXMRt� Wn�p��0�ץ�Μj��R�Z���ԉ��I��ww��>y����?�����g�:��0s�-M6�F�9Qb^�!�Qa�8�ƛ�{����p�%ɘY6T���&\v�B�������d�K�ר��>I>�z4ة6lx���OJ�U7,��6��{bn�Ѭ�3��eA8闞������@_�SL�YD y���'�0*�
���f9��lM���� �d�!��%�],>{���n�E�c���k#�/ �?�'����Y�˾M��&S/�^l6ݓ慠�\j:oA�$g�X�"=����R)��C����:�&	�M���71�����bd�(��W�(s�n5���J�{��RFc�#�
6"��$9�V��ښ�¬w<�E���j��P���9���$�EH(�ō+��/?ǹ3��e�=E�aS�*-�]�jn�#�g�y�������r�l'��'�����x���B�io��O��^a:NUD3J*�&.���㣌��$�]%���b��+_t%�٨�����"�-��5��f��9U�0��sB����i�.^�x�ˎݭmA�$԰�������W�����wQiZS�=9b�B^�ۧF�������M��%�Xxax���ɂ}|��Wų�2|wm�r�"b]�Ȥ�j���h�x�^^����R�j��������cXWNJ5ԬA\��t�\3:xZ��g�_�@�+�z>0��ǲm�9<���e��i@O���C�:���HÜbBx�C��)�385:��It�(�tqm�_.�ğ��� #S\�=�b��-���Ȱ�V�d
[�8��jw�̹�`R��X���|�D�ޔ�MM�����0#�̉O>06�GO���Ҧ:e�Z!��g_�`����a���������ac����M*=T>.�55��tKZf�*�)��aj�"$Ǳ���P620��0�w��8<�}&�9�����h8*ȑ(��_=۸�4�i^
�g��u��B�33��]�5YY���|dl���?<D0RJKVt���.c``H��SD����1)����+i�Yc,�*v7_c{�
�-!"��O�O�{�k'E�#��B6���ioe&p�]�I��<���U7�;��@9���w�ܣ*���Usg99<�Y6�N{kL�7Y�%A��)��**�@��/W��f�q��?�LM��M\����i�Nrkw=�8���=�Oʈ��ݡ5�]֯�p�\ٓ�.���`�,�Nn�u�^I�������^>�B��M�ݫ����/�zO��}�Q�&ţ���)cTEV%�]�}t�4����Wk�Z	f�A\�y�g�Ҩ���k��Q��_�&    IDATI!�F�Q�ʜ���Q�CB�;×��c� ���T7��J�X����+������0�	Y<�nl�N��@(�H���Pѹ�О�m~:"ď�z��~8�G�c8�x]f��������(�T�������IL���h�`w�B�`���Q����N�n��9��|"(TR(���d�Y�sOĭn��#C�8����D�j��XS����
�3Z1V�f�&0z��*[�֌tcrlX��|�J;{He���Z�%�7�$�>�U��p����� ج�a3OVg��F�T�i�?6܇gO�p��5��n��Nj6�֥NTrc��?�����{��|�����?��?J��NN�M|�aiJ�)��Z�o������e� �f�'��DQ�Yl�����Y��D��i�6�S�g$ǵW��N���t��vv77T�y�x3B��L*F{{u�,�`s��^)$Cv��"?����835�ŗ��G�d+�Q�����[q�}�M���o���Hܛ�؀�(�O�<.7r�v�,~yjN'(RnF�W)����Xy�͛�N�/S���_��C�{�QP�D�4MݰY�arrL��g�qNLL!�����:<n��{��0[�Ʉ�:�<ҩcَ�r�I�@o�֦�`#'�l6wt8Ǔ0[9Ҝ�*�po�:��(�?ҟC��/>�%�GG���/�&��WVp��)|��H&�111���>�y4
B�ꨰ��a��q!H��BO��9��_���N�	���@.�z_��\<h���D����Nܾy�s��H���/��X�å�4��*�2�M�}�.}�r>'�7:LQ�C�@�G�C~5Zl��n�dO'�:>����;Ϊ�$�>x�ޯ]� x�_/`sc?�������������:{��KS�[�o�/~�Dt���O
�g��S4�����Hf+����Y_����(�w4!�9�,�����F�+��Q�hG�V�f���y;�3FrVX�ܒ̑O�i�if��;��cmQS$�,O�ZWϞŵKcHy켞��!��X�Z��Ԥ���7�gO_��Z�M*Z�桭z	a��?�Wq�H�rj.��*�� zz;�7����Y��\��.d2I��u���4�[g���0^��� n��qՒ:�Ƴ{�����T&��(�]�S�|�=9��T���dC��Y�c�T�I��3W$u�Vc��BB�,b�|"O�T��k�1��-�N����{�JE|��)B� fOO����	�Ͽ���1�\��H�2��%�͌߿#d���s�l�ɩ��<!g�ݝ:g��D�$�1��LA��D��A����h=����de\e�����s_�Vˋ�FH6S�<{��A��k�hq��5�ό!�������0섵�hG�j`a�J�u�6`|lAbѐ�����T)Tx	�Aqx�X���Qd�=ձ���ۚ��LjL�?N�L�����!^�\V�Zw�	�ԗ��>ӛ}usK�4�?�x�l��p`%і������0���ˍH�#�⽝5LN�a}{_�ϣ��j���2
�hg�w�����~��|��3~��{Ɂ�/��?J�,�Y��^G�\n:�����t���q�mlo+ŉ�S!3g��×l���|^$���\�i�/?�B������p7�\,��P-����uw���Ȉf��Λ��#Oܢ&�rx����K�����$��<��%�uubj|LG�\Ѥ0s�,6������]$u��v�1 (;��o�	�q�����_
��e�(�s�Q�A�	"�������R,�R�j_�-:z�k5E�4�j�`�:B�|�v67$'ʥs853+����}�\tS|jK�.Χ�ul��	�09QLͲ�űh�&Lf����Lн�oЍ_~>���-4,F!E�y������gd���G�-f���<y�����r��	2y(�Hϛ7�+j6��ޥC�r/8�?��]0S�cj��Bo�B�Le<���8�y���]��UA�p�ք�h�S�TA�\�a8:<���ט����:�{E�{�`�j�� :P�+�Ӭ��K��U�	�du+���c�Q`���m�I�8����u$�e��"ƽ7ݬ���5�������	F���O^�u������JgU����{߿�@��؄��>�n�(�zxxP���D�zSh=�����^��)�Ն�MAt�	)B�,aN���5I<^�v���CHݽ}����;��%W��	�t���m2������V����v�LJ��L<��\
�Q����gc�p���zM�B�\�0%ӫ�밡3��@4���O��������~u�/^��p?�����E��U,x4���qLL����0[X�ZY��IԐ�2����9�!�w�U�Qɡ�M�����	�"�,��R^+�!L�)x��V*R)��=���w��XM�.z��,�G�Ь5������]�I��쉞�����yvx#���<vR�1~�F�q�~�33=:�l��t\���`�D����TZg
��G__��k+�D�J��F6WF_��X�l�N2)8f�VI�z���c�p�r[���Ϙ.Y���I���w��RAw���1C�'>�9-±�I6ID�ZkZCn�d8���t�h�f
4�!?�_�'��GY�Ӓ�����(�.Vk�犘{���L#=�(����_M�c旧3y�l�!��K�ʡ�|���	�y���upo��o���m��I�L
=���jyI��d�߸z	����1���b"Zj5�3O������n����*蟬�����?ʔm�Yn�V(���{�bIp��������i�8	���t8�H̤��̞����Y��<����݇FN:=8L�eF�.�b�R��*��f��,��p�oV	����"��7J%�F�9:D:_���!��&
ƶ�?:Ӟ^O+\$�x�}�8��%���<4:f�p�������+Pۮ��nss?�+W��Hf�����,S��Yl�����DTRW(A�&!�ț�΀ �78�z�.�����z}u�ߺ�J��WK����GOp"箆Lsdq���v�(脟:B~�QD�^��,u#��)��"lT�X��Q����/��U,U5��P!O ���#����vbc}��]��O���#���f��ʕ�XZZ�ÇE~!�<(Ǜ�Ot��z��SI��'x���ٍ�I	�:��v�}���tA���~�ƻ����	=���K8�V�h�{�92҅O>��}m8ó�%��>�u�T���A�%�a&s�N�cx�_�44����C����[�Q@i##"�j4�N�(\�PY���Uw,��fOO��Wb��������C_?fϝ�*=��b�]8�?Դ©��KȧsX^\[w�LUmT�����{p{}t��Y���6��jBwFS�^�� �N:��n�bȣ���u��U�sY��x�^�r+k�^B V4%Y���R�G'2�lH.�[AC�Z1�g���K!����V �[$�U�&y��x��B�^�6���o�d���(�zz��F��/?��ߺ-���7p��Y�����@�X��sx���|aQ�I��q����6��+�*�� J��X�5>�E��(���z�K3�h���_��.�{��e{�$W�Ȝ쓉�Yh�IR-W"n�_��_��ɴ�ʂ�ZX��l�$�+'����ֺr�ˆ|&-�$WV�O��ĔY�ۯ����@�6�M�B	m0����^�	4+���w��Ɠ|������X
����sp!ʳf����]���(
�"hRxa��������%]eA��p��S���S�LجN)��Gf�Cu����,x�hGe��ߣB�9IKN�v���e�Z���`�s�s�6�u]+B�t�d�,�r)/ΤӲ��ŊgK���@M}<�*|o9��������p� ;{�*�̹h���a���7X���j,��J��皐;W���6ӵ�AEY�Y�H�K�:�٠�tE��A6s���l2��3��Ŧ��,����Ox��~0:����v}��7��dʶ�0�t����kR�nG�Dou�m��G��Vq����Ӏ���j��u(������Y/�Oh�&;�N�o?�2�	�p���G������=v�bLg������>�JK����(��y<�.���V�ɡ,��1'0B��˒���^Y[�~��U8j���K�����KO���o������k�q���T"��3������=�R*�7P��ϱ���tZ�`$�"�bO���<A:'�����'cth�?�ѻȤr*��1�ۛ��¢�!Xp���|�gH5D_�~����$����[)�I���A�v��s�ml`� �?$X����ӯ��{q;6sdb2ئ+V@!<�!��O*����˗�h���?�5��ۉ��ettD��88�ë�/��[�T�c�`S�Ӹ����S��9�׊)<��78�}P�dsrw{5���A��b�M�J����҅s2��~�+�ׅ�E����B;P��}b�
�3s#ZSAw�=�N#H��pP�;U�<��%ە�d�^G*[�Sw�f����� �q�I���Y)���pjj�|��Ϝ�A"���#̞%��)�+���_-b��,��{�����u���+tuu�����_��ܼ}���KyBWj<܀��o
:�ڄ���
:��Z�y1����S�j����\pZ���pO��l맹o�G<E,S�[FO(�ӉSc�B�(S_�ʩ�)�}#��iI&�7���GI��63��J (�֥+��Y|�e�*v�vd,C���c��C$���!�?|�?���"�:eR	5)����D��;a��i�����^����ͪ�jrr�t�}��{Jp���a��!�un;L���{}~�b��
��s�Ɣ�M���.�k����3 _3z;����e�������y3������m�I�T�ȳ��^`zb#�]*l\{1����K���o����������5���ܹ��?�TH,Ld|�E�����Y���0R���	)A��'����
���PA������:����7rQ��R�{P*3���Ӯ�mz��6�m���s{n4U�P:7�׋��fp�b��	�2�֗q�N!�g�w)���i�:N���{5-�!7���:}K^��Gow��26h�b�_-���v�(�͕066!���E�1�?������=Z�l��<S~����V�D��F:<����&r�4B�1�Hr��(��F%?��?�}�'l�G!w����'U���;7.cvp��	��=8�(���}��8Je�eL}�_�}��,&�����B�����<����-��w���9E�k���S�ܵ�;ܓ�	w�4�WG͂�4�AG�4v��K���$���s�O!���1�ۋ��Y���}�h^�><i���Nh��-���ݼyS7�/��/E�D����~�?���*����C�fq�Q�b���_}�*�R�2�� �<@�ݚ�}���?���|0YX�����eG$ܡÞ�h�|��&N�ǯn��]�	����ō*.�N+���4�=�d���Pk���4�{��a<#��?�'�O�@��?����:#a]s�W���L���K�R��="�ϟbbl3�O���'b�߾}s��`sw����	�66���2�.?"��]���q�����[�1xB}*�VW��4��`g6�pr�F� �'���6<:��T
K�[���N�R�ڤ?<��RV�L.�Ya �]ݨ�xx���
gϟ$΂NB���;ҹ�-,� �A���bR-ᴙ%�t�Lx2w�C����g�hpjfZlޯ����s87{F��=$��o���ҿ�������=ّ޽���z�<x�L��������'"ŕi,C�B�&����	��$9$NƢ�s�-��q�����OEpd�9v�[:�J���#�É�ZA������۰�#V;��[N7�ֺ�#/U�l�d�BSn� _.	A�}pS>�#����R�Hbѯ�*(�s�|���\��aX�nēY+q��$��6���������Q�?}��xR������"���RV�h��*�n��b�j	��q��1�ҋ�T�.��z�d���k�� O��V���L�^�YP19t#<=9*�1%j|���Q�`��>�/a'���QB9�l��J�<C�:;���vj핈�01u
_߽�0���~ĺ��f!�T���Ww����{�b�I%a5����Zaqe�| ��U��r��K4ƄNz�l���9�>�`l �O�FG�UM]���!S�%���4<�>���=�GLwRڹb$4O�X�nѐO��J"<�b^��H0��?�u���X�/ ׿O���t���60�GU��8-�rv��K���X ��Gs��?�T��pKKK�˥���5����e�����h��� ��b�RS�U�����X^Z@6��'��~��M�(8��m��+��X���;����*�ml�������&��Tʢ��� ���µz�W^6�!S0���p�`���b̃,u|(���Ex�It�<�<Xd��%��m�p1Y�dU����/�x���5��N��Դ��c�.�GjM��Bt�{��X01�%����u� �_����U�/-� ����c{����/02>�ٙ32����S�:<҇��,�z-صk�����T��=�K126�gx��J]9w���v��p}��#zl��I�lktw�Wf,���HҲ��(�2*0�<ٕS�19u�\K���~��n�}�@"Yѷ�{_g�ݹ����_}����cr|B�:p�rx�j����[;0�]2�ZF6������Y�-�V�E�hhlP��/�&OM�Z<y�T�ɛo�FoW_|� O��[71:<�'�s�d���<�^�ϝ���.��P����Q:9)�xI�/'ttB���(*&���D%�Ģ+^&q$����B��Z^������r�Q��������)��V��7�\�@O7�w6q﫯Ő~��;��ٌ�lǢ��T����s�?J�\�F�Xk��ŏ02ث��=�(�,�q�-�����]5�.�G�#�B�A�4�I�'�&q���'���/�����3�<7�{+眫���sLCr��5��׀���k�ba��M��d�I����3�G��M6;�ʹ+�U�n�a����f�F�����]]���{��9�	?�/N��c�;���ʪ�����][�������^�н����+;t�y�p�ƕ]���N%�U�;l����^
���s����I�K��"6Ni&��������(������v6R��i�k"��H�cb���ݐ
!)h�i6����hO��n5�O_����ު*���������6w_��g�&��������bzz�xwn����.���p��;Xz���N���doS�>G&TA�
)o�k��N$�DX"��TL���9ׯ�G!�BSC=�ff��JajnA�*�fY �w!�>�.JB)���r���j^r��[jq� ��*��
��l���4G��@���6/�ԏ���[U��I���P�´���Z���S����+���$��
G�@/�g2rѣ̍�����
�b!�h"�3����� ��f�c��= 6��E���×�5|N���{KQ,P��k��:���-'F��D���4������w$��㶩c/�v��PDR"�d"*u
�	\N���d�����U�������1���ՠ���:�j��)�����ń�������_u&��5,��ɧ�1�4���k^zoY���a��+AĐߣ���)�������>=B8z��s��C�XZ2v�<6<�tr���O~t�������?��_��ɼ�Â�l�Q�����$�|�Ｋ���$�G�a�8��pJ�J���"���cQΥ3���|��;Ex99��]�G�1[�݂~~tg�z�����o�=T�c�;��|�����W����u���1�UU�&\��u�Y�" ��=X]^�A"ᇇ���<0���~��g��+���4�    IDAT���x���r�OD135��s|�<�v0�������*�ౕ0��Sm�#yt����N[P�˷?���JM,e�'}��
AaW���"p�����<��#���xe:gQ�킞��!�bMFN���=�q\�zE�JB~o@lOB�����;O����ɋ�E���h*����'�������� �#Oh���֩NILOO��;4��O�u�o]��6�V��{�������!y.f(�#�����n2e�@�ޚ�7�+��F`!gbu��l��Lv��z��������J�U��f1�Hf�ߥ��K�gE��3�jŰ�܄E-����`Ƶ ;@ĿɊ�|�5�N�zv<7����BWL���Q����f%3�$I�ɲWت��w8$Q�C �>���ˊ
�pk}�.]��e�����q�8���2�Qf��X�:A�u�b��]�)�#ɩ��?���eH�iG����ו���	!m���հ��������L�![�
�X]�����z��ө��dc��Y&2l�������P��u�9�e͂��1�Z�0ε��g�ξ���+^LϪ�p~\S���4�;:��7�̓Ͽ��h��-=;����Oq��E��>�y�׮�����)��zl
�x�9r�X�4���r�p����`��)D\:�$����Ѣ����[����z������&� ���V></*H\/�s�qO�y:�W/���U![��c$����N��~�c	�H�:<�#&Y����	��Zi��X�x�D�@�LRc
�����PH�|�����F9)߾����/?���P�Ǐ�օt�����7/e�M���c���K��Y�\cY8���=r�C�*蜌Y�I�%��w���ƕK�������!�}i�Z�܈ť�O���:���h^�Pϝ�(�������cQ�}��J���s�����`7���AH�.����w��a�T��\2ִ&#�5PU�p2�4}��a�Ьk��C��Q5�ˣ������ۘ�|�H�w��R	"
a�$��R�1���(����x���S<��PA/�m�	�
��@c�O~�Υ�nw��?
��bq��?����0]���}�)�@�`~�cW�i�͎�h@0R�'4�1|Д�PBD���#WY�H.#s��h��K*L�{�q=�JS:�z&�R��t�7�Q [��_�DJ�����M�7���d�p�F�i�ڱK�!ӝ6�t9�>����Vfr�Ғ�:]�H�/o�	�V��c��В����Õ/�q��S_�l�#���So-">��L'��5���.\���A���)��)x�έ����R1�s�?����o�P��	p��I�21h*Qɩ�����av#:����@v�5U~czq	�@��T�5����s���&��Lr#�
`�˲�Aș�(�\�s�A'͊Ia/*����.���`F����uM�88	�4A���7�Ӆ�
z�t�|\d�����]��	��#�.2#���P�s��e�2v���H��Hf�*��*���fGF����evs����|Z��h�ˉ�N}��Ҋ2�Y|[��j��>#M�r�bY�z�삇J�bQ�����*�p|A���C ����w9����P��J�u�Me����(哂��g���
�a5�2%���n�_��Ӥ�!�%�K���f��"~N�tJ���Ȱ���xz��2�u�� ��i�K�j�Pq��>:�[����}.��ڵ+h�jC�1�\�х����X\^��W�(�V�2ÄR�'���,�2:�T,*Ҡ+����s(X,������ݼ~	3ӓX_]�����1��h���=�r�<�.���$��l0���ڜn��iʳ�������O�T�ɶ.���;{I�<9���oa�S%w��tB��|�b�>�� :<�">1��ÍD.��ɦ;B��%oEX��i5���w��[���7��q��M���A��L")���h˛;��>��@,]�O�e�ݝ��l���O�B�{�]�7��Ž	,�^��ظ�6C���i�ȳ���DbQܸqC�ﳧ���M�x���:���������,jB_�|���gȄ�a'��bS���u��j�N�QA�T�\Yȣ��	Ã��Y%W����O��>w�Ltq��%��9ڦ�[�Jh?��ނ˗.h�N 	�l�Yę��»��&���'�.?�4�����P p�A-�Ho��6���������l���x��K��5�,-ʞ����WU#޹{G� WvmJ$a���Q�\�7��ϴ�L\>���X\_��gO�g e�$�M�������;����C������/~�G�����L�p��zjj59�U�ʏ��r	�܏iB�v��w
d�߾~'�CI�����)����V�S{������9��v?�,��;���f�j��4���X2|���/
�t�^IJv����v�ʸ�N�9}X���[�_ePC�*��,�2"�����T|�y�y�a FL,?ĺ�j���ʬ��(�52Y-d��CX�����;i��������+]!2'��ouw���R�}�	F|�rR��ki]j��r@d1)7S1��C��Դσ��!OV��%��V"�KƂ��A�OdMˉ��/�gT��N��W.�������5MX�`^0CF�2p�DI���k��z��(���i����ew����L
��
��/�3��M
	��No˛��:�@�0�d�;�SNt�-�����f2\C�P/^N���Y��G��i�v���1�=?��{�Ӝ�^�����)���	��-VOB��4 [4ɇ�P*��4��|j������X[5R-V���d;J2N����]լҜ�t����U���v��/�=�i4"���J<)�L헏�@>~ s呛l�������F:W��U��T,���*4�V���@�Y�]=ݸx�~����t��O����ޛ�q�Ʊ���p_�{�T���V��rBgq�EMD���(<��2��KRo�d�[����QH%�L��#/�`��2i����� ���P9?{�	&����f<��p�ꪑN����������i$�L�S�.�Y:Iq��]�ǰ�������]��E�x�<�R^���a��T_��2J��hO^M�dw���h6<h��xNB�n��̺����{w��P�w���_��qH�I�)�޴*�L��v<~5�əet��ZC�yo�����>�j����@$����*zŅ�����C^D(��000�ё32D������3#��jn�xRrp�������<����\�hJCd��{���VA��Ȝrq6(��U�{�������~��.� �b����B.��&B���d���fѶ��o�Q�\i�)�eSL�ۍ�8O���J�t�D��i9���Y�T}ܹsG�<��<��#Ix$O����nЇ���G�028��sc�|5���u����Q��_�g�s	�?~>!�;ya~����y�3�#Hr�:9�����Y�:�꯯�O�ܹ��SA�����?����GES�.���2^7�j|dM�:�D(����	#�5d�e2Y&�γ���\�������x���5t�l��索�O��I�	Mύ���]g}�'G�\&/��ťyu�L����E��yF�҆�,�ʧ�p;m"�0˗N=d��!T�b�T�J�E��g'��Η]f���J�5Z�~��޽{X�؁��Qv���=UJ�RA�\@6r�����fԴb��{(٫au�������� �a7��{��� �[D��kh����7�$���{�ppӀH�i�kZI,���n��,X���gE㘇O_h�E�_$����V�]�pO��L�$'sN��5J�\[�i4��0ZZ�5%r'Ll�Q���ɻ�/m'9I����G]��}������sA�E�l(1��͜�����	����B������B���m9�O�#��_�]2��Z[�(y�t8�l�M�!NE�R�AO2�Ky|p���h�Iy�l<��=��Ҳ`a��'���itN_,�4� BŔ/��?�{��\�x��``
�R���o%f���r*g�O䅆����٥���_VŔ���,)���X/�x�n6dk��v��Wu��?��,�^-f�������?�L��2��qR��3��̳Y�;��K��0��Lِ���]B�2� ��0�g�pS3�B�<�Z4��cscG�*}]�ǘ�ˢ��
�FF�����#o�`q}]��������;���q� �J:d�Y�Q"i��,�w�iv
D!��b��H�;�^�ҫo�dQ"��
����	��B�ȟ�(�a�t��܅��^�mo
=����֎������I,��^�l�R��0�RJ2$�ARg�4�~���lR�^�,���7!����Y���7���^M-�b2!w�',����2�6D��Z$3M���ѭ�(u�kJ%�BR��wt�)�A���C��Ze�Ϛ���������_ai�	���(q�9k��nt����� "Ek*-$�� �w��]����X���I8f�h�Ew�f3������ٰ�S��ۥ`�h���3hj�����Ul�{'߆u,�3x�bJ�`�[��Jf�[�872"���D*��?�H�_~�@+���/H�����U��p�<��/>��OKB*���,�L�����B����H��J[������ �\�|Vt��,�5N���򣫗��͑��r�����?��/�c����<�&�4�0Y5�������F�4�P�{./�}�'vRAw{��K�t�I{�B�{3/B�Q��fV4��x-�.oh*��"%qoCR[&��q��u''����D]}�a��p�RK)��dh\�Q���R�0����rG-9z�l�<�!��	~�[Z[�p9\�0���c�If-_���~�.̋ȕ&$���P8mn$�GX����	����갡R��_� w����ݔ���2�;62$����
:ڻ�x��?�/P���C����4hEPNGSj�ل��N�uu�l���,�/	z���D%>;ꊏNO����a��՘�'���+u��&��k��9�1c�/=v��e'��i�]g6��܏;T���uǔ�Q�q��]<{�{�C�dst��q<��_>^��B����r��L�X%ަE/���g��̋���'�0��8�F�tR:S0����f�|��f�(��������m���(��6�b�XX���Ȩ��{G� 羋DM��j�z�tJ+/C�ò��͙T�Y��ɉ��Y�����!A*��[��z���e��d�s�#���0���$v��:�Cx�+}���7��Y�$���<�~��s�YtQL��hlj�W!xJ���0a�P�d�K+��_�xEN�#��r�~f���/$�gjwy�8)���Q}}���I5>"���t�������4���3��[�n|妅RV�M�Zz�c�X��yp�AХ��[��ex��ळ��j<��Y�)��:���ծ��:�m
f?q'hA)K	,�⳨����?��t��i�ꏝ�}D�,�m�P%��p3åh"%ω��@w�L
wo�@}MN�V"�N&�������p���C��у�P;�Z�����f�/�Po�B�8m�5�N�k�(T��G��c|�Dٜ���3d���|�:#yfG���NFb�I�P���g3�i+b��},M>F!~��;�+�Q�5����P�ԣ�ε :3x߹�.�N��8o3�;�CC�������h��Lf�g��\�7�}%w���gG�ക�47���1�������He5�7��=�,����!	kBg3��!6)���h�"CA45���u�	��y�vu��~��4:crE����TTW�ww�f�u㺆�g�^ ���r$Z[���T�@�v�3Kx4�J:I�,�uS������\��o���O�����~���o��䲚���������.N�YdM�9�����!���չJ1&~�C8>:���+״]�����.���L�p��d̂΋BnNԫҵ���T���pOɆ�RN�,zkk�5�S��t"w(�7i��EOx�;yf�������CIX�{����%�o2�Y�yi��L�#��Hle���tA��v���q��>@pc��x�7������]݆�`D?'Yl��K'���E� �3::���0�_Mk
��8	rB7X�2��0�I*2��;[�p�'�GjN��y������:�j��Ӄ��%l��kjax?g���Y�
D���<�V�I{f+<�����[�Đ/Y��8�(�T\�9���ǋCz˧�"2�3t�2��L��v�,�� 6���:q���`��(��s�K�S�P�>��ɗ"�tv���C�X�{��٪F��8�ʩQ�e��S	/w�xlP�u�gv�U���������G��=x��$Ɋ$��?}��D�XF�%�7�2�M2��^�/8/�X���jjj��P���-��Uz�ّ���'���Z�"ћ����3���E,N=�AA�,�,��Y�m��	�Z��ѱ��;�i;��w Q��l�ѿ�M��cCHT���E�p:����W.�C��.�
~�TqO��zui��f����2�����ٔ�%�I��I��v�.X��c�$�\&'$����b��ҰY�p�)Ob�I$���������/5�@��P�l�h���\��������%�A�Y f7zG/j������(��Y�	m���U{$����A��
M�B��Ag���z��	:�-�LF_�ǭ�W��ͩ�I�����l�J�h3[�9�i�h�;�IFAg��Wc_��!�$;�AMOO�X0���ן��*x��&��w�g�1O��N�]`sEy���!�-�`kk�_����Tfa����2)Y��]�k�{�t�秤��́cg%�:��GH�}33��;���7����]2��}aSDinC�WFdm�2�!�KԘK'�2��煐���܎d���/'p+�������5���5zw)�#��0x�T1'��ih�����.6|��mA}9�jj.O��!���\��#E��fq��ň�N�&}���X�\ǳ9&_�5��S�0������+��w*�<1��g��͟�R}-Mh�Υ�H��c��+9�p��w��u��"�$��n��Y�F��@O^<{�*�uu�=v8�X�ڃ�D3�%i�OMi	id��]
sx�җ��VWk�&�I�s��O&^>�!��k8�����9B"��rRLR~��4I�х�v`��E��x8���^ւ��s��qQ��鈐Ӊ�u�C@Mlu���3#X_����<U>��c4#�8���78\�Մ^)�$Ž]�C�1�� _�����CwG+�}�$��������sbz^(��mt�*OLo��Z��8�3��y��<
��	E}m-�������� x���kڟs��y����oqUA؍&$�T�����7���;����vN��e:��+���^���T������6���ƕ�ek��1}�*�6χ&[-j��T��&���,�\u1f3��l�F�t"�����	��슘�l�H�!r����4���g���D�5<�ٔ�I�#��X�t��ۏo��B�,c�^����]Z>�]Hg��7+�O�C��t��ڢ!���y�&�m%��!-$h��NE����.w~~VѢlTΏ��v��ꦲR���S��&��=UA�9�"�_���Y2'�WE�B1��XP6�?�'�Da~>��m:3s�b���ErP��hP6�7�:�ِND�Rg�)K"���]6�ѻA�LU�� �9f��ln��,9���i9�v�M�3��݈	#D��*SB2W�{ix���<N#�Uȕ�ɜC8���:��޵��ƺ�b}S��uN��0��s �)�RA�L蕂N�7��.��h�hH�0\
���O�/E���Yg�L��ϟ��U�qN������~�"�{{?��dMD���ᓰ�C\W�xT��d-["9�h���jį�l�@�L"bL�Y�Y��Ar*ItٔS3�YȩZ���gC�HZ�̓����`/�^N���X�+�Dc�
�ܫo`J���K���AY�����Y�%ߣ��{����i�w    IDAT�`��͍�Jv���J������aGM�$�4�1���HqXcC�[�T�wISM@�H=��8<�i-@"��o��8�?@�9�Q�O��FO#�/���R\�pvpH�2�{8	�@��h�7��a__[��(���|�M��"�rmE?6c�䩜�*�n�����;��j�<Ø�}��/�N�	|z�K����R��%����߿s���]X��tr��~��O��+Q���,��{�b{z/�=�-PN)��H�K"��f�N�4,�	'��g�� Ty���Q}k���$���F�92z�u�Z(F|��¤D�<�tT#|h�C߸vvSNP�ᮾO�X��Q�S��H2�҃H?�S�=]ݚ �_#Q6�������_��ʋ����y��\���07�`�P����hnjW�����:!���T�9�{��7z]�0.��P��iB���	���.Y>��[�vw�������J�  �ǃH"�Bd@�\Yχ�>
�tv��}i���x�bA"�pX�l�Z��p613'�I;k�%DO%!��=5�T�m�z�hZ�g:L���f����~����I-��ޞ-}���1c>����.�ׄ�|j
�'	x�A��ȡ w��YЉް�7�����qnG�֚���=��)����C�N8Bo߀�,VĪf�Ȧ�Y��W��;�r~5ϴ��\.�����?�ŋQ_�E!rA��WO�aeuK�v��Ryd��٦uC�s`7O�^,��$φ���[絩�kk�"֨��L����'�e�A�a�t�K=���e���#�͠�{���O=F1q�ð���o��[}-2"�J�ig6�G;�T,���A�^\T��Ј�.�����/%�pN�+�I���zB�l��f��$��'��Lb䙓�B6��s��P�Q �ޞ>��w�a�x�����@��EP���uOU�N�i"GB��{X����"�}�2�a2��G�+�z^�����������}6w�n�K���E�<��T�P�ې;z���btS6�$/N�U����8�w���G��r�׶�Q�؈#�l�������l{�U�yz��U�TG�b�=L%�
�{_~�>_ '�cY�Z�y혉���[��a��7T�q����Ai�dxWX��P�ɻ�Ѽi��%5�<��7���ߣ�3����`j���yv��M=�k6*��(��>|�
:5պ��ɜ,�|ɓ"�L��G�,������X�$R3��;x���!����k�N\�p>�Eu�Ѻ�&��)��)y�p'Md���M-UFTj��t*�R��#񄉕�8�?@0t�v�&y�]����#?4��¯�7H���Y�Y3�¢j��!e��ȋa���EM}�qx����L�,bjy��tS����/~�Ε��nW��?*[���S���_����|�S.;��������f�"QnV_݈��!஝�h��K��,���\>]]�["�,-�byuS���D���U�SI�tv��c�c��r���
�l��	��Ə��N�T���W_\Y��֖�`B��4�d�I��{wojOE(��&,�4�`g�i||��w�&������_J~��&����LcccK2��=A���?����}����\v�b7��zP��������7#'s�P>cK�Y�i�H����NM4�t���B$X�� ����y���(�,�d�V�����*�tn�{��%c}~qŸ�|�X��*��r�J c�^T�orjV�W�||?�}����b1��>8���!�ܼ~C�qL}�*D/�Ê��4%}��`���l,`��;݆͖��i�U��sT=�f�I2G�.�l��M�uB:�Z�=M8�h�W����.'2Z�2���)'ϒy�N˥�{K2d�P*Y/�e���E��sFr���m���(d�$�R58�ܥ\���iM?Y��LML����,6qOo�\�|�~�l�brz.I^Q\�rUϗH,�`y������?���HJl�h��6�
K��`J��M�f1mp�ub��MX�M��(j�����*��7�^E"վ/�(�xd��W��dkw��⪬t6�
��/'�F��w��f������ܿH$J&�8�j������	M��L����Ѩ��|m����iL���ldID>c�����gCC�j1�߭�hvv����S�İم��큁��I�N?VA'K��V����+�cAg0�U�M)�F97�8�Z%�{���>Ovz���z�l��WU+%��W��pB��	R�Ն�鱦1�1��D��Ã#�}�s"���z1���H<�p"cL��!�A~����P}�xќ��4���� ޿*`~ȁ`�"�~2ѳYx���ˉ������%	���~\��
�	81��&�|	[.&ȟ�_�h�}��MԵ���K"\��M�T<|��~���k�u�00��<��l�I:��*�1qT�ݧ*�T���;
𸬸va��Ɩ9=�~|kg��1q�kS�@�]&/R2M�T�ڒqGRa�͉:
*��P,"�����`��&�h�uKT�j�P=.�⪕���H��a�g�(�-?O"�U~z;�p� �ǧ_}�p�<��� �j�%������\�7w��CA�M���_�Y�`�����Y�{�n`���� uE������)��<��`����5k�q���:e��N���Y�f/�J�dcCf$�?�{v_"=pω�f@;M~:�����pM�������F}l���Lm�a��C��î�_��$��"��d���Mh��4{;��و������"Y��Hn�u�lm�Mx���"	be�>6�^�ά^�au:�]�ԏ���>�y����fM����%�c�4�"E"w����ojS�o�����6R֌�<������\���x��3��F����he���%,�B�	5��J�`�����c����U�;-��������,�^�� -_)5�$Nq��)#rEKk���}�w��=c^+�#��!S,�ѓ�Z4�����_ z�CU��L����1�����Ȼ���j�Ć�ڕ�h����ޖ�qD^�����{$�㊇|	R7*�F�������"�3`�"˼� +���G6�.z,������^xDIx��׫�P���i�v�2��ڢ���H�H7���Aխ-�:{l����)���}h����}��'�"�p:^_����S�2�*�<��UM��r%g ��A$����$���;:p��%]�4��;I-�����P�dE2������m�+��o���g�6�� D�<��ϞAo_��#��4Ǒ�NN��1J�H�"1��b<�L����xѡ���+����s��Ӆ���2�����*L<ӄ</_���3'-�0x��D����x11���=��.I�V^ae��G[��ED�V���K>��M�=�|~څ�=)d��ނ��V574e�}�/P���M鄐5L�АJ�u�x6�j����c�sŝjX��=,/.�$H��(nߺ����#�z@"��y%W(�<� ���֖&45���/-�b��P,w�%��l���Y����>��׮i��d6�}8{v�KX]��3v8Ͱ[�{��Ö������);��s#o�S׬$L�
yy��Z����8u���,+����i8�����c���ɥ��!5.�L>�dpҶd22a�s�9��Z3ŤY��K�%���'T�n��7��'ǃ�+\nXK&��ڪ������m5E�(e:U���	�"�tо?��P�u[<�Pݐ:��@�ښ�08С �ٹ)l� m�H����;̙��������X�����gZr�.�D!�i����$]�B��W���m���9@�̰Nٔ^�I���Sik�����ITM1��,J6��!D����{�b��JoK�M�E���/<��L<�P�X,/w^>n�N7c����.��]C��̀z[�$-�]8��bcmS{�_��g��psZ�����Ύ��gΜQ؈`�� \>7���Bx���%��B�
�^}���p�D㭂^�<����E��⨕&I�u*ÍK�N��j����*})'�`���n��0K��mA�6��Q�9��A��K�l�8��W"��!�J�Kv��.l6�|�Į�e��\�鷦�Ul:RI���>Zy�*h���GR}]��c���/pO$<<B2F�@��cY,�[^i���m6!�����_����e����}g1|�=��nu��g`By"�	��}>�UW+AizfV�9Y�"dfd�o��/�rSD�CNc�B�z>�E)�~�2s!�qiOhH��t��^���뚐,����5U���N"
��!�Q~}�^ t0�ڇE�A� ZZj�fD�9>�-mveAq��?�����2������I��
z�qcW�A��C�,sIa������t�g��R����� ���.mmٸ�31�Z����5VCģR���`� ����Fnmt�#^BR"Cjv�Cp��zD@�:�P�e.:mi���A��f�N/��[16zF���|$�@�U(�<�dA"��ϓ�O4ǅ�WKf��kH�ی��i,O~�dxWa)�"�gղ/>w�&�jtyl\���b����nom���a�i��z�|+�bi��t��U��J5�U^�m��3G�3���D,��M���,�Y0��ťMA�U"9W��́��p��8rلк��c5\K���َƖf5�V�He�x���?�v�Ȏ�����j���R9TWS�>����̻�a7
:���L��׻��@m�0��j5�p��ͬ�-� ���F�����X�T6��q��{zv{GG�ͦ&�����h^���|N��&�������@���Ⱥ�h!�LA;�jԨ��Idse~O��S�	E��Xa%:h2��y�K[;"�:���.�Ww��������>�[h�?��x&�,���p�X$�ϊd�Ύf$'X^�E$zo}�LTA��ݚ�o���^��ont��;�7��<�?����_��'E��b�\�i4(�d�$� �q�X�Fpz�`��$ձ�m͂��#�[Dm���eZa�;�����S3���U�ҡW&t�����l����d��(�8S�M2��n���u��թ]]�<��S�� w�h)�*�0��Ӳ�I�Sq�Tl�ņ'O���V�dN�\��QL�,�Hak�P� �]���	�b�%�W'`�]�[��e���Y�˗^��/0��p�����rB�����|�v��o�D�l�f���ߟ�%b#�Q�j����I�ϐϔ/�;$ei�IJA�$��?S.��1f�b�Z�e<B� ^��\\�X��?��$t��/�A�a(�����ڢ��F�-��@\�9O�T�&ҰSל��?G�tO�z��FG�Fο�"5�44av�Ū�i!tVʣ��	-��z<pRS],`fv�6At)�*�a8$~�Zp�����\�r1WagL(;�tZ~�	�N�C7��4�]T2
���kdx��j�+�y���h��׵�gIM9�tf�����jy�\T�gį͢O�Z<JRS	'E2���}^�o�a��p�bp9�}��iX:\~t�|�����&c��z�޻w���#����tg�)'s&��J/7�:��`A���r�,h�j)7�q��񼑀f�+�"��=t�2��؄�l���Zt^xdwv�v��ssc��kB3�;�����(\-1�ec���+�!�䬯n������Ԍ���^o��s����ۘ���clΣ��@�d{SЇƯ#U���Q�p�<��0��>'��w�?�/n�|�{{0Y�0�ܥ�R���S��0*f�WJIP�8*��W{����7qi�]�����7-�+,N�.�߅B��83܇4�%'KH�3Z{���ECc������b������䮾�~◿���:RvH�{~��e�(B��6aq�L>�K:*��&�:����d��"e��l��ܼ~�Љ+ZԶ��`?���!�>�>�L��J�� }i��;M�h(V�6���j5��g<��� S��DI��|��=9��$G~Y�lr�J�4��z���j�k1����pD+	��R;��֎���fҲ����OG[�Hu���q��Q�ռ3�f�.3���=����lB&��}}G���V���l_c�_������;�?�r��_�{����~>�M��4�K��^P��>�!��w������q1y�k�P�^� ؏fkc� B�G'��*���⑰o�ԥY->�w�@kL�|��xʓ%?$�r-��v��u*B�;c�.k,�����	��s�������
��Ȉ����Ο?�߳0��?�l폾�1�Ǉ�jm6���+^�P�RDbqx��p���X3Ŭ��]o/��9vצa�V��eȽ�}���")��E�ٿ#Q��&FPR%pv���NHa��H�dZ>R7��'�`9�E����&�m�ƃ� iCO��
�d�����T�^0ڐr%�l��*�l��0<8���}I�דX�JOh��!�P�A��aKs�����Up6-���m`�g���]��E��e�����O���b)�К\�8oL�f� .~]=��|�gGpnt��� �SӒ�r�Ν�;�]�h��v���%�.*H��LV. NF<7lR�}�����9$a1�&��Kȝ^�t��o�v������41����p��=ǯ��Z��w	����Ù�_��f��9��9dRy*E�9���"�&��-w�VA�"�8��W�yS�y��>>9Qz3MK���ꧬk���^���@������g�a��&9��6�z�p$�#�_����J�� ��ن��F���p��"$O��'�2�Pg3��˩	=K�t�w�φh	'��pH�i2F�`����������{Z[W��qzH�dsj��2��+/q���*�]�d�A��E�]��S�
�?�i�HW.��Hf�J<�P�e`�9uL�;@�^��~�O��(����6cA�/"�{�*�����d*&�QSs��K�y���K�j)j@�Iޅ�M��kq~Q����(�ojj�Z1��J�sp�'�6����#=g�{"m�r�{�jǡ��6�ǌ���*��TDֳD�*�;w莪z�#��]���'����k���濫����a�˫��܂��|���yJ�5�|��b*�����{��O�����A:]ԟ����+t�dɱ��lwj�@CO��� vV��gB�˹98kj�����jP\^]�>w��W��¹�X?x.y�Y�{�z5�LN�p|2��Vd�a��q��5���������߻q���߱��(b���L��ׯ�����RtzǢ�4
�L$��30��q������DsSv�CJ�b3�1h�1���z�t���r';1��*{�l�JA'��Fr�����z��]]>Ɵ�"��润#e��Sa##�/w˼xI���t^�v���+
�p:�8�"ͮ�d#���~��������)�	O�K#ăK$�B��L���%##�;)SɊ��^�~���9X�i.Jf�zs�9\��Ds&u�4a���j2Asm5�^:��c:.A��q(��㕵-x��˺VÆ�ߛ>�2T̟[e!����4�6�">t���H��_�0���D}3�c,�dm2��2<��f����S������]����V%�3�s%�I[���5=o�a|�m�ҡ�iĒIe�o��SY��З_�
���VN6vd�D���*��T��H �������)����dm}3sK��	�3ԇot���*�*�z�(�+%5urڔ���%��I�7D#9[Gs�l�-dw>��У��J#��^��o��g��w�a��h����MM�Zi��⟗�屵����ETU�"���x	�˘�| s��MAOf��,� ȑ���gB�.����X/�)%�������.I��5�
D�������Rf�Ӟ��93���nB� L���2�݄tB��BG�4/9�;�ӱ��������<�z)wcb����z�ݝj(ɸ&3�s��˃��:]�ܣG�1�����6�����ח^bs�)�Ǜp���t��7=Iӟ���d1��?Nj�k�}`�OP6m^7wv4��P�0�*�+CY��    IDATĦ�b��oh/%cB��)G|>|~����b���#(��0����Wբ��U�'�x�
�z��z�hnh���{�-�q��Y�B�xױ	b��Ĕ�,ו�r���ѥ�Gi/���f�qt�2ĕ�͚���#L�0
:�vvr%'ʤ8��Fg�<����0r944T	�e���������!��dԍ-��F����}�!���V��
:�\��������>C�]�	�QW�U��6�ǀ6�6�\:P������L��͒n�-/���dBOs��l�{(C�K9[��D�JD��p��w�S0t���.������a��Ncx�W��S��O>�n(��ov�\�Uۭ�ކ�����K��;����/�ͣ�l�Ռ��Y =@¿�ӧ�.-�b�T������H��eފ��cu�Կ�׷L�LM���nZ�Z�?8$���g�p�HJGʽ��N���4�p{Rɋ!������ˇ��zE�l�b��D	��" ���zT���u�֔e@<���y�	�� �`gJc~ ��%�������@Jo��L�XDr�L�3����"Lɸ�N艼m}q����(Z��$�����h�`�YE��-ͨ�����Esg����d4�N7I�=���zeb҅*�e�ؑ�-�ˣT��mjiVe'�ɞ�X�]�.6M�?�<X�9������Q�6'�c=߹�1��kt���}����\�ρ��Ei��&�x"f��(�pJ[�jf^M
�xs!�xx/����Q���5��U���%�Q�/���Q"��GŐ�g)�2�C�z��j�z8f0�����]���!xr�G�0���:/a^���c$��H��v�� øY�>�Ԓ-Kn/:c�3��,_~Z�q����~��sy����#��{ﾋ��u���g�=��@go>{$d�F;D��6W0��+X�4��g��vAg>�&���m�EB:k���h%B>�������4{K��S�����Q��C�;Z��ߚ�59k�Y��2Ad�l�N�Ő0eT�DBf$y�d#NbS�O{�e󼿿'$d��9tvt���~��O�jm�9�އ��OO�RD�Mn����(��D��yt�4�׊��6�`oc"f���s��	�ۂn��h���T"���!����"��Q����i8%�V�%��Y�Ig>@�@�ʄVʹ*��u�|��b�&��p_��8ܭ�����Әtڵ��z�O8��>���n�E΢39gMLM�N������"^�r68TI�^U������G��=�"h��� ���o����1i�i�J|�3�n���PN�;?�@�%��rz�Y@"!Wqt�L9LFG\�d�{��@CUbx�HrFFz� ��'jȿ*��T��$�qPr�"���Q�0I��s��߀�l�C�,��_-.j�OC�$h�h�W�F������z��$�V�qJ�76��Aǔϣ�ևt2���5�7��T�?{����\o}��~|�ҿ��������Ͽ{r���^����?�Ȥ�H���ڌ����O���'O�"b$�0^���ēN���ᒜP̦��֮˕d$�EYݯ�ܻ���"c�JwZ��iZzâ%/���4/	K�&�h��cM��%����<�)�e�({Ԝ���AE�1u�,b��)���ϝ3�:�9�{��o�<O�6���dؿs�C�������j�i��<�N��Q�G��x΄��˸t�c���(�jJx@�Ka�_6N8Ό��p��	��$9�Α�;s����oC�T���m3������ǃT]UkX�2#�{˲)5�|iy	�`pH٫��T^0�"�R�b���z����e���k��]�tk�X�_0$2�z��186����������9ؑ�<���7]�d�	}h�]��K{o������ę��/1Wzvnk[��?P�;!��h�m8�����Ɇ�X��i�Hx����B�t�IY<VEJ���>�������}��eSD���R����I({��
Zo_�������4�՚B�70�߇s���ͧ�6��iq�p:=x����ٌ����W�&�<��ܱ
:�)��ɀܯ��'�T�x^���f1��	(��0!/���V��2��k
�̤#������W���0.K=�Mz�8:8T|���FKS��)���}�I$j��
20����q���QERJ��0Z	ao�@�K�Uɭ!3��,A��M��e6������XD�z}~�.,b}g�,�4'��$v�g���L���J�&{�ot�-��mu"rt�ˌ��z|�[��H�[X^�͉4t�:)�K]a�8P#o��_���uғ�"�r�~�n�")��F�*"j�}~?����ж�5���ϟ=��A��:m>~�~�}:���G�g�h�}�cs@�[M@�=�z�y.6�vawVk���}i�!'���y��l����ѫw��+���#��5���Ȥ���S (e���}O�T2��3����
Ht��F$��E*�B�2e�W:����͖��S��J�ϲ���sg�'铀&%pM�mpz]r̦�hk�G�ӎ�����r��W�_�\���6�G]c6���r9:9V}��q���Ω�$�ϑ����>��%C���&�k���?�D]} ��>��}���=���Ò�m���ߺ�?|�������_?�`A�$b�X������lFkW�<���k���!R��T�~;�X4$�۞�6�UUk��%M���/���ň��L�bn��	�%ӣA1����m�\&-~���CIƻX��
e��E.����N?���-d�"�t^,��tV1��P����졯�W�
F�K�_�Q�$�]�z�L�3S�o�-v�mcy��
z1{S�cY�s�
.��)ؑ�>�	�����>k}\�0n0,-&�()[���#|FӐU�����W�$�{+�\�R�W?�"Yٌ���N�c9���r���<	�S'�:�7�|���.Nwp'DM%�������⢱������ &&_	���֏�Hw?�P?��ʊ� f6!�Մ���{��P>��C|a��(Q*h�E����Ӂ�с��d��{�ꕬY����"���j$�4��t�{^��J�!��|�|�Dnty�S����ɤsz�����l��K�ͯA���sa��NY�}x��wp�ԅ�?ogsKύ���6�o<@M�J^�tKdC9:6����H��k���*f_>ЄN�m�OɜU�C8{��
�1�[�N��6�YM٬���ϔ�-B�߸���Щ�(���%��*�|~���_�as"c��B��D?w�4:�YW)侰A��T�'x���&Ԑ`���q�SY l6O#�.����q�v��/�>�r~&W.^й���6v�V�08r˫��_�ng[��X��
��!,Y�.o
:FR��HX��yuq�u�AM��hH�;���.=����W|hG�8�~P���]w��lFQJ&bB�����(3ޝ*� �U���#<�DXę��p��(���j6س�sZ�x��084��I��-��ڪ�yMm����~���kuA����n�m�b~q]=��R!���ǘ}� �LT�jw+?��cg/߅��E��%me�c2����062�?�`���;
��9�~�L	#�5ܴmN����RE.?3���Ap�h|E�[�
��)��Z��Resͳā��/��hniB:��K(;���̿2�":�����.X���9q<H���n\*�Љ�cg9��w�??���S�ۈP�p���ր��zTU�����{O�Du��t��x�ڿ��۾�N���/_�����[�#t�)!���	ζ����f�M���@�yV�`�;m)�2�!/�1-V��w�"vuvʅ�nP��<\~�.d2�+;���^�2+� =�h
9�HH�S���<����;$�M�<�8���Op��yM��S��4����W,�`�&���dP=��E�
�߳�ӵ�Տ���GsS'^MLbcsݸtbI�#GX��:x����#Y������� w�/�@�[��<M*�:�P[���g�X��;��ڎ`$���ؽ^DbI�Q2���6���I�'&J0x�C��I�6.���}�A�Y0&��ݤ
b>�)���s`�:��$��B><
�;;>������.N�\Yp�A�!f.�����YM}u�`��V��?}j�'�Ua~꩑zݗS!w��
]�1v�{8�3�X�O�f�f\:7&y����n�?;:�l����-��2��{��������r��:
�)�ǅ�X̲L��>7B�V�Mϔ;pB�ULP
������s/�sԯ��^Ng���2E�w�N����u	n�C�:u1�%�bzi�h\�3��W^am�&t���rRy+j��`�����<H��[�E�F�r��έ����{`}s[�?��i˪t>��sOk<�
۽Ҁ�8��Rޡ����0N���QP���q4�~�<��.���ǐ
�O��y~	��Yr�E�u��@��\|���yWp��UZ.�U<;2,2�ƝbB>W��~�݃ �O. ��lK��u���"6w�v��cW�y�D5rg@��m���nBC]�
#�?:.�kk'%�e�8r0�j��d�o:5��]h���a	��lth\�g&�?Ϧ��D<J��{wo�m�v����!���d����W�]w�����:�HDcʡg�a,-����ciqE���[Z��=���䢔�%r��}q3���QL����fsr�Fm� F.P�ޮ��Bw<_3�z[��z����?��3F�<?{*���s���CN�����J'��lܧ[}0l��؆Ý�N�.�g��۵v�;���d�l�s�9VuUWN��U������p8$��}��_|�v�l�A�&��)�p:ZE���e�
r=4��\Q�WZɑJʵ�ZE�fL��NJ(|����6��ꗅ�Po7�*0��v�6�[<���M=���V	2��5��b���3פ�nLH�#�ϙ�����p\��ވ|6!�Z2i�)������^l�l[���~|��������G7~�h�O�p�1٥R��ίQ����O>���Q�b}q��Q�m��C����ǃ��t�blh ��3�lmn�ࡥ�C�)x�e-[���.��wEތ�)�I����84�!�$����� m
�pr�`�E��W`&RH������z%�h$b�j��§�L�(�l�����NC��z���!N<����yh+�_�x�����L4t�f����>bY�:XV�-����f�uwh?�j��4]=h��ă'����� ^J�%�A�8���Ŏ�nLCD{�X�d����j]&l]0��eGˎ�#<B��	�i��V��C�7���  U�u
�T@cХ�;u:Fqd���m�ײb�����,F8����)���ˎ��UL<�D#�RB7����u	CW�G8�U0S!Cf��cRr�����������P�}��2bB'}�;[>Sɾ��߭v�"��D�☝��A��6���^�Hx�=c
�'������ЉCOi��_'咂�;��.�ħ�{+�N�:�I�yn�S���G'g�� M��E\t���42�Oԡӵ�	��y�7�A�D@av�Ujx�3ĘP��TRee$Sq�wvcfv��G����&�jdy�7&�R�e���aB�q	�65��&���,(l�[�t't;�Z���~�*�^��g��r%F���	�?���B��9����p�^D��hmjTw�����	ZSSOB�[��>5���d��_�tw>�"࿕��f�T�=��IM!c�|�f\�2���*���q|r�	׃��!�5���Y�Z�JSJU�MC�v��_���L����{,S&~���W��n��������8�e�J�{Z����cem݃������<^��Sqr$KP�=o�u���_h}�I��ܼV-��w��}���%"��~�0��>�8,�r�:�5���.߁��I6�.�w�$�KE��������dz�᯶�Y	�����݇"�R��<-���sF�ա�XI��dX{��2S\F1����ɼ�N����{�8素�VfC�|=���=��L�����8:һ�o�:�ϐ��TI��ą\$�>;MJ��Nł��u,.,�!!_=p���	>��|���#$H��Ѭ�(��|����˟ܽ�_���X��������_<z�V�����nW?�w��&�47���^t�v��q����������$�|[�/��jA��@Y�{��������h����vg^Z��*]��n��ɩv��bQ\����͈��N١'�R�aB�^��]Z<�,^(��g@	x}�*�\t�V�$��P��s�YL�a���r'�{������G8�](�2��̆M]Wp�ݏpJ¤*�p	Ka�@Ķ�z\�|I�q<�������G8|��¼y�É�"�K_R���j�j/4ꩩn�AG�����q	jL�~d)�J��|�X|���&��ύ���R��dJE���� @\wҧ����
�����7����l�像5r'm��t�����.���E^���g�i�c$��:��+t�r��L$�x55�}�>�n!dK�7�7WEh>o��j�+�ݿ��D���O���gRϯ�*���1�c
�J��s%e��^UU�_#���#�/�42�PGK��r���?'ւ\p&t�׏�9/�&*$�3O<�{�%��Cg������u�7�A8u�R#cb�4���+�}S/��K1%����#��Z�5�Ƽ�B�bd6ޜ�;%��&�Ϳ��d��Č��\�$1lL���ɪ�G�L��u��\�~A]M���Vb����s�E����fm��$��2�k�Ŷ��ahh��C��xW\#�5r_Z�Swτ��1���qn-������Imb��5bK6��pGkf�_k��f�������	(-�Lў���FB2���$����X��ZH<P�P)Ԅ!g48��I��G�WG��h����㒩׌�U՘����b��eG$����*kq��Mٌ^\D��+#��W�T��r�FH���������(�Ͽz�.ݖ�)�����y �W��W��e�&��A��YRE�:�U�h���\A��<�D4N��QDQ��a`Z(|U���[L��,��'<Lʼ�6�MkN��|�xF	�̗���5����E�M&	=�9͠? ��Y/�/..��g�ᙖ[(%��Y��`��ό�l��xEM-������PmmPE5G�-��x<�S++�ЙЩ���r��_�ޭ+������ߚ����~��'O'�����iK]>x�&��c�l��s��wޅ�����>�c�����Ywi�A�$��4���=�`���v��an~Q�$�9��Jh������V,	DC���(�4s)lAa*u�'=�7ݒ����n *ͦ���
��<C��M����0jT����u�2�v��y�x�w�70xX1C
�A�/H��k2ga���e��Eq��:n����J�]v��,������l5�hinT������:R%��+�{���\��~�����31٬�� �">'&'>7�S�`H[a㈜ܕ�C'Б�� %~^R���2ق�ϳ3�ΐSo�n8��j��Q���wvz��E�dV+�n�Ά�c7aos	SO?C2~
�n`/CK�e��E<ie��	Af���sۭJ�f%e�#ޅ�e�r�5�(��v侭(�YJ襤^��K	ݠ������$)_t�"���u�D�F�~ҡ!C�ަ��ɾ�?�s��Xq��?o��"����lGSC=�YT$�2��6��a��F��J�I��չ	�.��)u��Ͽ �\�����$�UpbA��,W�ą:��.���]tM�m~���z<}�R��r��rCj�9��d��w�(z�yCn���i�[Ԯ�h�W^
�f%����*%k����L�Ѥ%�Q�K�o>>�Ӏ�;�ֆ��|o�`�mA�MQ�2�e�*l��4��z�
�;���[y���U�X�f��^���K��u�b�	ݜ�����
�5A�,��`_񄫲���.��صڽ�P%<��m+i�ӡ;������^R%��FExv(;=�y6�Sq~����р��\P`���.�������Q^Q�4Q"    IDAT���x�b��G&��<�? ����0�g��g�{���]u�LNGF�ٗ�5r7g�!ot�5-���6��F	;�j�4�	����W�8L7���3r�ŮBR�,	��Ɗ�l�6�Y�}+��޳A���p�h�	������ Z����[���XS���VX�9M4���0���	���WDю�c�5��MX]Y��⒞�;o�������FA��+�Ӫmh�f��`�݉�r���S��?���n����wF�~k.�����w���w�[�kB������=�\��&���/���w��a��&�������C�^�A(���O�At	�:{{�#-��������xxqi��*D����"0G��b�2�H�T�FB/
�P�� 	�|�ҡ/%��:6V�i��D�`�*u�D���Y�b0���+] ������*$��f�?E'9��Y������^}���9��2Fn�ÍӋ4�/��Ko}��I�j0��:D���5����ݷo#
��ڍ[�=<���*�O�G�ыbB*Ip��Q����h�f�<����<t|�G��\#��Q�w9*������1x���Y�������e�]���'��1�w���ʕKn_D��aGK�"�tmV%���5	�dRԳ7h�L��л�n#��:����I )/,(:�ۅ�Y�{��?9	龱{�ۋd���IZ�r��0�ݡ�g��E��xRQ
6�״�Eϟ޽�(N�a��8U��hS٬��@��E�|A�9Z9r��g@:�]~6&\"���Ƹ� C��Su2K��Ƅ�I1���&���I�ɬ��71x���	���(����2)�=���{w���$1R��VW����0�ܑ3)0+�
WR'��5���q�JS3�k�g���C�#a�,r���3tz��P]C�ٹ�1;/�;�Q���g���$�{xt��ǵ�r9��(e��^�_��'�F��;������`���^(%��ٯq��� ��2&X�uh�C��U�пI�2�%�b5�02؃���)*sp ��p$���_�$�c�������C�[�b�R'�w[�T*��j��b�����dR�%S;����hc�ŀg�[�!NQ��L�����ʑ񓉟�w�g��������dV��A��5)@����p��(��<y�$��kw�*o@�l��?������6��ڑ�%���hh�GGW�ZL��#��jz�3��.�W��J�ȶaYbD�-�@L��0P�L)Я��o���Й��P�D�|��{��8Z�l�����Ů,���@[S�&
++���nm<��[R���d:!�a�o��>�W���@SS��}������O�tr��`�P�9_��-��/~���?|��e�&��g�����?��< �x����������h$�Lށ��(�C\B�=�������s{}M�?�$��,t���]Ѯh�t&��-�]J@'��H�C^�TJ�bL�&�¹�.Uio��"���jfL���Me��y�*#x������L@;[�2�ר��C��.�p�14��MU��@5�ĻN(0x:!���ϡ�Ţ�p�:��0r��zg�� Z���B��\!�k#C��
�Y[Ç��@`us��_Lh�dq8 K	� '}7)�Y�2ZJ�F�R
F���?�V��LR���K�N	A�X_�`�+�k�59��������V�M�\�
�@��F:�T�˧��d�O��+`�p�0ʃUZ!L��8$e�|
��mL<��L���^
��:+$AJ�(��QR3����b�%ed�}���S�j<}9)�m*k����"(�	�ԉ�C/���WiJ�gc�YcL�w ښI�T�Q�]����rdhX�TvP͍M�d,�Ψs⾐&+��p8����V ��z�.��t���}Fr�����;�X<��OIЂ����ݘ���_�:G���]�L��iC��i�j�	N;G�簙���f4��beeY�P�����{�����t�vB�%�kQ�,Ǆm3��̖�g�n�Ϝ����Q!��EĐ����8==X�I�,"�%MBVd6��(�d��`�q1���_�`�7ơ�L��B}�C	��9N���>V�whU�<� g;��m�g�['����+�rgB�a��ڊ*��2_��|eЋѡa��C�]$�����ܾ ��:t����E���W��t�����D�S�(�$ʢSS�����%���:�+;O���i�{��\�ѽ��Cc�����2����gw����L#��=�h�XJt��n���ӯ�$��l��u�L�βz)52������TI����Z��N�������5���(q�f&s%�	�7҄E�˿���5D����q��Љ�$�2�I�a�4�K����t�CE���^�mE�Sc�{~!/>cG��H3'��M��u���Ȍ�i�j2F�m��;t�͆�:��4~��/��������C���Y�h	������~z��k��&���_���O�7�O�������>�}~TY궽�..��w����6��:�\��J��`P��'�``pXA`ec��
u�^���.Z�1@+����1�+rZ%.c$o����S�g%C�J�UT��~U�!�΃\U�V�ݪ�hY�$399)kJ\rW�n���<oy �R9VUj�'
��6����	�`B?�[���O��1�
GV�{I0x���T`%��A���=��9j��u�@q���x��F��>�ꁂk�|y���E_�AH���*V��8�/=;�z)�B��4:�o�������5��҄��,�M��� ##C��.���L	��DSx�� j���-���M&�@�#�6���eը�����^LM��̱��J��=i�r���C�����[{�#grkU#z��Lc������{�-��8�ZYAOO�.Ы�,MEx�,���z���v7^Z]�p	z�4�`������V�k��D�#�q�ƃ���ȝ���?�!�^�c�Eu��:���Ā�,-�8 `��e����I$2X[����!N/�Z�0"�b1�쯽I��q%KYQ�4���!ar"�3����?%���s㑐�-�W��gbr�G�g�q��GM�"Z�A�k)�#�k�Q�1��0�g��3�yh9!��v�`$t�z�W�� �Y���nt�Ē466��_c��������1�|yI}���3*힩ϕ
t�������#2}�{m�Z���ėHF��T*k��S�&��:t~�g@�H�������wVsO=Fcs#��q��1ڈH�IX&K�s�z)0���M����k��)i����8��y<��҆*�MH|���,T�3�zt�FL��m��:�N
�n�8>KC�tD	�ϐ�,�+�?sy�bɄlK���ă7��*�fj[���݁z5%�k%G
����
�V\�4$@��yX*����\Z݀��r�G#�}��ʧ4��f��"�$�z(��n2(�D���Gm�<�4��4a��*PY�ǩ�A�/�S(w5��8�����%']S�G,2
z�_��� ���Æ,z�W��l�Ȁ��6�;<�(Q��4Ѫ�2�=���p�	��R��h��\��{�o��n_��oM�����������h ��m΢��
�MB֦L9%� e��8��`1���v�kTH�U�(�Iu(���<z�瑈�e�M%d��`�ʛ4�l�٥8�+ڦ��S�<��еW��=E}��A-%.v3L������Asc=~�W?GksƟ?C� .]�,�h2��,G���	��`�ͪ��ni��C�����&���P\#��hWC���,M~���y����fy��@��]���Y��>D�#�l>��,�_*qϠ��\jv�f�S(c��T T$+Zc�'��,B�7T����J]�:���IZ�K4]}ilD�'_?�?rq���v�=lmlK%�&4 :�Js�>$]�U7��cÆr]�H���d��%/	�qm��`g?�1����bBK�`�J�]+'1�t\��L��x��&�mxx�/_���"A��:%NExƸ6<���EuBV�~�hl���3�3}������x�D�r��5y�4�H&qixX���ϟ��d`�<vINkt�����4jfnV�"�h[g���a������[k����@={!�si$2\{x%C��0���q8��ʠ�PN�8&��p��F3���WVb���'�u����qy�S	��/L�T�"��|{�'~��_cO>@c�w���{����xa���׹��:��7��PB!����ԇ�=����*�U���UG�V�4'�^�膌���%�����'��g��{�W��������X�9��jJ�to�Sp~��Մt�#�z4w����i;J@���E�,�)���&�w��ٓG�riL��;�Bj�l�A%��Ɉ)��˷��q+���u�F����2Ϡ��?�1�d�	�0���+���gs����}$`5��j��_�y���b�K`w`mmE,r�9U��Hk�a�
�M�B6s˛8;k��g0���v��B�L�S	��m�����(�V<,�l\���:��(�������Vl�ak� &�C �x�9�2�(~~#?������]�PV50\s"���˨)�'��?:F,�VwΘI
��\�Q��6�S?>o):&� ʤ9��(��qU��ڊ���NN��U+L�=h���Sj��!�`*�-�O�b3!k3#ʆ��F2K�U'|�,��?�{����O�ք�G���7����pxk�T8,���{p��wz���Z!S���9���1�+�v�@��	Y��H�d-�Mhl����"g!��4k�u.Ot����ϴ0 �
�ؖU�����U��Ob�0�`�ȕ�蒴'6�,<w�.�1��9�U��@�=m����7��u���KU)�Q(�ïC�^�L�(� 0`�mDO:p���-� v6���';�s�NIe(cv�s�6����p�=�U\VR��[������dK_�558�ݑ /%���i͎8O"XQ#����,�h�w��)2�i��u��2䉲�7��������C��A-�>��SuU��+��{{��3�oi�}#;N���������#)x1������Fow�e>���}��!�`X� ���v�����0�䀴�� �8�^���tޅ��+��.u�|�*Ŵ�EX�>���������jgh��uQ8!���@eE��x~(Nr�@"�ci�-v�Y2�>��B�C]����I6�K���\���&LL�T�2��N��h����@7��S��`U�:���֟㯵�w���M�^6ZZYDm]����Ƒh:�@0X�d��@�%t�_#����X��=����.�&uJ}Wn�*�9�%u)��bS�J�G�Ν��0F���y��T��q���KD��'�O~P�Ƚ�}Y ��rb�^��jο�7�7��I�7�Z��.���$��pd#؍�AD�/���,��)����_b`�_�$�"��3&u\, �|�˂"Stuu�A"Sk"��䔻Q�A���p���噯>�^$���lAS�Z���C�mr4����4rr�2���F@��Uc�~��������.�_l8!@�u��qz���(̻��)6	�C�[ʥ121(��5I ظ��^�&�=>S;��D1�ʕKRZ�[����dsI�{UT�����d�ϒ��_�`�R��O����֕�f����spZSX|�T�9�}q.ol~Դ�o�-��ME��?o�)!��*q�҈@e��7��b}k��s!�3��d���%		q��"�S����0�*o��RR+��?kL,�ȥEڥINk�����0O�9��'.�
���XG��}3ڵ�+�E��D�H�,2��Nr�*V��$�

�0���f��k��X�l�F\���`��y�K�vsA�M��߽y����L�����~����4���0����`��~���|�8�����WH�(2���.�*�a�¸3+�ֲ��C��,z�Z�qG�EE]���w{�K&�<��8�V�	�1ِ;�����&��еR�0Db�=�"cg�@��$��R/���ET����l��{q�8�x�w��Xp���xK{@&t��hLR�ǌՊ�����]vZ�T�C������2++6��	�}�6�.�A,K�LNz�S\#�2;�.8�n��W�C�))%�FTTD�I���������A�>�>WnV�J���'�P���U,rύ)�q����Ο����#f�3���ʘ`Ee9�~���0��Q=�z�.(:�g?5�`PmVz� :E��֡�jkr4\( t�j�]��Ɋ8^L� �$�?��;�S�.�{�*�I����|v�K�K, MI݊߃��J<F�9\��p~z>��j���w�ս38���ǋB}s4ƕP�`х7�qY�}p�b��\	x$ ��	G:g�H=/�#pd�x�8�ݡۧQ-��p�L[ś�n��ubqis��C�x��[����,���Z+�p8���-�noj�g�H���=�x�)����X�%2V�2{.�B�l34�Y�ҹV8�Vdb)�Ic@�$a��7؏��]M��n���o���˫�n�T�5qߜ��1xfw�V��tdw˩GBL���r*܍�u牎�ʉ��P�����������MMx�b�}�JB�^j��$�5ٳg�L��F42��qz��8cR��*O�Y�ϋ����X|���v��X�@�
Ɏ�1D�99�1�2u��3��wg[�\���"vv�q��u���a|���y��TN���h4$\i�C����bV�h%���Ϣv��d�`,�\�.�?��pJ���!��hi�g��Xw�B]c��oo� ����O?Cwg��B�w�6��4Y��}z�L!U���Dï�5r��_%OJ�Z
X�~.��B�L+�ف�ū�N:z��T�� �,��l��W:�������8	���1��.�Y.���f4m��SPMS8�}:���STÆɜϢ�E�8�3�t��aN�:�Ϟ m��wa�Y��nE��/쀯, ����v��5k�eR=$�̝��a�I��2p�����˴n㔃�,��<}a���	הy(?L�Vv7qF�A�'�S�A�����o]�?��$��/~����4��U3w�V���0���T�����=��e��8��p-�ϛHO^<�9K%�t�!����ىk{C�\�(dppx�}��ի}q4U]S'�:C��H��A��*'+9������)*��Ғ0-R�D9�t&�Ŝ���FOg�4��W����q�B�Z�0I�����Er���������R�!�A*~����*�N�}��V�o.cs�z��0�o)r`r�k�.�Go�l���E]h��ĤD9�)X�)�Y�y	WT��5z%�|iyA;��~!N��}pt&Z��=�)C�۝"�`�*6��!=�
�����]-�]e���.?�GcC-��AZcyu���v77�|�z������p��'O{]��Ɔ���<�l&���64׵itId�������-9X�I�O6�CϦ#�|���UB�����CC��j#J��0��L�8��<G��t�BZ�d	Ѻ���LC�����>��1Cf����Z��\�,�~6^Tk��h���XDZ�nu`�|��@�K��,<v[�u:����/��6v��K�x�t\�r��%�x�'g��z\�4����/1:؇��VLMM�dr���3S�;ؗ�)�#��x���L�(C�]|�Α�o:�j��Q�!�n�#�;,X\�EeMP璝���%]N�Da�>{)3?-vM9%qi�/T�Yp�C�bF:g`Q���؝+�bb"O\�LJBAE�����щ��6�����_�~���G����Z|�,�yO9�g�纞���	�%r^�gtfL��+�2�ll-Ob��W�'°[MH������;���+J�en��`�w�,�t*.���yH],;����2��'��($�.�E���o�z��1�e�
�!Lb؀�{gS���A�U$���-�"m��Uἵ��Ǎ��h|O/i��Յ��f,-,
�D\9�L�/_�B[{�l��~�`:;3���ke�    IDATx˂Hg-�٭|i�X����S%t��YH[k��+�e�A��d&���p�ͦw qW��19~��o0<z	�lV�S>?�k)�ʢ��E�j�"�0E��a�m�"��J�`>{����Xy����{PQę@�m�*_�?��h��;P&���GW�p3s�3ڙ3Qs���������"m�9�`B�_�}b�W�5g���
+c,l9,m�!E&��&���2%tףݹ���t��;�B�`�G��?_��'y���{��` �u��C��U����k���7O`������צ�]���1�c-���!	Ɠ�t��a{k�M��C�*�����'OZ��h?G�
���)/_�l�5�����Թ+�z��QB?��ю��Դ�&��ۻ:����D>0;��>�H� ;@Ŀ��g�w�=u�,&._�g������5!��I�	x��^���CCq�t&JR����D�w�1�.�K�H�3<�U�;l���y��칷.'�0�Duu%::۰��m�Q�v���EG�FRM�MKW����-���[���:�aq�Ʉv������]��ш��l��^��"|~�$�����"���s�{��wv��u�&�?EkK�|�秖4����yX��L�~�E��g��|�9#�P������.!�b�u�{��m�ŉҦ��Y R�X�E�!�RQ����m���V;�`y9VVWq�"kva��V�G3;n��J^V;��Qeg��G^�I��Q%*E�S�A���'F6���MF0�ي��zu��#�V=�|�����fg籾�%]��w޽���U,�,cxx�m-x5��G������(��S�3��S̯��4�ىG�ْ�{�H'3J��ev��@R{wv"y��B&[����9dQ�������ORV��ޡRmm��;�t�9v��5��q�Y�04�j��%��W4��g+%Y_%y{Q�8�R!I�T2%����`]�8:>���ԼhjBCc=��tx���x�u����D͜pUR�\���.��BD[>\����9���	6_=�:��9tY&tN�r�'�jV(1͑+��\��Ac�"e��mpxD�Z\ݰ�cܣ#�;1��W�fP�F����"�3�:V�x�ƈ�T���"�8_ ��Z062�/A�tG�J1��\g�V̂�үܵG��MW0;Ae%��3[9NN��H孊�D���Q,�z��WaI������aB�vO�2�dZ��	j��ObLq4�7{����Fj����:���s����������&@�dKbOT�cqS�0a�Nf� ���&DyӇ�;N0M�ݔǵ�A�bcmM--�]\ƽ�}�XR�����CL�|!3�g��p-����"����>��bLD�p�.�G:�ֆ47��岃ċ�	L-�HȦ@Z�Ʉ2�	-ף�\���w�~{B��џ��0����SV�lO���X�ю^�������ɼ;!8]^%jL3�@Ň&���䅀S�@�C����Z�Ң����M�l6�]��W�3Ec2���¨��:`%Q&k^ R�K⸈���I}|���s�ژ����u�
��<v6V���]:A�洘�r�D ���:LR$�޽���(;������eut��,���
���5۰�����_UB�ċ�:L�7����Q�F�p;ݰ��t	�rzF�\m�n�O�iV�N�W�F��G`��PV�UG�ŧ����]�}R�ĩvDt����{,�!��عh�n-h���-U���ֵ��eI�'j�s7Dm��n�D8t���=�U��wm�%�^�˫�N����,�ff���#�������T={��5*���rg�Z�p����0��g_�TH �H�ᡷ����gɔ���|��ۡB��Ƚ]��PYU���|�AuU�hN�.`��=�n޹�}��W��*и3G���.��;M�J��!�2�կ;����Z���,�4�3Y�+��A6AW}5Z*�Ng!Kdғ�n��˗���e*2p9�n��H���'(�v�e�W����k����<���N�Ne��Ϸ���չ@�e�H"�wH6�;��Ձh"3���������/�E�ș�b_�XX���~��ei~	��}hji���6&g�T�G�M%��Ɲ���,���E���8�j9U1Y>�_���N����PSU��&��uܸ����Z��t�y�y���r�1==��@9�ܹ�$O{�>�P`�����1���T��æK���$Ώ����Uw��=����Ǔ�������tj���Zu���?���	H)v�����W�	%&�P}3F��Ψ2V��o��	���"��K�vዊZ
���C��8�G�? UA��:��o������͘Z[S#�����e�bdO��h:�;�wʂ�������e��	��vZ�$�0�5f^އ9y��HxN!���NB�ũI�fj"�b���A�^/��>��Ҥ�B�͞�f+y��)(E�!�	��h抒G;_Mw�;gQ�.��EҰT�4��*)�rmKL1���e�MP5�\KG7���W����@Gs�
:�v�<���OU�s-�<Af (��E�e���^�$�k�*���cnv
N��LY6�l�8�*�ܛ�\�~����[w�B��_�ɟ�ݗ+[�;<��f@�������E�����D�y�F�WW���)e���m���agoWc
oY��r<��Ҿ���������x�'2���ӎ�^���H��x��y��@�H�V��%������?�M� .|�V:.��^�Jw,�C����%h���Np��!�hmW_gXG��a�Ɋ��R�<0���e%ɝ1j斖q:�.I[+�X�}������:(����!;���8��F�<<$72��v��z��;w�T∜��T*�Rp�{|��"�ל�]�J�
n/�؜6ax�����5PEЯN���;Bz��}Cm�F7���?�YUPp����\�
�.F��B#�D4�J���V����JA�U���"�w%,S_G��(�+��m����@%���p&t[!���y�~�9���1��}��	��C &���e�ܾ�`E@�����9��9���\��Q]
��k�j�a%]VY���}l���Vg�O�d��wjEw+��H�km�x�,�m��kD�$��b��
}\DP�u����^���<�_9n���<[�/_ѹ�t�+	�8혙�V��+���=,C�a�`mc�|J�������"�_�%��.P'\J��c7��9qA9a�t-���t"�ɋ�γx�'v '+�֮��뢛W%��Y�͢opH�4"҉m�@S��p0TI�����t�r���W^[S��p;{�t� ��BJX�9��ۤ<93=����|
���]�=Bw��'
�����܊/>�Rϛ�l�y����駟�����~|��}�QTV�I�q����F�i�+��;t�}�8G�Kad����0�1�!��u2j��I���A�*�}�Z���+�׌���\���!�͜�H�3���0FDl��W�'?��� �7
��R_���F#}��k�����5�X��ה���Z����X]:;t>;69�4����$����3��ڷs���?gB7%�Z�����ik�7ȶט�@@O_���NU���QK�B��뎢��]�M��<���mo���sc�u��ؽ�Yr]Y��Ԅ�9~a�H��H�]0.���*�S�#��cC�ZA�J�M��M/.���m�k7��ܠ�D�0����]�#�PcJ՝��;���"k4�a�@�nE�W��k�DO��W�!�N"����&�7��Ƶ?��t��'�=[��_��� ��\�ܼg΄�=�ص+�\�9��n��%��064���n$D2�07?���]�݄� ��&)wm�o�2�
�c<�;��b��@4�'����6r��(Ր�����C���R2���G@T�⃊'�����!��]�uc}uQ�-���1��jnm��e0;�^(��
vc�zL�Lvܝ3Ry��&�����������&f'>C�`E(w��`B��CԵ��"�A.�C:�ݛoad��L
�l�[똞���e	ˢ��mmMr|�E����]s�K`E4F�v��q���p֔��֦fW�,�>}���+Iϯ�?��Hf~f��x܈�G0viHf��H]���m�������\T��\۔��d��崦,X���5ux��&P�����j�,N��`2�V�;�8?���_�s�@�:\0{*��:��	�"*��A�T�
��x9���5��w/p_B}C�{�8W��P_��������cڕ�2	X̜�S����E$ҟ����A��W�����>P2x��r�钦���ؐ���Z�`O�&�Ħ�W�<���}uuukJDp�X���P�c!Ʉ���	�]��cqq	��Jy���s�Xo��|g}+��a˅Q�})�����w*���&]��R�f�@%&:���hX&*�L2����iu������2B�8�z{��f� V���w]�/T$� kL�H���$��{FKk;&^Oa��D��^A�]eJMy�����wڅ�!ր����F����V�@j-ba�����bhhD��:�"�9'�1���K����qtUa9?�}y���c��@���t�_AK���,G�$ç� hU�dB��=DP�hF�������x��Xg�&g���ƄNЩ�'%�"�Z��➘S&&&v||�Z3z}U}���,�c~~V��c~&Fv����l?z�P������z��vz~ܼySy~��� ~��_��r��5�F�XX^�����Q���C�ܭ�(�*�m��|�iD�%j�7
��	�F�朰���`�ËdQĪ�܇l<���V�U1?7��l�{�Oʣ����I ��7e܎��(��g�E��IY�:d����ۃS)6�NS6�(?GUePxv5��%�Z;���QSQ���w�%�sx���B�$�.�j	ǻAt��E��ge��q�P^�C��)a6�5���-��q�xT�ˣ���ݺ��v��w賅�������'/�7���;P��V�G��Ã�?�������"����1N��89�������چ��zQ�٩���֡�kn�y�B�D&H	���|��ν���!�O:��A��pT�����3�/~���֌L&���l��(�p�������ӱ�8���PeU��t��A�ߣ������������K�i�vadv�o���0��Ԡ1��Q&�����?���hke��p~���+R�<R&.��#Դt#AhV��$n^����&��];�����Ҳ�g�u��=�v��h?t"̞����S�x�V�Sժt�	�P�3��*�D����]�@��� �S3���{*b^O͊�1`Y�K� [W���ƚ:46թS�&t,���L��D���� }q��� 1V�L
Q�*P�{+�x$&���HB�S�ē��:��_>�͛��p�a�V)�׷(�{,v�\�1���:+TŚ�]Qq�dm��q9�F�ޭ�'M�����<�N�~�n1���e���B2��M_o��;\�8P�5���������	�,v�I���.r؁�EH�yA������d�9��ʊj������H���O�&������ޟ:��~��	�h�ōeq[�n�����<&��C'ʝ	��@u�����w���/�(f3�{�=��H3�3Bh�'A<	��s<t=�i���H���z�|���U\װ�d��̎�_k6z:���j�ϯ�o -m���#Q!�R�q�O�`!�ǉ��9��{�!p���Ǣa]�vEw��.�4�������wf����cwN<8��a{�'g1��\6�����_�@,|�	M�`���m}h�B��l���1n_AM�Rr�sˋ�2�3`�pe�u�@sd�DC�ƺqq	�����əy������jQ��Lpo�ݦ!D��Ґƭ���^�v��?8�������h�d�>�k�Y�i����)_&���v��ǧz��0���\˾�M��ܱ?{�#����ǫ�,����0���a���X�|g>�L*��`'m�	�-�Љݰ�v���f������[\�R�(!���e.Z�QH�P]Y��@yV_y%�1��K�x%m9`�i�C�@���"�99�#�9�b�,G&���25+����io1��t��X���3Db4_���;p;5��P7�z�v���wp����j����O�r��_���K�������|~�p��cr�e.��$�p �f�0�7�y�v	}�Pp����_��������{��[ܹ2�:�����oQUQ��C<5%u8rO�Br�"`kt�_�=�
�n��f�E��������I����W㰍���f�Iiӝ��;��r?:��PUШ�ų(����/�ĵk7$�q��#�\n� ܏��������^.���PU]�gϟ��<d��0WT��׿�L4&���1%TJc�d|rr���V���cfqV������:�_~���6\����e2#k��C6�#Aκ׋�Ewo�Pp�>��r`y}/'����(�2G�g�0vtu��u�2}�Z��(
�uSV�,�)���&�u��,���ꊞ}4���W�084�`e5��W�R8]>�] ���ȧ`��jF�����u��������pzx�N���B��?P�N`em]��<�N�ZL
n����&�--���J�>6���5�?�5,yr�i��T��=tum�J�.&�L�o^w��cu���k�W��tc�p���7����v��٩
��&2�lCyyN�w`3�Qp���յ5hk�����_��Ȑ���_=ƍ[�d?�Z��,���S�\9ԗ{�u��d�󱓻}t,���!N�=WI��tV����5���p��%��g?Z��Q"r	
�|�*�V簱�.4
z�/b����Z�d�J�;t*�\�E� ��3)=Yd�|�C�R�ZX^�"�!?�;7F�ӓ�졲����X\Y���~/���h��v4G4mY#�َ��h´��_��q���u�6�&��H�G��&xn�	e^:���6�H���,J�jk��Ѧ�J����ɴ��������{4�"ː�����Bop{+4�'�q}y
��?��]i"����־�s�%� �}�����N��t`~eI|}���Q�ﵷ�GkbU8��~;�L����$���֮�W�8M�����(��K,�_u\%�=}�W�]�������e<�q0�W"�9>��GK}k+qr|��S���I�ziyg���8�`q��SG�x(,:2�0v����j�Q(Cye�wN�a�N$���_���ԡ�r��Y������{�y�5^�H�&Je�
�wѝ�ݫ�WJ\{�}h�� 2q2!�����/?�mݨ����܂&Z����^��I�ye������l6����.�J���A��{\QR�V@�l�]m���H|)"�WV����ޝ{��vU�&~��*���F\����uu��j���O�ⱷo Ss��?��E{{a�μ��gG��$mq�R�lp����|���?��H���ء
������[:���)��Ǫ�roz�������F��bfaV����ɒ�����>T��:�|�T�Z������>�&�ƇD��|1�Ƥ���A�%G%��&��
R3#��nG+G��Uh��j<���)l�������z���̺�F����Y$�����Ȥ@ʊ���9X&>/�!9m`gD�qr-����䠖H	��Ѡs}�G�k�R:;9E}}޾�v�ӯT�W���2��W��I�2}1[��y1v���l�PB�֞)��ի����*�n�?������{�@Y��z�t!#�f P%�W*SP�`g�J�[�`���9)�t�">���:�=~�����[��g�����@�<G$���v��jy��u�˨&e�cc{C*N|Vm�����+�S"-�Ѽf����o:�-�?����!ɛ�I��ǿ��Z}��*ʽB��>4��<U���O5�+�=r��L��`    IDAT�y��6��!ܽ{C��{;�fG��j���,��+ ����^��b���!C ��!g����dɥ��ڀ��^ѷ�n&'�0��L�n]�$D���1~�{G���O?��%U�L���9�8=����>�u�S% ���Q�ł�����Sp`�$�D�Q69���׏%)K�"���Z)ʍO�cm}�UJ�k���X|[.��Ή���������焋I<{����e�K>�j�$�̜���9��I�����p�؏\�3,�V�V2�&8�ד'O�"8��O�5�qtN�u��Ra�;��N�#K�]�*xZZ����k,,.
'Apw��]�|�G'� T�,�����Cq� bKQ���LN������:��Ql��be�:t��Z��������>^��$.u���Ј�.U���j�5\^zg��v��QB�1��ɂ���i�Lgҹt;\8=�+�U�ѽ�mt�����-M��,����3���F�����<�@���$y��N%�J�MuUڟ;��To{gO��0iB�b��p�!g����]���b����8�,��v,�p4��Ʌ�4�)��}��n�d����P�ԋ��C'�cns>�룽�ּ�[B�`��鹦t4�8���
��j��nQ#��Ӈ�PXL���d��(A��Z�ʥ6J�'���}<��Y[��?����1&��Q0��A
��dB��2�\j�4Y]]�@0��P���klIQ�:'��������9�Ml	�#���w��,%`�k��u�����Xa����
�n��E]�|5�?�v�?�m#w&�������|�o�f������ۗ/���QG����\�؉D<��㐺6&t�����
dzf�;�y�6��,/S�N�c!9Y��KU����e���-���҂�nT\�������mo�pV�T�潷1�� A���A<|�5ַw�l��GLtE�H
:�Kƣp��.�/&�/Sg%*�ݩ�G0��������AP�'�������3��y%Ѓ�e�L�G�t�9��$�Kw>2:; �wr&ܺ<��2x�n��^MO����[B�JS=����_!�9�s�7��\�����Ѭ��<ķ��a��U�'�%�/�+�ooI����44����~� ��QQؘ��f�z6�BSc-z��qzr�U����\G	Jщ�v!�#Q)����P�߽Y��7��p�#Cڧz.�+�Lgp5t���s�C�x��/�$tr�١��^WB�@G�Í�E�o_U��.���ر�w(iQvpN�M�r�:�(ڽ�4���v7�9�{sZ
�lk ��ʁ��u,,�kZ�N��m�[7o����h��g[�p������D�����i8I�u�1:|��	��PW�B���,0#ј{(��������2��{���q�0�����+2���C�yI�ZB�R���wm�W�V���)z;�p�Ұ&1�e������K�}������SB�H?y�>��T�d�G������09�L��d��u���Iʃ���ݾv�:>����8�z�&�����l�d&vĤ^�����63<v�bYe�BgSP�4�	����?Dd+%�ϙ酢9ˠ3���ص11ݺ~k��x�zNc�B>���i��c��ؙ$�D��M4	lt����ՋKTM#%)�C�4Î�.�ѹV��#H��hR���V�6p���b.�U�0��]���N^``��2��r����������AyU��[4�D���㜢g�q��V�#gRQ�����m9�QpgucS46�����lkGks���~�\q�SP�;N+�����)bh8:�Y�D8�͚�Ǟ�����y�n$��0Y�H�lh칤���B���$z[jpilG�(L67��U�8W6\��6գ��
���0[��`x�A�v.̯ r3D�� G` ��n%�H3-/('ut�css]��77�195HZV���iA��|�}=�
S�:�	�H=�y�βT��u�Bg8��]����	�ۜr�2\QQ�B�9�<�#1 9�aX@0�����Y\���� N�Yj�a��{�K�4K�\�ox���>+�uM��i�F����F�EBH ���V#v��E찳��e5�0m����EfDf�ｷ7��ιY���N�U��Y�7��~��<�9&�+J����h�'�����:�\����w��w���e�h�9�	ԕ�����bquE�]�#�<�!��2�T}=����9����A�=������֡�~;��漢j��|-��?���:`R���X�e^WU���V8,F�NN��ģa�����3M��PT�_~�:^wA�.o��w6�&�����Ǒ��Q�C���%JK���֮�K���ř�;"�.���� D�Q\_�d�i���-N�n,`g�"WG*��H����������Bu�Mf����DY�uM���{'���f���y1��e����w�P�Jm%U�y��py�xH���cG�ˁ��w���Ɋz���w�q�on�������f�uN��'��kc��")e[Y!		Q'G���n��TH#K/on���U���m(Ю�;Ӊ�y�ae+���dws_��`Z&.,蝃wP�ЅX<[� s��}�9c���;���	�P\R���b��H"lo������OiM
$��/�\:�Հʲ�w4�<�;?�����[�����`w���3�b�z��>?LN/�`"�<�4�zZ�v�_]�t�,n�{��/_����}�N�O�.��[qQ)�[[dx��%��6��*��"����|1�3�2! ���{�qsq�VM��tB�Eo��P�{wǐJ��(�������d���6���I��x�J;qNP�%rRxpE��e�:uYq��NcmJ�,X\X���;�O\m=��g'Ǹ8?Ɲ�����Α�8I��E-C��R��$Fq��no�P�?n^��9���D4�$C���&���M���7o'��'&y*��w�����ڎPA!�����W0�oK�A�2�y���v�S�&7�b����]�"�N	A#�O$[>�@S��������hD��F"bN�3 ���U�ch���7���͉C1::����h��Biu������
z2�O�'���*-t���Q6����N�{p���R24>��ق��s�܉$i����/�"t��=���?0���,,-��ԋh�;KS�X��)A�+�`��}��&��э˛��,�ў&t��#K��g��Dvl�&	��d߭.}���I�,�(�zniuv�3���ae(�ͬ��k:���"}r�RX����
��v�wt|��yY5�q��:������D8*++pvq!�KH���Bm]�N}"����BwFH�k�zV�Yﱼ7
�(�D��p�B��<?����+q�l3�H���|Aw�M�)p��x觿�
���M������S3b4��q"�G!C(��<1�fBkG��2��fț����'��)=1z�:=�����SF���ī��hm�>����kr8�IG4�����[���'�{�ۅ�*퀩�f���·V{5uu��;@cSv�����kJ�n�����r����=X���̗���UD�Ņ%�6[�;0=5��O؉.J��yi	5��iRcZJ/�hLl�x,���bDS���pX]8�_��ҳaA~�C�շ �L�Q��x04���*����Z��N�=��}L%�/����M�oj��ck{Or/e,3#E"�Y��T"��*Â��
4�V���/_�@>x� ނ"��_���(W7��
G�t�(s�bny]����h���Wr-��ܙ��7�V����"k��΢E�MO^�y#�,v��b:G�@��[Bf���b��qXLY�Џw�D����+2�]����*��ئ�i6�޽!���"\n4bvf����Bf4�����ݸ36���3Lͼ���)�%�r�3Z��gA���hQV���$ч�߇��9\�
+�r�����_��#���$�Q����]m(pZ�`aNghhi��ѡ&��.��\��I2��$J��U+�2�ǣ�t����`~�w���e�Jf���&6��`����M����̈́�\����S���/��a��+�4����I\��VV���8:�G�ֵ��Dbi�)X�r$�(!s{�^dS9��}�Ņ9]�z{�QVR���q������H��٣�4�BWe�
]6t�6�w�U4����
�|W*:�hg��MA���	�r7΂_UU�����7Ǆ��W�X��A�~��v曫�X��
�TV#�,09�00��Ս��3�����C���S "����0:�:q��]����ʪ�*j�Dt��ڒW��Mg5d��4���	Օ��E��>������РI��種�GCs3&�����Z1֌fΆ�N�U�E(.t���{;ۺר���?F[G��ة���&w��Yȿ�&:���U�`U�>��:�ֶNlퟫ�W�~[��'�-�\a��N�w����� �B��?g!<�DE�[�y ,�W�7������Q"G��ww��%�>>8<���B+�j�1�2���Ռʊr�x���lW��y,�l��t}��"�bbz�,�C5W2�WA�!���ؓυgvF����!���2�LB7���GH�������;ʮ�ܹ#9*�>!cT�8\x7��S�vTT�!!³��ܹ������;�J=�����~����_�w����S�a�hr�K8��*dVwZ���m()�G�C���J��z��PV\��ʗ��_�Q=$��!��+J$��c�:Ė׷`�ڑ5�O�Df��@KM���	u�wF�PY����V���M�32D����H��n��=����#��߃۷_En�U��m1�dmu]yԍ�b�r�D0lx��R��O"�^͠�i��_�%R��9��h�Mpy���������{y�͋�ǿ���VD�U������~4���a5!����؛��j��>�ß�����ކ��N�bi1��ַ�Qք4�ڌ�tXEIrg������B!h�k�K���U�XEUGn�؅��d*'�)
���:w�#�b���iY=%e�ܶ76QR\���Zu�쮝n� �g�^��ʂN)/SN����0=5�dάx��	��f��n���_��'�Wt��\��{$���.g�>���&�����E4��� ,v+l��3�T����9;N�����	��%�$iٕw�2202
o �߻��Q�r�~�^�s�hk��G=����.�p��L���FCװ���픾��
	�3K8��@U]-��w02<,�;'\�C�Y��/J���ǂ����h��׿z��ivY�-�P�	�`{�&��ؕRA��I����{�B����7�~��G�-������E}C�3zzS��O�{�FE�L�q0q�̀��VTp�g2���ہ�������"�	�����tubz�%�:�p�`r~����Q�ܡ�Ԕ�pzx�d<����6��ˋ���V������ryto��v�����y���5.bVgI5��F�`�2w���K����lv+�7&�����
�k���dY�owub���TJS!����y��D�Hd�&Ҙ��i�� ��_��PN]4��U�"f�|9*���.a67Vp����e%�x������N�?4���m�l� k�#�e�k�F$�ME��R���j!�V{޼hmm;;��r����UQ����=��	S������
�B:(_���#@~�pZRX�|�����y�$�9d�n�5����?��^(�|�K�x��i�R����oqqu�?�L�\0��n~qYJM�d�g�W�"��	`&����(o�\Q^��3r�|�W8�?P�mkiEUu�={���A8

�pĒI$35��8όH�M5U�:l��,�y!:D��/ѹ*+,FmM��x��2Hf+�&�Z�2���WV��b�B<��[��0[ͨ�*E$r��U�;)�d���PRZ.䓵���h����?����ׇ����7���0���9�
�!���;�4��h���hl�B<����E.�&���z����n����	B��|19�
M�uhikU�CHvb���l%r:�67�F�p�c�<�WaA'��h�T8,�*F������K*lL��nO��:a�PLX�jBkC-�������ٹyi�	�TU֩��%�f�m0����u�μ�LYf���E�2gx��g�}���8ژ�+����?ByC�
:#,�.���B{m��Hlno�p�#'��B�"��_�L�����c�V7w�m&��ds	>��GS�o�md�&��hml���lV#�7����K!w<���%,����2�%�S�UȐ��Q��Xt��T�iI�-t~���K�J����ӫ��5I_Js�_7j0���2���GT�#��4�e�N�/Lbe��_)����T�Ñ�v'��@UYѷ}jrJ�+>�XŐ��`$����.g**�Ꮕ��ӗ8&@1Z�\z�hy�����dTA`� !��.�M������B6���mx�z˛��Z�H��fG��9�ΆJD�W�/�-~y����6vw�b����s!���NA+>��W��1#���NK����*����Z~��A,���P�{ku;k3�#C&�mAo�/�;'t1o�����d���a���>��_���5�������XY]�o��gjL8q���������Nk�<�EC��:�ۛ��� 3>F�^^^��������q��������S�*�dȇ��b��W8����&Z�Ӌ��.|��k�X	C�B%Dt���[�����i<������H���n�����єA{w�͌��̾�̈�,~S��}
wq%b�����@K3Fo��@�)��kz��%��|K+�095�}�Ï>���5����Ꮢ?rU�\�a��uF�KϢt��0s9����ť9!��=����/��Ս��+��Yd�뮥� �y�.3���L�z�U��l����O�_h7^\Z�&�u�g�faCD��+ף$cR�ƒHbLV����XЗ�^`q�9�Ƅ�}�,��rִ��~�K:r� �3q�����*��i��s���?8
ϲ̓ ���o�wi����g��Xa��'�N�!���ꠅw�� ���~�+�o�h�`�v�l�Wd.��ֆ/�=�M$��Ά����)���m���y�=��6���5ee�O&����{\W�5��D	Y��J��S���)����!N�/`��PX�ٔ���	�K ����tc��.W�)�ԗy_��ÿ񽞦_�C_K��?����I$���F��sQ8��pL��SVa*�`6�8�������B(�(yN.���%��?v�l'���\׀��6��aM^s���;>G�d���v9���k6�r����1f�Gce9��.d�B=���*�-��܃,wN���!ɤ��CP���)��zqy}�چl��i�ojiEyY���`X����:M�[[��2Ȕ����1Y�|	�\��E�n��#'"�y�,=G��X;t�UȂ�Xp��o����H~I�����@?����t��)�[YV�!͈@&X����6y;���;XZ�A6�&2�݌�"�i4�3�Ο���ou���
A@d;��of�a��Dϟ:u���Dp���TǌUo�p��(|��;�{�:=a���������+�dx�gD�
9����;^T�-JڸǦ��l�Ƅ���'��������,蕍]�����c�V;*K
`��b���"�&j]�N}$��_`hhՕ5��ɘ]^���%�f�|d�C��\Z^$�|�:��cFvmyZ��T_���Қ�/�A�
�&�L��9��`�O	r��t2����{E�������G2� �s�3�����D4�D0��Y����'{���!_X��P"��Ek�r8�\����S*���gR]SW~B�]��j8�3wgtPg.��}B�4�m)	cr'��MY'}�m$�X013��� ±�̜`�E%w���%7+
*cV�=��8��Li��LDă�d����$sD�y�T6��?O�+񢻽]���(t��GX��5!O6;��)<?���Y���x�c6��$�L    IDAT_��a||R{�¢2��FE�ҹ��`+��	�鳓�bv������U\���]M��--��"���/羼�V_~@㬒
LL� ��6�^��J��ʤg�Ϣd�f��	��`�U�q���G�'���5����Y2���[��x5���)�I��*�Cq�]�DbIF��b�P:�� ���<�q�P�b���M�����xW��^T7t�w���aw ���"�?���<V߽�=E.�PAwz+`/�����]d,�|�$�hHa���-����TK�k��ݠ�o5��҇�����$���%���g���V���5@9�IQ��V���Y�%�lP���4���3zW�������˯��u(���V����9xm6:ir$�hL�U0�ƭ��ZrLYC�q�5�j�ěI��<w�n�w��,��h8,N�
/.b�[�ܕ���n�n&9 4@˿YH���_|� ��Lf�-��:_�p��?�M����P��/��?�N��H:g��bM���DP�p�!�ā�{��������2hn�E}u̖��������y�@�.�wR����s�tu���\d%�m`k�T����!��D �لL:�d�6zf� *E,S\!]�jʐ�����Bqf	[�B��Q�I{^�uiZ�����7�������;�y�S��}$;���7�Py�S�Z]U!���H49;����\%��dw��/��9����	9{n�#�J��N&�E���AKc2�
�v��|��?Q�6��B��z��hn��Q��v��1���D�j��:Lr�ӡ=:�wZ���v�4V_Y���Z�����{�z;��ڟK�A�<�S�+Mq����<?V��i��'I̽!'�f|�7Jsh�v>��Y���ҲMk'�`dL<�E<�x܅үfA.��0���2j�L���ފ��9O���{�<F�'��L��e���C��h�]�?��!��CV�ff��1�r�� OPbl�)��4M�b#0k�!��JA�P��H�֜r���q����X�`u��ĩ͐����
�F��f8��c�}�S�ң��I��}'d��|�L�ca|�1���TUV&�����ǧzv,�cY�)�aocN^�v]S0ZJ��� ����cr��E�����+?�1!��^M(d�f��EҖ��W�Ø�	��6vO���<©�T�Ny����l�H��w�p%��d�Si��ބ��C9C�K�(�o�fd�*=S.����T���9�������N���?�Gye���X��n�}~}���MM�,R��prW�cy)F�d�sus���s�܅"��}9;����$�ק2���]P��;(�i�iVdL&0�܎[-�
�af��ɹ����5�r\Z��X���Qc~����U�F��I(T(XF��b��x\L��e��3��b}u�������ߗ�}ffQ�P6Go3�gA�GCmU�n�i>��k�R�<E%�}Q:Iu %�t�$�M�+6�l&y�Q��������9�NO姐��etq �+o�67g�6�m0XPPՊ'���4�$�Q��u�p��եH%R��Z�9�[������W����T��W/^#�ex��J�8����n�j��ݻ(��������E��u�qpx����n�b���H\lr�7rY�>u���� k�,�Lw?QA�\_��$�!L��FI9fT�7�
`�`_(�ֵ$:Z�BcK����eznF���x�(+� ���d���Ǹ�����t�g_|�D2�J�������oԡ��W���O����߹�&��h^�UlNF�RI���RN<�&s��"��d]m�0���d�a?�{�ed�BHvz�-����\�X*,����k�b�2��3f�(Qp1!�t&�pد���eC6AqQ!ƆF�N|�f7���fH��@UE2+�.���g���-�=�|Ado��G���Z�Q���ڸ����
B��k������acgW��T�ڌ6�o/b�%��c8��5����uc����YR+V/s�Kى������h ���x5��xw<D*�T$i8����H������H"[��^�D����/5�A�.�B�4/8~���)	����U�p`u}�W~���X��&#��J�_�����)�NUu5�f��ܷQ��Їd"���z�i��Nkbb��ڨ���j���)ȇD���+l���塃[�t{��X�{�,sI�rA/o�A���8>}xG N�|!_�|)D��;*&<S�@�^Nʩ���L����6�n��1͍��̒��>����$�V{̠'�����pL2/^ �'��'��[�bQx�.X���ޛS��䮨���Ξ�Mܝ*4U� /�H<�g����*��t�wq�4�'V��>U�uʜ_Z��e�.p�j�Ja��0	k6 ᛂ�����/M�$�1g3h�*�cC�aqb#d8==�x`z��!kiy�� �F�����]!��O_��)�M4)�@޺�{�$��w�q����^�W�btt�d9�Y�z�L�l�6���#~|����m�X[�DUe�R~�˟a`pPꔵ�u�.�|����AR=���$���|n�U������3.�-�+��$�6�2�T^D㲰�ST�mAOЛ�Y2���vv��ec�W{��������cJ�"{�q��'&�>>�3(�f$������� v�N;♄�Q�g�@��(��G	a2�̸=2����3�����P3�����JC�J�-���˚�n���1�Z���8�p{03;�����-�y� ����5�Q�ˉ���9+�a��[ĥ8=��	$��sal,����S8��Φ�Jf��VZۉ{}�卸�a��P�ވ��"$)���y�F��'�b���u����!������5"��B������*�A�	��
�Y��ˈ����d�TYU��;w���Vw�a��%9���j4�M��޻�յ�nf�Y�{'����B�˂�C���Q�Z��o{[�P�j��ҹ'B�Ŋ�2���ain�W()�G$���9ql��	A�Y����@E}��������!�*�k�{���î�]��#p��5}��o���g7Y�[7�����"��hL�"$�q'��މO!.�o`��$+p��܀��Z��Ti���ߓl�:���m�e�E��{���rtv���w���
�n`~iSz�"��$x��`H3:π�FT�V� �}������S8,�����82f��y�4ʊ�Q����p_ݥ��=N���/��RR@�QB��!,̗�ݳ9!�˜P����"ᐬ�:{�t���	�cA1bj�+��#vs��.�,���·?VA���9�n��Mg:�GOC�2uO�/���0$s�ڜ�G�*��ݒ��RQyyo\���6FҔ`�8~�N��PS���R�9���齅��H��8>:@yY�.m���Fԁp;/cBDT�,-Fks=��6�Cm(ճ����B6:�MY���TI]�D
��hok���b��G�(/.Aeu���^OO�#\[�4*-lyf�D��Ɣ}3��/�v�dx8ҏ���AxΈ�Bxtw�}^�U1��^���YWY*�9�� ϯ��dw�F�sfA
�DC�T���ݽ]y3�l��B� ��L�I~|ֹ���p"��Nx�ܒl"�Φ*�v�(�������T�<�:��Y<wlJ)�����L���-���.6 7>5f��Kd��}���5����������R�aA�IFů�F�h�(��ۃ�H��K5Y�̼�����x-�[\��أ���
�|��L�.��&��ъt����DcR����f�� �K�%Y~�V�:��a�ٰp��9��v�JDi7+����^��Ŕ��*�aqy�������ںB^��wBH��m���g3�\_��~y~*������,��%�8����>��^#pu�<lp�'���&����؆��.5Q��ή�f�-�EUE���Y���N)S��H�~_�dƹ?��S+H��gԐ����i�l"���EQM`Dk{k+z��`���h���>�旵�"��Ƅ��wSq�Kde�Ƒ���VQ]���r��ۏPRZ&�`�o�ٻ�og��7�����X.��k�6;��cB��'�4�.cJ�ZSGSfT6��w���/����6��#�hk�F.�VA�>��:�Ϗ+/6#\�LM��.)�d�M4�Wogq�HV(9�r �%���Z�ۆH��[���U�ags[���}���zj{�H�P�oR��x�B�]N�Te�����,f�e�`ay�K+�R_73�CXZ_C�?7-�9�U׈���nA9��p9�2Ժ�>�������װ����5Դ����Itwv������������QG��_[�箢5�����e-�6��De���2�q{p�Ņ�������'*�4IG#�~��4��n	����k04<���R&le��y��5UhiiB(z���R,�ncfq�f\g�v����/O��ڊ��6M�ggp8��6��!���>�R�"ނb���
�l��hF�҇'��������E��%�LM���B����p'�d���LF~Ȝf�)��8��1~���QdR�X�r)�u���g_�Õ��/�@�Y�	��4˅�t�f�hB�-,���*�/��>�&�~��`_=}���^�גQn��+[r�cA�lm`�u�P ���Rш���$9��;[8<>G�H������HpS�A:���*�7���Ņ^��*����"D�â��%��s�ʳ���ц�B�d#�H�K�zQ����҉7��!
z0`����Y��1��h��|��7���6��I���c��G/?/���y86*	
w�,��'�`�����Y��n�~����SX���� hp�!��u@�,V�O�������P]���3.��m0���3;�B�=����٨�n����0[�HX\_W�Hqq�H7�b#�)T3E&>5��~�$eϿ�J	d�Т���:{��}$NC:����ake�\P=�H������7I&�Y�[_^���*��8������@/*+J��FKѹ�e\^�����n,n�aneW�y,0l�l��9=ȓj6�� �pv|�U	^ޢrԷ�(����
6�K4!w���l��mݝmj�7vPYQ�tֈ}�"6ج�K�j-�\l�4�"I�bn��qIvw�=DN�y����I_��>H%���Z���x�XF�����9��>yPzsG~�����_����[<FMU�Ѹ>:���4�I���G1�nQr^��8|C(��a2�k�)�ٲH�B�I1Y��L(r�02|[ϛ�����G:��&�'YЍ��F��a2�tkG�d�Kk(𖡩�E�g秸=2*� ��>>o��TW�j���Vv�V�6��P'��&ȝ}}�H ����"����7u����PTR�\2��m�.�����p����Wو��7��*����Y}?�ap][�j���d�ԏ3�����{u"\���c7���8��ш¨���[^�����,Tl�e���h��;?C*rq����J���O�ܿ����v�����%�F>Cr6x}��@DY #_��Ȼ2��,T�4�:�*˼(*����˟c�� ��B��Y�U;��©�����Fz��ڂ����������Y���L����>�� m��b��1Y�(������ڵZrY������^��虩Y�1�SX��?�ׯ_���Y�l�^/�7������]zG#�����Û��Ļ�Y�Y,
��)pKz��ddCW���.rS��F��i�ɴ�P�0�z�L�\GG;
�^,/,jo.+���&I�dHr��!��$��88�Ӂ�^$	I�SYݠc ���3d�8�Y���+�w$[S�0���=�,��Д�c�Vn�jC:�;���l���?��Hfo��3굯�O�_�4�&Y�OUг6����ca��~�S(&�ɜ�`��GyA=z�ٹ%�Xb�!�I��ewI? ^"�N�A���П=v�.(��}7��EJ�m��ID��(��R|-Me�����ỾP6��`DK[*k�brR�]2=ˋ\�����*����Ņ�#>EA}�9�0�"���Z<�7�g�Ɖ2�_-�/^��gCEI�sy0>����3m]��C�!lY]V�,��w���Y�ݑ'�P�	u�D��ל9Ϻ����a��d����3!>�C�(��×/^ F�n�(ɗ�`�.op:���������d.�|X��k�$S�������ڤ�Z����^"��itS��G��PAg�9�Ae�?E*�w��C݋W�E]u�
���*Nή�ɓ`EV���ъ��3�
�%=d3�F�r)�dS,t)���]���.��hkk�_X�Q~��-�)�#m�g$\�02ҋp�&#�D/N��sk/''a�K���g����jR��Z���]�ln �L(����'O�`�� ��{:7�_���N��T8o�c��YX���������K�0��)�;�����rxgD��SY����huł�P�`��u �k�R�x\B����� �OJjWU]��Ϋ�3�/-���
�eUR�d%#� �`gJ�X�V#
�v5C�秚�;{�U4��Oa��UXXY��^�-n��d�0�{��A���DEi��wN��u���S#ɂn1�TЗg�Þ�����=kr����=��֋ k��#����0e�����Ɇ���@i�K�["O_�����Uk_�� ����[@�h ��4���ߜ�9U��A�J.%��G)	��HEE9��$���iB��!�v�u�e�=؇H0�������� �mY�ݹ� &���Gy���G4?
j����ޜ�;F��` Í�C��P�q���
�E.8]&�o,`qc	F[##�����6eE�߹=HR��-�/O|���Gʙ~/���Տu�B_{;gf�"˝u_W?��A�\�Djc�xWK�+������9�mlhV1�x�?���yB�\6��8�/�mvϐ���H�½zsS�X��X��U�yK�ѱl��� �G���ί(�F�h�Gm���c~��*����.���;��qzt,�8�|dr�.�*a(~)�&�;Z��ޖ���)M���ё�`���_o�&ty�����9ބːo8��e��3��q�<8�YT�ᓏh�m�E�4?�x.-��\<���T����d�J�CmV������	�;tzC�;��o��;(�8�p��@|i���6k�!���x6>�ˋ�It��Â�b�׭�S7\��i?TY� ��p��Bi��ߒ_��IQ�dJ��s�g(p��/g�M�015��!�Mpٲx���p��@�Ml��������162�hJ��=����u��iJ��R/'&124��86&߭bq�LE�盐{2r���'��@������wu��n�V�~�p4!��YYe^�I����,V�%N�$�y�M[d"B������&�\��ݱB��4!�f�x���I���
�eH2�b�w@V0	M�x�L/*���č��cl.��xwY�,��df[�
�7:�%�C�݆�~x�dX����!f߽�,m79a�Ntai'�����C�9��t�?}�
���ǥ�Ѕ��m�M�߿�u�i��s��.-Bks366�ffF�)r^x�q�J��b� x�ft���3Y��� M��`amS)���Ɍm}��"ٞ2�f�zZ[1�敞�!�����nx��.�@6���,O}��Ց�_0X���� �o
:��κ&�D"�����L����nk](?o&��j�>6L#����;��]�/C���d���K^4��Î�V��������d~�G���Y�M��!tHM)��������:1��P�!��n"B3���zJ�@"�J�*I�0ӦI��nSSS���H�(/�@cK+��δZ���7��1��sM�`�#��[;�;p����di6�O�����!kjc���.z��S��bl2?���-tz�Sqp�ë�wj��L��a~n���&"��ţ�$���G~���l����v���I�nR�(,� ��V���~�tuau{K�WU.=    IDAT�J�#g���Z�������$#�t������L2%'˭�C�p�TS�xsu�ã-Dc7p�3 I�F�S�ȉ,ʋf�s����QO����_��4����;l0�n$�1��)��5����7�TH�7���ƭ�~	��������!�gO�H&����@oe��g_��b�*��[X��CJ��v�$�D �FC]���pzr(����Cu��$+�C8:9��~"i��ʺ�_Bd�rB7��M��!0�YD�z�I�aZ^�,�<4lF�j�Х��#�p5ٌ���zRG�$PK>��z���E\���dn#b����[���+���gz:�������)�V�;˂n`A������GiI��@ڈ��	�H�]�t���B��bg}�&�����X^[���>��cD�A�l~���斖��{����h�jBbD#t۽��X`6Q瞖��id<���{�d���ĝT:OR�r8�b{\6tBƱHDY�΂��Z�Âb���<���[u��t*F~Gz4AH߂\"�͈6\җ��)K(��ݑ�5��X��sD}E~7h��01�/�L�Bu@>驥��G��矫 ��G���Ҽ�ݽ����a��=���-,J����Râ��n�J��0�u��b�C� �ݮ�N��Օ/O�2���������C����A���A����8�𡤼
�PRDT���AA�+s��Cwڌ�����[�%��cZAk���}()����&ycc�z:�T[-(�l�)Z������0e�S�?���7�L5��3@*�Ю�}��<D6���Ңv��~i�S^��{t�����e�L~�W�����������Btw6���+��h�oBG{/��(��aw�ecLĀ�l2��4C��,��<y|g�'ZϱI()*��gD�Y,.o�g21���=�?��g�`����>J�)�FP][\��c�aL'$-��;���<>�?&u	׀��f"��;÷��R�c��?��S�J�csG�y?���f����//-h�c��I؎�����-�m��3�E9�*<�5%�����VS}��}�-��'����UFk>G�����T'dR��1*�]��PT������m��ckg[Dh�9��w/���+�,��a"���DY]����)�����=�l�]�h�.A�	�o߭���L�2tN�dpB����� �f2m���%f�W%f�9��9ݓ��M��Y�$�:Z�T��hHŔ�86C��w��q$�h�Ld���HE��lnD{s�.�0>�VFi�X'�pY�q��0WClB��TE�b`�A�5���:$ѐ��J<}9���ϝr��:3&`2g������d�v�2����	��`�{���mM�~B�s����'2��L�T�,��܊��fA|d�'�I�Y$��]�T��!i�RWQ)����	Vu�������J �_x����JjFh̆��}�l��E�!-܉Qo[W[���B̼���=a`E�"��3&W���S/3���f�Vb����=��l�id)��W:�̔�ݢ���W>T�p��f1v��;{݂����<]ZOWKNqys�O(2ؤg�[WA��E�DR�����0z*U��gL'�r������ R� ��qrq���bL�����5�2�����5��am�s+[*��c�`�R�_e�S�ƑM�q��~.��iY]^���>��GQPR������p�;���^j�4�A?*J��O���]<��,8��.;"A:Ĺa5Y�Wgb?'/6|��'�� �`�9`a@Ky�]n�<ʚ�����Y��W�7=k+|_�[5�s푉G`�$Q_S�{wie����[q/>����0�W���x��C���(Ҏ�ɋ7�X�9��Q(�!��\6|��c�~���as���X���:M��uOL�A �PA����.��:&2F�����{,Y�ɄN��mNx�K$9:��7��=���]��OF2]�_K%�٨�� �-�5�+��� �W7�!��݀p�ǻ��Xz��)�y��Զ����b��+�F�Ubh��T;{ۊm��hEe�W��|7|��"<���x19+�T�&0���\���C}=���/�����nGkS=f�g16�H��S�3�%/�2�l&�Z�u���Ŀ TI��S���!��x��K���D7RZI1����Yg��`�ZѰ�T���"XZ��?g4�q���w�D:~#5A,����mAg'�e�6'>z�P�1凌�i�?zxW�3���^�y�"�`l�LB<�s_ogVJ�i�ͮ)����������X��Ӫ�Nx����!�4�x0����k50����O.��|b�IrSz����cw�ȹlko&�fʩ"����g�9�FZN$� ���_
�1[4}��� ��+8:9V�y"z���g�]�D�ӄD(��N�{us߷�����
�,�Z*�PY$r,����k�?<£;#J�㚆k����*�5�j�sF.|�ZXD,�����.�l@ecJ������CN�ee�"L����iwɆ9ǘҜ	6�#l���	5��__YV�
5���h���f��6����Ҋʼ�i&%~Umu5:ۛ��̈́�D�VGg�ӅǏ?�����~N�݂�c���QT����^�L#ER��q�XM�.r���������m��B�OWO��?��x�J�(g��cd¨�xQQT"�i��@���X{��b�q/@!�B_w'z���n����K�x5��DD����1E�h���Ļ�5l� ��K/x�h�A���i��̔$'�|z�{E`��pau�<�VT����������"��ry�B4@.����c;�d�_Qw~y-#�p("�4��h$�n��̔{�dVSY�����WW�ņ|��c��`��U3�%ǂq�o/�hm���9h�A��W)��@�\�g�Rw˼o#/�,B;��11��g�x��>���ׁk�������!���|an}��{�yJp�
"e�'<D8p�wo&�Gf~gw��z���\�RCA?����lm��1�}.�c7h���.ۈ(���kB�kj�e�Nf��]���2���b�~�o�L�� w�����5���D�����]�I��d)��c�`m~{k�ȥb�H�c8�н�Q\�$�����͌H�Z)^==�������:��չ�{�G���ۉ��5�vO�v�sk�0ڼڡ[mF8�����}B0(:;?�w>�Օe�};#s6�>��c<{�\�r����P �a���=V]�� �N��H�S������2����	��b���$�*�e6�Uu���_a���ee� �P�
ק���z���jD6mD�X���OQ�ܭ����
<<zp�������ꊠ�[-HD#�Z�X\^�?Q��ݘ'GE3�����f�
�ኋv���5>��L�f�g��ю��MzTL�55���$,6F����O�F�Y��i����*�
�ـh�e�N\]�*��ns��*,����E�K��;�We)P�e6
IˤS���P^Z�PЏH0���Z�o�ʘ�:<r=c�m��qv��噯�����F*m��U��{���QZ`��M'�dF��dj!�k���Қ��I���_�b4�Ƿ
���'2x�b
�Ta�`��GbJ�jolF'�/1<<���"����?��@����5������_�x���Uc�¢��HP���p��BH���#��CGC&<��ǈ��� m/����ܨ���ى�c6O�F���>�sO%c�$o����8ؘ�۔֐�����)���6�+��焞���р{����O�jc�[��b����}O����32��j��U���{��_ے�.�l⸶ Ɍ�R�|���P�ӣ�����'����߯�]� !�R*(�T!3������
�|�L���'j�y�����-�1�(����nyUP�ƵEoO':Z[0?7+�^��8�p5x�V�
:w�M(,���k��|d�W!��x��Ɍ�Ŧ������¹����=㿡��6��?���: �0�3�y�ʫe~q0,�#;���.ܻ}�`���bѐ�#Z�q���T"���6x��x�f�f0|{Tv��XnW�V���O�t�,��X�In�Z_UAoh�S'\R^�t&��m����&���s�n�"g���;��؜ڧ�� $�BCk�����M��}�yH+�k4��L^�������_wd���<����
�>Z`:���I<�]������m��:�I����#�(����I��e2��iǝ�~���N�ɇ�n0*u���/_>GGS��%��l�����T�<�]��>�7W�x;�奅�Y-:�.�G������PV^���g����$!w���oK�c�������.�L*O�K�qvr*?�Al���"S�ϊ����Ԡ777���H�26t����R�?��M��l�efLy�o�>?!ȝ��g��cO����/D�� �!�h�F�XyUe��b�a���#Ol�D����ނ��:e�^���Q &{�j�l�hP��镊_�[�0�B��uX^YÛ�y��~�_��ȁ{G��<L�3e���6#��
%[��HJ�2�.,"g���r��Gڝ����D���Φ�@$3}�䉌e������>�@o/&^Ob���No1����-r"`�y�yc6,�0�k�;�h�RA�͞3��yrQtu��od7�9��v����aܡ[���]�A��!�Fc��L���D��5!f�j]#�F���8���u�h�3:��]N�{�[�dM>��w�6������Vw��Q\D`H�k.�#�;
`��qxt�K�w�Jzn#�:�1�/��]�i�J���҄��S�ל^�K�PS׈��=%3r��N�p�C��K�/�W�ѕ�͂����K<��($�H�����u
o:>����<F�{	�U<_���1��l�$*��r6��A�0ک��Y�������!�d�ÂJB0��WW"s�!���&,B�00`(+} �q8,4���D*�E�\N���k���3N��t�1��h�æ��2 �Y��d3\��ק�}wuJ:�\"�,��MnT5�B�Q�5����&ǥ���}�:/���n�j�����ß��Wo)u�RAg���U���c�����Wԣse���Itwr�ⲉ��N��y�=|�����U���T�6�u� f���A$���SÕ�%�(������'����
�N�l*e�M����'�*��B R�QC����ݝ}�V8�V��bcs�U%&�x>9�$Yt�p"�����n������6���''n��0�ɚhkz���DR���DMuj+ԡ�5Us��J�-�TJ�������[=�pZ��s��	�����j�P	1��[VAO�?���w�yz��T�� H�`&�sw����43����k�=���$�?��`����gd˲d�Y�	����9'� I�*Tλ���b�����4�$
U��}�p����7�q���R)c������V?��&�'��Ԅ����מ��;�-ڙP� M�"ꌵ��!�^>��tqCA��ӗ�_j'v�u�n���\���Y&7�Μ*������}�H��3h��PH�ӫS�����Wf���\�bm�F��?�hװ�t`i$\�'�3/��d�K�fA���'?�@���Jr�n^�j�v찭[6��0���dB�{2Wb��γ�O���=���Ѡ?vTz#���ҳ�����п����+״�c������662�DR�m_�`�k�j`o:z��{zev��"P>�
W5���m[���Cv��!;���8��#���]c�����yO>�n!o�).U��mv�Y��[ݠ��+�y�YҎ�3������S��L�P�o2~܇�����~�@�v��={��D�d�;=�O>8eS/�.3U��{���H5����v��Kb5S<}�:����Y:�n�Dס��6��GG{�����;}g�����0B�Eb*,Y�@��Z��|����,�ûw�đ�KAƓ�v
u7_�2(:v�,��N	}i��U�o5C�����z��WJ�A�$�Ǌ�u�h����4����C���ǂ��E��y��P�?<��N!W����Ɯ��el5ۺ�[jp�/_�r�l�pD��nCv��m��,-��ǟ}��IT����U���ŖG���)X,�C��]�M��L�@�x�@��DA�9����+*ș��C�L3	�{�|����ﷅ�{�j��.�����7l��c{��Hq�ku��Z6��S�X������[!~��+Y����w����]X�W��o�u��8����wX$��{F$x��r����[2_�Z�ge�0-jk�����%V/��ymǞ�����H�,��f-�9~BB&S�o�V	ZGQ !���mV��9V�z�u$ԗ����@FN��HBD�"���E��b��w���n��ȘM�\��XȚϲv���J��=t����!�	gn��X���3�����Aw<���<Z��:��ʍ�r�۽u��^����Yu����t��h�`�>���%&_<�SǏ[6�V�=�����k��>�1�� 5(�Vk��T%1ˎSq�����B9�j���@ݒ��^�H�0م���'�wu$�7/4��F�`&���	U%Z�b���E������̪��xQ�F;[�Z�}~�������ܡ�������?������~��T�$�����'�"�n<l�,��)|�W���ƂD��=/������u��mld����:++K�Og��?k_7�=�Wof�jq�j����!S�H����5��ܽþ<���{�V^�G���w�1�z�,��(@�� ��^'�F�A�����&v2�p$(�����Z�Y�--/*�3˦���:>T蚨 ��N�x��*������_�e���M=�m�o���񞺶���k�[O��3� �a���=Q����&��vH����&����svd����:҈�o�O�˙��Q��]��\�N���675!�m�P�WW�R��+�ڕ�'�;t�=�����5n�FrE�U4��epPb���b�;����@�Q��*ǶmWe��7B&�u���?W����`�N{��h�d�W׭��[6�?yj������u{����73��C�v��Ϭ�w�ֲe��%�/�O����Y,����c�}����4,���o���c�wt��H0�^�mX��<�O����}~�#%t����.۾�b���Z�q;wndD���~h�.~#�='��!HH��KYV��E'(���8,I�K׮����:�Q���ոg`pP������Y��o�<���H(h=���a`ӝ=z6�y$H�U�[x��߽bar�Z'9���A�$t�A�V��`�
Ļ��ߦ�^��#�m�Рy$��S1�h��O��^�*U�ٹK7,�sJ~�@�R�+�o�6Iz~��/�9iI$l��ذ�����e�
s�B�b����>o�T
�*	{����6:�٦�L��浹�w6�jF�Ό�p�c�
��Ω��#�[Ż������ߛ{����_�Hz�qe�ޢ-�~l�n��jnE
��Z�"m�6.��1Kc+M��� ����:��������1�������Z��=6d�t�"-����aw����\�ʞ�Eba���"n���W�����;|���w�����~r���E	�$�0H�s�Ob	Lmfۉ֨�f[�9����m��k)doQ��!纷�Gn{�Ss��٣]k����+I��Һ-,0�+�C�
v��W���MqF@vP����=����;	j}e���c�n���wD:���*������+7�����ǶZ��h���_�˷��Ԋ-�S&��o�ɓ��έ�zjR��}z����O��;0(��;����5�9D*(|�Қ/@�`V� �Yg��D9ףVv.||������a�����5��ĺi�VS��8�G
����Vf�kv��m[�f�
���⾚u��}~l��~z��oN����֟��/��J���l�.U��N���;g?��@�ӻ����lcͪ�}a+1.����"
Q����U1^�;�e�I��\p���B��kwڛ�y�+3K�Aeg���}��n����
"�n��g��e[^^�pږn    IDAT����\� &:��*}�TZ�*V<�+�O����j�3yaᝠv>#p����ڔ�Ixt�@�n
���*�k�9{��%�}�: s�o�o��_Z=�,��^�4_k����-��o�"��q�����'��^�0u[b�>���:<hu_ծ~s�N>h݉v�Ƒ���았�OP,+t�?��c{��M>{$	ݶ�xC{<nkkI���3S�yd?���K�}�ּX�b�I�Wc���0
��B�}��&ɜ`�}J��n���XĶm���zr��-8���!���?'�`�Xʧ,dE���'���y"��,ڹ��O��h��<r�bF�#az�B��C�)[<��xĆ�6��yx��m�l��b�S+���G�bz�|�v�m��w��{gmvj�&��Pw�+�mdtH�N�Kk637�����;t`�]�􍭬�$!Y�F��a�c�]Y��۟"�����6�6�f��̔���1'� <@ÿ��j�k?95e�m-Z�۹cLɒ����c6��,l�3��F<��<g3�Omq���rKٻ�k$�M���*|��W��2X��p�_z��;w��;-D�W��Ru#�UB��r���re�x�$`=���rz}���a��v�����?|Xֹ$����O��6�`�0Z:��Ŧ�e��b��g��θvI�'�h0j7��uk��,A�Z�J�$�6H���x��_H{�5M��Ǐ����Xk��9v��l��C{|�y�)I��D;�؞#X��v�(ŷ��dۊ�?r���E�\�ث׳*��ݦ��t� ��+�^Z	ϊ�F![]y'?����Ą��(Rqr$���|w��V�`��P�HҘ�V���߇�k��ﷷ�sJJ4	 ��mdۘ��(�I2����S��翶8+����2ļ�7�k�|��1i�?z��֒i�T��G+�%Z��׾���;Jq�zX�{��NB�aٶΈ�o����?fO�cϞة����!�W�]�"E�C��$r
�ljn�n=~a5�O�zp(n��vwڍ�����Il��j̰7]]Y�����a{=7gV��I	��D��g2"<b���f�d6;?oAܡ���QO��3-/���
��;\N��$BEl��b�>�B�l=]]�D$*6?��Ba�m�r�+�ݘV\&���<�)�����?�������3����p�/����T+���{<跷`��X!��f��-��Ν{mǶ]���嗅�q�t@�"���p1r9�$���d�pc#c'O���R.�"�ƕ[,�O�/�*��N���^�ЁD���b�d=�����VmWg�}��Y�p劼ms5�==bs�uuK��^�n�D}�/e��z�n.��D9 �|��O�Ee
��CFBg���T�XU�${�r/���]����[ZSB�I+��S��C��J� ���AR��G0qMJ[K�����P$d�K��ُ�'�2YA�����U��Kp ~��Y{3��ݽ)q��*y��Nמ��:�CY`�`P�Rx�=����-�I������)[Y[�=�C
��
��#�� �F	,[upؿ���d�|I���zR�=mO)mw�}m/�_��7(A��x׈�9���;��P�oኌ0������Ke\���-T��#b����^��=;ml��=%���G/���9�Y�����v��1�ս�Lѩ�7�˖��mv��پ��鬽]^����X��ծ߼��xG��K&x.
r�-=2���&��'�@�^����?�Y{��YK[�:���ӂ�򙴂}'t��޽u�	�*<�������}�ĞܻjQoN�m�<ҹ��Џ���V�b8�]oV�+��aGU܏0֑=���S��΄ݺu��RI;}��I�+�]���R���w�%ٹst�z;�v��E�k:R����>{���$��������v��M+U}�Ε5G ����槬�1��n������wf�/�o,&ȝ���)�*�g�;v�RB'qFe:��T7W(�mzvA�;��J�^?�c/\�zi]]n��׹�y��m�eI�'�{g��a����a�g���v���3���r�kl�:���ثX�o�M�����lnC�<��`�l�O�Z�����]�Ĉ�d:���w˶��l�=���+��X�Yr0,	�
I)��α�Z����Q������kieu�iSHv��Sfgg԰�l����5>z�\�JUki����c�]��M=�i���f�t��{��(�3C�P2�H�^�LrͶ�w۾��,������;-:+̵��pY瞄������y��*g�@((2/�&��̼�A��f�Q��Hf��]���f-�.����z��i �7������[c�1������1���%yu�R��l��T*E�zdA�߯��;��P_.Ś�@�Ċ�OY���h=4��nڒh�l�-���=���]��	��~q����j?N�JԹr+k6��Q���+�w챁�!���)�
4��i�z]ںRȪV�cW,�Q�E�1it������n�o޳��_(�KԄrO���+���KU�;zBU��Ĥ<r���t����+u��y��*�����ޟ?h?b�L�޼��lљaط��b���� �GŅ���I��{n����jRUWG���r��0`a����D��^=��Ǘ�
+��;��]2m;�ۑ�O	}=���9Z�0K�1qp�li��p9�N(W%�����Û�T�p�П���*II3��V�N)����O;���Ҳ<�}5�VX6o��MCv��-�CFbm�L�������c��S*��[7��ˊ-�38h_]8/�H��t���Q@ù���^����S�Q��C]�Z�+���C���j�.���ա��y��[{���cY(��re��APc�)�`��Wp�#�[U��M=>O�����u��4�x�f�5�yH�[����}�����G?��=|t�&_<����������W���?������y�����8Ε�����3�Y_��������7n_��*x~�����1����m"~�_�܁��ٽ��ݽyC���-��(��[^c��g�@UZ�o����(�e�^B�w�'J�t�� ��5�ǀ�ynA��B�⁠�=f����7��A�Sǭ^�P!��-	�L窖+2�X�[���6�=��._:�:���=!ao_��|�L���n����]�v͢-�{-��:/�̆�c~��o�|1p��\�u;����꘻��U0@�D$��]&�f�g9��1�H����n9i�mQ}�On؋�ߨCW!YXK���QH��ڐ�CȦ���G�S4�o���^شɺ�z%����aw�H�mp�{>��.�zf�
r�}<ⷣ��J������y$�k|��
��.!he��	Gbv���pCB���
ҹ�Ժ��A<�&w��c��?S"ޱs�����[������B��~	A5@B) �e�4E&���w��������A<�u� w:�8�Y@ٞ!�������[c��=���cD�E��{��mG�1�
dnrf����S#�~)|J���.�˗O���d-�� ��>8�����'r��>&-�Id����>�/eJ��������7��h��OB'G|i�C(39����9����P���F�1���~�����[N'�sS�-&Wm��ak�E-��,V���4�\�fE��nB�o?���?���G/�ք��~�������{^��oۮNpN���7�ض�c�b��y;��B��yA˳o��Y��%�Q�R6/����NAe@�����MC����;v��3E�Z[aV	Y��f_�VG	C{qqI�7CCC��X���;z����+�,�\�I���<;/��nfV�`�UM�>x,+�O?�D75*-	������{���N�:%���I���!uf�\�$�L�d�3����V�.[�ϊM��2yk��b����T�R�5�qAcW�S$�dv"�X����L���ul��V���餽���"��x�өs��7agN��׿�Ut�?9+��H���Ç����߳��5����[z��&�0A�W�ƽ`T�E�ɳ�{��Y�C""���٠ b�����`!#,�rⅠO��U^^KK�T������m��c)�A`��m����>�Hǀe
u�Hx>DfpE+)ز��Q�PI��/$+qQk��� �{�g_�����.4�����E	�N|�}�v������ػ��_�d�ָ�ݻwŭ��0�y�-b@��}�V��@O�*���S*I�s�o��tI�?
�V�g��D������|d���eS)��g��˗�b`Gc�v�+�^���.���#{��k��-���wؾc?���q[$�|�}/W��E���N7J^$fB:�a�&W-�g)�mtt�>��+�R�N�����������0�Tx�����=������۳o�`{�ko��x�\�����x����uX��S�k�=��G��k��6]��E¬{����[B��|�:pP�o�޽*� |�lf>J��1��8#X.w�I�I�r=oOn������$�R6Z{Fml�	�۲��A+I�@�O"�e\��w��{�������3��?���OQY|�z�~��em�@�Bx	&���;�=��W��^�X�ڑ�8�?�؇��=��b�bWoܑ�H�|
��{�h�K��ƀׂ�bjJ�>q���W�~�ײ��m��z��t��֌��	�C`"q��_S�T���`W/������tR	R	��Dﰄp�!�a�B�юQP�l�tF(ީc�lh�_1��y��%k�F���1�ϣј��gW�?�b�.R��)k M��drնoiHv��9��ƍ���<y:�.%��ϧ>N�vlӸ����a5C���oX����x d��}B �Z�[�ƺ�B���ݽ�����Ƕ�ڰ(hA֭V�U���bm:i{v���ڒ]�z�|���I�@H���z������'����	�Ͽ�=��|�'�@�A���&������J�wd�@6?�l]����rCC����{�8���k�#]U>�� ��k�u3]�zM��$
�؇���y�����D�s�����҅�ldt�m�aw�=�Q=֔�h�*/*u
�b6m��e�2�'b]|~~Y���Q������qP�s���K���|�_��mݲ����a��J�����ƽ����WK�^Y���Ƕ��U`2#%�ۻL��#v��ߵ`�˒ɒ�|n7���:F(�
"*�D'Ұr��!	�k�H��7�)�6�9�V0�	JX�n�V���ON[!���/���>�D9_�_��K1�Y�{p���Ƭ���Ç Al������/.�:�aٌ����M:��,��ג� �g��p��Ʉ�I�~`�f��Dm!� ��]9���z��@Udò,ֻ��?k�ĀD��V��_��T��#�5������D�o��T�j��V���w�����֘���[�l�62*H5��;i���w�L���?��z�x�m���)��*E7F>OUs�<ҭ敻 D< ®�v�=aM�R�(iS�ۺ�я\e��u����cIu2�o��d[Gv����] u���g�l���S"3*����g6�m���"b�|e���%�k�)����6-AĂx�I
�r��fKtu
5�p񊽘��(!"��;|p\F<w�ޒ�6�����:pp��ܾ/і#�NJ����$�%�)D�JŬu����@��^8�t�[��������ol��]����$�p4jV��nyI[�h\�8Ik�(!�f6r�bj������mٍE���k���Y��`�BV���?���{G-��X8��+��\��s.[�\V�]���V@��6�)h���=��~�β|�z]�.<����vٝ�7�RK��p��}��|�A�R?~����鹷�ZX�lh�D*u��uĢr�{��P�\� )�*��.�[<�0��Z�a�d��󉩆���Rk����S|�'�)$Z_(f�|M�^��rnMkkSOnY�S��;g)_���A;x�c��٬�LC@D~*����YG�3��3�� �޹yK���n*� �-��onܒ,�K["!��4��}��0.�;��#�^f����FL=6��o�)��h��Q����)0Z� �����1�|�Z�W��u�۵֗�钿:v���	��miv޺�:��>��R�?v\��ք�Z�]m6<��b�]�q�n�O��	�Y\߬j�Gg�������_\������W�W.��2o�c[�{�n3=����ߚU��k�^�����e�F:miqU��
=0�Y� �zCV��6��kqh�gp��gT���]Z[��90P�ZQ����H`�
R_Y^t�,V������;v�w�v��ck��t1���!�Wn�[��E
d��%uJt>�m]63���ݑ�kn�2��bPI�C�x��I�n�%����-���mǮ=�yl�=��K|YkT�Z�f_<���W�����L;sE�ٺ�N~�9e�����JƵ����9FVw�\t�#V�H|h-g�k���Z�7�)��&X�%�������3��d�:G���97;/�ۃ��������&�s���)���~��0�jOX������s��~�0�+�H8װ��[vm}�<�c?���I;��z��_N^���-���w3v�ү-�4k~/���#�3d>��ź��@�ÈBB�.i�̿�����u�H�ͤ�_7I٢��%�1�����c�a�ݻ�[<�7�����[�_n����X4�f_^8�y9�|����S����shS���1���!]	B_�!듏?����k���}2!�|1��Q'F�K!���o.��ꚍl�m��=���k[]]6?+~����m��M��G���D�?�=�r�U��=>+ϫ[w�ѦR��~�9����Z.��
�Š�ok��l}u�Z[�3s���ƶٱ���g?���!g�~hk+n��"���۶sǸv�����ȅ��q�CF����;��y�ضQ1��EI&�`����a4F���1��5�Ξnmk>|D���'Omx`P�axTw$z���+{6�Vz ���-O?����[��t&3����m���[k�6��VdBD���sͪ:{��+n������d-���x��6=����y��f�xEtuu*����?�{����/�������?�϶o�ۼy�֮���mc;����Q(hy�dH嫕���Mʈ�L^$��[XZ��o�g?�L���ד��4d�N�򑰸��!�����%؃� DLt�Y��܈x�_��׿������WҬ+�|�o�F�m��3��Զ
�I��ͼ �SPI��b���:��m��_�+�\$���E�b+������;w���B��&�sF��0C'7 D�����Y���/�;P;*v�6��u�I�ؖ�~	B�]NZ�Z��7��nuUh��w����6�S�6��N�0��0N���i�5�/_.歕x��,����n%����9;r��]�}G3�\ݑ�bL��=��O�����~c�NB�W���?/Gc���́��#)��c��m���A[^I��"���|�u+xV	�9'I���"��tsJ�* R������JTw>�E�א��GGF�{g�j݀)����������0׈�Y��TΘG���S���Y	�����:���唼�a-3{�]�o�]W��ss"���c`P�sK$jW.�Κ`�vuÞ��q� ������7����s�+e���h5W���=v�ӟZ��d�`>4��s%��х (�;Og�e���Z�6:�.���X=+C�z�'�  D~�҉�X���u߷[�k�k"Q�<pH=��O�<�Ì�b���Zb �]�%&�r`_J:�n�tZ]J2�;��LeܑhSgI`���D7��,�R)g;wm����'���[�X��
p)$���b�o���'w��A��8�E;6ۑ3?��ޭ��ʺD���|5;r���RQ����,�3J���t�3����nz����Q2�"���lk+�6�uئ�mfa��V��Ȅ�p�
�E�������;����I+4L}���YX�|y���Q�ZC @�}eqE�N�O    IDATOO��Ŵ.���=;��b�{z�oeiݦ�ް��;���rYV}����Ϭ�n[�W���kS�QC����exj�s@��o��f�C�O�.G.3A�|��\�Y`�	��#���.ك{���|��q%a�~�c*&�OL��mh�Ke�Vȣjw���.F�-��?
�&��g2i���Z���,:'H�3��3���ʥo,���Pӳ�O$����?���u{6� m����{���������o��~�k���C�$���!	rӼ8��g�TB��#Oq�xX7$��x*�g�_��~s}x�s���"����3u�g�|��j���B�K~p�V�sv����5E`H@ӕ\���%B��L�2����lr�T��j�Yo��ݕ���]^�#�r<�\���)!-+�IKgKv��I;� f6QjŔ=�yަ_ܱVE$F�7h%Yϖ=�}���v���J�G�ӰZ�����Bs�⚑F]�
x2]m�T�Ȥ�S~�/��^�d��]����1;v숄d0Rڷ#��]FXft��k׮KY�&�ޣG�5�549M��A?�`�Fm��A�j�|����-�g�֝�����Z�㷇WoZ[$��52��n>�o�K"�&b1�j��d�Q�@��WJ����r��
��M����{��uu�Y�W�t�*�\�Z�T�z{���c{���&���؟~��Y��?A�	Y�z:o�JE�/0���#��[[{��}�jܒ�i���
�ЩN��c��D�j�N����O�A��6HW,�#̋N2��ʒy�u�hkw��D�F�l}�뷚$��J�٧[�/�bc-� ~>�?���9���V���1,��T�(Xn$Sg`d�Vf�M�fV���l׎���~���V�md��j4�aʶ%���5l��-L>��wΙ����X�J�n����'?����={�t��	��Y���D��9��TJ��P'�Q�!���V�W�Nn�6|~�JUKgVe����C�F�B`@�ؙ�D�:��[���?�0L�iP�a3SS"��&���u.+a��#[}�s����H� 3��	��������=$Q�gS�v�#�Q2Bʾ��olcqڼ��!�Y81`'���Z{��~�#�f���\g���5�%�
<M7@�@=�'D��-�>g���O6��gg$����:]���0����jv���\j�.)�_��pv�{:D&�"�
G-[b}�[��C}R#����.1�X�H��E���N��lx� �g�Zq^p	r�E�|v��X���o�t�⭽J�=Cc���db��Vt��D
�KrE	iyS�_�nt��Z(�H�FRxJ�BB��*i*�uH`[G�u�={js���KGF�ivK�r����oW���K_ni��:��~�r�)i6�a��=y��6�l�ޮn�ta�c���]X�7������G����f��>o��v��I��𱌍�m�nx��=��s����/d�|{�4�i��d6�D���ֵ�VP>��4�Q� K\:m\�(J�� >�� BҸc�t�"��8yL��믿�j׮"��V���ж��/�8g���P�F�� E૊�T�f�|Q�O�����KSx�Y5e�<`Q �3f�������ʜ�w�?�+�ҿw�c�������ˌ�B��3oe�ݺ`�/�Y{��f辠�<a��m�{�Y�s��,�#�5���{�Sqe&͉��<(4:6>��b��sJ����uu�ؒ����0;#�͝������W�R�4`�.]�Z�W�����u�w��b�S��ְطۊ�m�d�U+�=��լ6���-�6�e���ڮxGs���%s	Rm�j�7�ؓ�����F���R2i/'�-����Oa_�&_>�dj�*����:��XX��C��g����	�O�������?��c:ra���!$�QJٲ%ڻ�[��b��X�*���-P#��p�$ғV�� �N�Tw��V+P#�c���
�y��٥U�Y_��Y<�&����]P�:�����s`�#�G�ɗ�qIA^R�`��"�����S'_5��x���r��d�\�b'�����U� ��\Ƽq�P�W�Tm��6�,��e�V��L6�d�c�#{�ȇ?��'�LP�0��0K�C$������U�y�ur�+�����zdA��^���2�J��5H�(q/I<0T�@�R{�E]H[%\�|n���Q�������Z[(Ңy�濎���mu����$w9��o���Y�԰�D��.�$$��d�ʆݽ~ޖg^��k����X�f;y��r[[\ˈAM�$��F�vݺ�cl���>��`G��H�߈����Qg.Z�|ra��Y'��̰�q�%�Zn�,��z*� ��$ߪ�ѕ�+b�?`2&!@Q �[�?3����E�Dk���ZZJPx��C7��6.to��S��V�[^�g�Rް7/nٛ�w�B�!�Q���&;p쬘��H�[m�)���q�������%��R�� ��#�a�Ҹ�2�!a��Jz�$�94�{_���<�U�\_���i���Z��]�՚*`r�ሊ ��4%Wj��ttuة'�s''&dR#e�|^g��8�}�ydr���sK����O>�d1e7�=����qR��_<��g��[H�@	�?ڽ�v��b]���u"+Kx�{�>�-��#�I���A��Ļ�Y""�H�EEg�Y���2R�ه�	'e|�n!tw����`��xa�بݸ~����6�o��E';Z�J-�Y:���o@fK�hT]���9{����1j�C}�Gk�ć��y���4��m���i���k:w�:�m۱ۮ\�-�VK�I�w��"�uE<��K){�ֽe�Fv�x�Ti �1B������ t�)�q� �ɵ�\�F�n_)�^�,hLW-���=JK,g���჻����-vĶ�w�����'657c���=����ֽ�W�P�V�-��zgw�-�lX��C������Gl�첁�.�9���o,�������N��7n��R�v����m���v��s[]IiO�<��e��1�T��۵U�ƢV�b����f�]�����G��ā�L����Ww�٥��b�����X+����v%t`$����e3��"���IIB!f����qӊ9���JE�R���G���*���	�$~^�x���X�����ϮA�p:�і�<~��Y_�眊?���Ҫ���D2�k����dk�D�������d��!�֨9Xt�T��v�Px�mҥ�Չ`I)�dS�o���C��W��[o����w���߷b��=�g�zu�� �^4X��p$$r!
d ��;~ 	��� ���|/U>�,�Sz��R����� �|V�$xَ/��%#V�WK�Gت2g���d%qM"�����F(R���4bH���q�.H���H0cymE;��ת��]���VL/����_֚��#v�Zk�� �|)��o�`A��o�['l~�/Ȇ.ӑrFkV'q�����D~�*0�Z�d�ؠ֊*���� �@J����r��.$�)�j���T�A��aղy��v]ٓ�3�������=��!ӿAk@R�~W�U�Y�J�^=�aӯY�^��D6U���Ͷ��YkI��h$t�An
���)�q=(����!	_�a�C���gձt�ｂ���V���)p8�2$(;���9��:�O
w�	Q��U��so�*A�����p2�⿫�ӖW����]Ϲn�{0���g(l=�ݶ����
�KF|s��Vc��d�;���[6q�%�H�%��v��#�-��o����,��;7�u�������H�*.��5T��E�ی�b���y��	�&*���޽{tAI�f�5nܸns�o-�y2"-
�<s:ی�2iI4;rD���S��B+��Ɨ�ѩ���m��sw�ص�r?L�����%9rvzF�ꃏ���ݾ�P�v4e'e����f�ݲΘ,Bx$�gx�F���. w�Cs)��rș�2+MK�B����ae{噐5��"�x���y����J���q��^�|A�0$W<G��p�� q�[I���>_���#���ׅuIv�9���ۻeNC��D��Tq<�XĖ�I��c���}dľ��լ�U�W.ڛ������r�ޠ	������]v������Ö����K߈垫U�Pżu��3����5����k�~����ա{�f��l��e�s�淕BŶlUy�fNу���͛)v%[���`��\W锜�?)�����7�U2���B�<����%*Vw��V���7�dt�<dT������� >�ZK	��K�Z�Z������Z[���f>�CW7�iV��y�TxT)GQ�#�cLz,_r���#ު2�v�_��Y�(� A�u`d�8��m�k�`g�Ae5�K�/A
�n'1���u=�����]��
���ê�3O�W�&b�|Z{̬G!`@�&�������W\��:�9a
gr9�"'$��16�N	�`��/JVH5�G���Ƞ#eF�������L�sE%,PTڬ^c��ol��ͳ���J��|d�X�.�9�sqG�".���I$�f�����k��b����dW�T�>�0���;������@ixG7;Z�jR�Y*��񸂌�-����W�p4$�P�@@��9I��T���g���p^Xs���+Ho��ع�Jڞ?�f��^��Z��*YO�f�{����{-_!<6k�8��k~�Sp�ŃQ�itU��:��a�P䋳�s��v��xV�{F��0��utu˾MP�M:�����ۛ��g���y����BN�#H��^EZc���.�d���ԩAH�2@rb�$�*���l��={p��Z��t���Z�����G�~!��f-�q�ȱ��)P*�$�g�/�?�Y|�9�}�=Vȁbl�� +XO]F#�>B:�[]%'��FH�D��<�I>wg"��Ami��d�"1�{@�r������*��.DӇrhI�g$z��A#����Q�ڰ�7�r�m�P��t���uo�g�����\ en����\>ڂr�1b�r��˚
A6}
p� I�qE(O�7���S�E6}�zJ���<`w|��W�6_8f%��~Lc@9+b�3}�m�o�q�%�	@b�]��z�Zm������!�8T�b֦ly}Eg�����)W-�����͕�v��	�����+@b��c[���/�̙��X�x� �|�ۄ�����٣{����-��Kww��_��_Tc�3�jj>��>��ݾv�������w�h��.:������܉]��l�1�!�8��O�h�و�Mx�D�̜u!:fV/�a���dy�I�]�n��a�N��b�u%��x�E�
� (3��!h���C���r]']9A��`F$p �3tJi��
$����g&��8i_UePR�@?O`��B6��=�}��՜#Xy�T��?������TF�"<��8H0t��yŢ�@�E��� YP��T���� G)(��$)�?;�l�u���
=~��62N��ș�qz��F����U⇹ˋ�P������\@#I�e�4�Ӟ/�m��Ԭ�<�� ��������%��xlӓOE�*�X{װ��:de_T^���6'��}Tm@��hUd5:r����[��C��HƑB�3y!y�gt��h���pPA�����2'e����Y;�t��)9G�tR�˖�( ꇈ�<͕�V/u�p���y��,1#a#���<�ݼ%{���--LJu/��[r-o�݃���	���-����(�5��;�N�I*��s��[��p�K�9�"W��(�,Y��QT�z��Q�`��(�^wm6�5֪��s�+5Gg�s��/�y8�޼'%�㚨���g��

I�=7���gr���o(�꾀m�a�X�R�^=�c���6��[�k�Ə~h�N���QD:!�/�<Q��J#ߜ�K����"��V�� �q�#���1��o	��u��M��dr]gÍ�ܸ���^vr#��(��rQ$I~Q��E��� zJ���<ʹ��)�U`���^�|��A� yx4$zf��
G�5���WOo���(oX?�`�r�un�k;����4́egAЍ�3W�XI��%t]����jm�T�Pp������&�Sn�V� �v:!niۭ��K�	������L�-�w��9V��<��F
��h��{�����ݽ/���{�d-�-�Wl��]�Vm��K�{�������A�3h��zZ"�=}�X����c��u����+���n����Z��{�������'��IB��k������C{������x�~����v���p���.�?����fJ�S/�;�b�uy(�1	� �y��m�i�q�����2����̤��Á  Qa�48`��[��"�ù�:�%صUcd_%T���
��y* p��hǘ9 �^���L#�*J*TX��Y�p�@�k,��E�
b���@�ɋ�΢V��}�j�C�3��~�j1g��K�t�T�T(X�R�#�'�xG�t�Y���HQ��:����<�BE���kE_�x��T.W7�g��A�n�IГ�9I�% �mSO���~��Xު�g����"I��}�og`��!�+v$�fB�1Ԗ���0���"�QP1;�j�V�lqvJ�4�3�a+[���[���2��E %H*���`���K(R'��q��V��߹Y�KD��Xm#��E����'�4���Y��/R9(�E���cp�8+�l�.���f�o����q�A����p��<��e����V8��ձ`�n�O���C�mm�˔��ۖ�����k�״�KQ@�(f�

D��y!1�2t��3�5V��%\A���k�&��g�Y��:��W�e�Aϼ_�����L��z��4BP��a��?!�t'(�u��R�g��J�K� ΦS�o�n*g�iأL�Nt8ޢ�0��d=mQ[�����[K�c��U�����c{%7����4+��J�t��"i��>��-�BԔ��;&4>*��4�W��6W`�Y��4ߗ�nHQ�d���g�jL��'$^P!^��EE�\��и������w6���
#V��#��;Uܘ��� �#��ꀘ��ޭ+����Ik����Z����v�w���vh�"0a�焆�c�=�(�t��n@����ƞ^�3�)ৡ*
A��#v�Fȹ^±�Yvk��ɜ�A`��j��h@(,�;�:��%�#�Zu1O���O;��W�8d�Y���|��u�^������D�W���!5�G�צ���}y�+��ZY��B�B���m�zqb߶?�O��oL�?;k��z�ߤj��^_H�<j����ɷ^�Y$����w�R�A9�+ѡ�Ԇ����禭R��^�y7�	��P������)�-�{�2�p���ڙ����+~@����t^5�q{�<�h^���^��А�q�aEA�#�Pw�����	�u-���%T^�o7����X���F�y�Hb�RY���Hw�k�F$Ѝ��`w$5?��ϣ@����1#&9I��q�P�c�����A���F�XP@�{�k��tSHG������L<z?���\j���|\�g��]{^���	X�&����g1� }��T�J���ԪD;���Hf����-ot�-P �1BK��\bo&G��]�rp$��%`1Éx��W���5�ytיĥ3��oZ�t$<^G��yc�պ���f�Cwݾ-2\g��>�7�F�{�ܴ���Z?.u������j��S�l}m�j��3]a���K��o`�Z�;l�n����oS_�3^Z�g!�>I�8o��\���Z���I��F!���&�еFB&p��I�|5�Nps�L�ٹ�\�.�Y��h�u]=���X�"��v����}�qY{V�[p��T3��)��ȋ���Ogk�f&�H����O(���Ͷu�n���D._���7`�H�6�i[O%�D)&@�=6-Β���.h�����{\W�&bp��M^�3�~:�ɚ�fǎ��~2刂*�"�4�׷�^�����pK�m0���L�j    IDAT�ȹBl��/���[���T� �Z�(>Ƣ^�ԭ8ﳂ�y��&ݴ�DL{V*�N�ݺ����@�]BL����"�LX��b�F�L�&W���ؑ/�>��t#ɴ�,�H��\q�U�ʕ�$�A��G$}��;E@6���c]<�OH[3vw(���q#B��Ӻ�:��@��
c�X� י�HȨ3ni��{2��_u#�PH6�Ľ��eiK�3�B�Vj�	������m��zyj��?�'����� ������.^���\�7^�y>���H�u��ݎg.����QLZ0���LLb��9����&�{dG��Tr�2�5%�J�*)O��b�6:�~��|A	�R�3�/��O��.�x7(��`j�H���uh��C�yU�ό��`����Ы��w3%w��!�Cř��,�x�"��5,c5�s�!����A���/�l2�3���u��A��^���`�6G�� q}���o��~>$��n'ש0d)�Hf��� #@ܿC�	�.��5n@V�"�����~?6����ܟ7�������8�GA� ��<h�"�k��_���-t�/�ZInX�=!ȏ@��
���u��t�}�4�l4�η�Ģ�i��Pr��n�cC�zJ�Ƒ��Ї&D�g�뫸@�H�0��uc�ʹ&�4�mw�V5��D7�;�0�VwIn���R�d�P�3�	�-�p������I�rD��	jU
���H��D�Eb,�\��ܔ@��Q(��v�`R��\S�"΍}�_�9g����`~7 }��?��3!mè�n�@�{]w	/�zM�k�&��i�m�6;��*��?c5 ^SH֧�n��QB'ȋ��;_(`ɕE+�׭V*
���[w?��V�kD���ѩN4����Rǈ�u�XĹ��@<!.Ppp�xv�s�	���L����،��+)#��3"ɿO%3:G��N��q�!��ăl�pR�;�V��+���F5'�5Vג���j〢��X�x[v���Z�����|��~3�nx���f&����Sԋ��,m�l�o��>غ�꾀$VY%���0��ڠ�����3onMP�qO�ŗ�*%�=�MQr+q��GCLw"Ly[��h<��2k��5V��$9���K�#�]G^"B��d4�Y�=�q1��8��9�ܯL6��K�AR$Q|Pp�3�b�ys�&���]���׭��Ǌ�G�E�W��
�K6��1qr���?}x�ߘ�������+�v�Z;�l�K���Xh��1C�д�F�ă���భ��d�x���ү}�z�6֗��´�-/X���Z�`�|^�_%f>���\P����\v�0j��}>�;v5�z��D�$@Dȡ�Y��{�g%~����:QK�K@bMВ��z}�V5����tz5�2CJz�������vX2�M��n\�h5O�Ba��ba) ��b�YP![T�!DA	��	k�ஓ"3�(
t������ۗm&�M���U�^K��1��1��zb7`���F������]�a
q�qm�]�[W���� F��XAQA����5�.P::�;�� K���(��$a����&��4�p������`#E�C�67:`�) i�][V�R��v�Yɼ�աm����	�4g�U������g�}�Yp�5�8����J��g��W��-��������TwO��<+�2��N�V�G�r[yur�ו�B�e�Ba9�3��\]����v+nߞ�oё�X��>Ss��|^����l�k���{4v�5����O���"v��F���zX�Q�<���&
�b�G��P��(�_6�(�%DVd��[��`�����	� D�[
K;q5�ݍ'$���;�I�˿3�it��q��9l� ����A�����p��E����������Z�+��l�>di���b�|*U����?�ow4b2Ex(&�z��p�p�Qpd�f��s��e��s�*]vc�����Yz�Z�b�hk�<M`�&ڶS�2H�O��t���Uk2����w��Ů&ٚB��^YA˫F@ES��ɖ� �.���jR<+0dO5H:K:��1��郕�x7�.6�z[�x�B�:�:�#�s�����$D^ժ��KZ��Xʬ�����`�3��*f$��$t����k�z�F{�'v������ɿ��	�g�/������w�*�R\MZ@�����
�]ɉN�c�J&-��!���#R�joiׇ�y���|v]��>8�-f6żf ��H���#���ܤZ�ܤ�ˋ��^�Ե-Ń�$K��`�}ǥ�x�G���y:y:A Di�7�f��w�y�����V-�t;�kvm.h��J� �Y8�%�H&x���i���x�]���¡>�{ȁ�8�.S���U�}������R�3;��f�v���?s�����ё��5�v?�������� �=����.��	8�����p�R�rc�|!+	LV���L�	Pt�ε��UЀ�8Y]KY[�Ӳ���é�n�4ߦ�f�h���q�[~���C����1��	jE���l�=�����u��$�f�*[��S6g�B��~��	��kp8��9!�VX�t�'��MHc��r�����X�^��0k��Uk9�l��[A��G0 ��C�,x��/�54�0�$�~��$�
_��7�f�ߎ�P{�N4��w��{$��M:
{:����P]#��y;.|G�kB�
�c���w�3�;}�E�.�����:{�>1"�sbT�X�����qs{:A����S$�s�����Q�f'ݼn��^�"�?�t3#	y43E}�f"wl���{�;�u������ �t�l�~�,�+6YdK��J�ZTi���m#3�3_�dEm�ԴU1�JK[B�7��0֡�ú4W*[(�.a�<�˓K[�i�ꌵ��8��Hºu`�r� t��"W���T֢�p�Io;��;�]�yf��#��tS1O\��		��)	�s���r��+�6�t�=�*͇D�N��1uWX`��c	��yV�nB�>״Y�j��5��z�V5+y��Db!�[zg��V˲��s.~->�m}���wl����3'��7&������7�u%�W��-���@��!=�$�/|G`���H3B}��F��ɉy�����aH��y�64�	a1��&c�V�
{j��gk¢���0M�f�XM"���5D<a�¡13o<�Tg��5�O͙$sxUau�d#�H�$4��	y��?��z���\�%!Gd����tzC��P�]����ąz�L${���s�@)�A� %b�Ԡ��<��	Zt((�Ԇtgcf�$e5+P)J5D`���<�)x��G3�@��Lpl̄yx�g��+���${���̈{*���F��!��ϗ,!�;BA�]lZ.�<to��V
%�-Y_�����{��u_�߭�{�V�����f�b�(1(P�
�my䠱Ɠ��gv������؀x�9H�9X��I���&�9T��M��ί��ofV��#�fW��;�|��%%�����]�5�����b4�!{u'��w濋1�Q;��<t��pcʽ����V�H�&y�\��Xx�k�A�n�[g�,$���s�#n@�7�i��\�D%%�=5�f�/��(��JM�"Yj��yU�q*f!�� �Rf��xD�D̢�%�(E�Bu��)]�i��4�j��G;���m,�	������x��$��O��0C5��#�Y%Uk'N�\��U��jD��G�z�a�]7�H��BA'E�d.#�D4��iHT3�s�g1VEX52l�ȉ��븜�Y�s+ͷX2���c�E��Nt?�j�U_�u���3�H~|LA�J��qc���F��a�������,&<W�@LTUv�ʔ�{��i#)�Q��H�JC�7� $Ş{tFas���� �z�Bo2�d�05-G=j5�ͥs�ڞ�N�qʎ#H�iPV�f�u�M�5e#��o���D�[���������;Bm�\#�!�C����ue��K�#���$�3�+ �h�*��F��r�+�@�8��@VT�)��0� �|/z������b��Ѡt�J���\<�=��J��o�;,���)mp�a�pc�֐�h,�Wv�[���aA��^���w�~�K��Z.��*�3�
A��a�b���⯆���X��]�	%03W��b�,��ܷ���u�|�MsRP�hv����߂.��6�"��N���l��m]��u��:�1< �hEk�;9�g�J*�ٓ�t��/�4�H���r$�ΰ��S�;�:m������cx���2*�Zjw,F��@
z���بQX��4*6!��⽽bh@'0qi�B,R��.Y��]=8��]%_YC�0���8�s�kց��.�[���*��]�?7ˤ������b�G1/[�X�s�*	ݽ^��v'1)��k!/G��+\� BP$�I	� �'N��Ɍ�JaQV;��K��<<�\�Ȋ�t7
9���H�6UЅ]߹��&�б||Yw��JB�g8�	]��yp���:�~(62�T�<6{]�?������V�p���P�i�P�PV�4��Ǎ�l>����!�Ø��.^gj�i��5����Y���C�F"�:@R(M`�,=�����A����̃C���]��Fb$�vz i^;HP����O�<D�h�<s�w�:�pJ�ۼVt\TM�,�d��琇nWsMވz?䙑)]�2������_w&��z��;���E6�����k`l��������pջF�.� 0Tqj6j���5�=��YD��q �5Q�������q�$"#v՚x��r�攩
��w�a���P��B�m�� �X�i�U��Nҙ�|N}N�$�NB�s��~^��*D�z�~q�����l��̴#1,���]���6PZ,�R(�@�5-Io<��{!S]ۮ!aF��jb2��\6/�Ar#�q���=�wz*��Ud�s�s�u�c����b�s]C䉰YU��W�k���b�T�6dU!�J2ؠ��t��+�.V�y���ђl6aE�媄�Fu5�3V|t�*x��J%�A��t�+�	��k���~��������K�%c�N5ch��´����k��n{�ߝп��ۻ}��-#����������l/ٵ+�T��@:݃5k����p���fJ�8ECJ�ڞM�����%��@N���S�o�CUԴ,T�������$�I��Hu�*�O:P=�7�tVM��"Х�C葢ہ����7��^�q�TU7H�MK|���]�+V�%L��D�#��Z�Le
��eXL���)84ka(A�C,�C$�A8���1�ڗB�e��!����;�!G�����ݦP��IFM��ӗ�z�h	E�3�K� �F��1;�^��O��*"R�;��.\χW&��'ۇ������+�N/���	^>[��E�	��Hu�b K� as8/�^�bYv�=�Abx���-l�x�8���zl��ݴ���n�麢}\p���b�H��n_�������V(��|�cR��N���j�!�\7�ߝ����3.S�"�u�A�}�3(Nc����N�:���#���X��=�I�^_���F��w��5З�U�Mn��#�+ӄ){��t�׌^]Y)E)F|o�!QUVQ�jX5w���U��-rG~��S�iK�0\+(�)�vȳ(�S��U:+awlC�,��}�?�&YU��'�;|ɐP07o���ul���5�Rг)&�]E6��hXN�Б�,�az\81qxe2c��{W>����g@��^[ `�M�5g�X�SSyg��=Ө����6���I�#���"��\oM1�iL"�-�Z9\v�I^G������F���A2��U�xBB�$�3ϑ��s��xZj��N"�O��/���Y�>m�B�ct,�@��p	�G5��h�����3Q�6d�w͈�S W�_�H���MT82��^,�<�e�����цn������y}���$��Ib�O&���U6p]<��J
�Ra��A�B�x�A�1S�0�1Nes�0#Z�U��4J���s�bA��|�8���`vnK��D��:w�l�RI|/|�H�Fz��^��;��������{����xz��jKb��D竦�������ɚ���-�"����+��UT� S~(��G5T�p9�ƣ(����ų�cIW>��&drY�g�[W�|;22B�9:;F>�\yip�z�{B�����n��4d``P��Ƞ'|�l��b�O6�L��>�'KWΉ[Z�9����By^�!�v��W�Сt�<o0˵@��M��x�V�W�K���`&�h'�p��P6��_H+��rs�I�h�˰��&e JO���~��,�<l;��l*x]�	����!��Qp	����Yζ�H�B�T��k��!��ah�*Tɠ����&CMKD%��x-�L¢�N�	�:� : �<h�V"m,(i���d�� j(�'�2+&�<�<T��$�0Z�%�J�����}�#_��DvE<��]�
�Z#�<��1B�������,�;D5e~L�����G�##"��:�4��`&�O-T����<,�H��}����P[������Ga����G+YcH���"RTx��lR���=*\T5[<�b��fmZ���F�j�T�c��㲓�Oҝ�\$��"OT��������HH�(�D��IW�H�I�J؝Ո"����D�L��]�C��+�"C�<]yj[�����ĝ6'��DNһ������7��;�`��p<"H���·��f��c"�Ь��p!�q-B����@kj��<;4) �EYD�@2����rxD� ��P�/:����p77�A���:�!�8���=��.�%�=�.Ӣ�gGK�J����ϱ-Z�t�)uث��G�Sk%���	Y��$��3خz0hy�,&ņUC��:fG"E䟉�* $�\X-��Y��u�z�2�׋3h�ș)�,��r�:>�%����G�O�;�ߞlF�dZ�Z�����2���ćÒ��߃�c�%�@I��q��rg~o��8������3m0�ۇ\(�<TEvݾ�w«P%i��<o,�T+�M��Òz�Ƃ
�l�W�@��+�%EM0>yn;��H,���I��"�m܄U˖��D+��@?
�
&�'Qj4�&�Hl���E��7?�w݆�������OO�������xj}�I�-֬���Pޜ��~eA�����۰Tv�Tl�Q���h�I�UaGFY(1~�<�jYf��0F1��*�H��s�{t8���g+��	�R�@/uq�"ە�ז-vO�bQ�EchhD�v�La�	+�&��bAW0�b�+)�2^ac��;0��b]��Tj���d�dFl�� UJ^W�C{�D��u�L^��6�7���mBb,%��M6�p����%� �%j�Je���j��}�ɭ3Mr¦��x�p�����q	ip��>�/�F�@��Yh���ʕE2�W���.]���H�T��<X������� _
G�И�VόκI^#�S}�f5���n"��C*�UM�%6��	i�*=��A�4�Zqh[�3y�~��̢иG�pN6�H�A�kI�>=9)Nff"#��,�'�+��jM���*\�!�^&�m�K�{!ex�G��{��E5a�#�b���T���A��ݔɶ�w�f,�_'�N�D��O~x���ʡ�	����7`XN�'I/"ӺG`���d��ۨW���%�-�{�f ���fF,tH����.yaPr�\5�"--��a>�ɞ&�OR���4�vU
(zZqYN�N��*�0�]���(���&���Z�|��2�ӴIr���=��vM�v�!�
Y��#�F62��d��DBM�h�.�4�%/>f�9�Q)�˵�V�D���@"�Ed#kq��~K��ڈ:�#�FT<0��H<']�K�y#��J�I�����<P.�N8)������޶�v���{˗P�����+�j3�Rh��r^BA�*�?/�Q�|�� �q�	�a)~�*����ڒ��.=��2
��¬�H3�yv�s�%�V    IDAT�R^$�Y@��"ҤCSdXϏ*�p��(n�F[	���d���'IL�	]/e��)�:� ��ߎ�VPV�V�0�kX-3��>
�5�Zr��{ϵ��ɤ���i2��EA��!��J�2O���Gʜ��0	�⩞�4�lؽvf<��(�2He�[�}�y~� �T�p]ڑ�֚�D���8k��	��XЍ�������}O�>���Ll�X�AN���3!!��(�q1�ú�n�鳓p�(,��:.B��^&�N.:!)�"\�thԤ��.�����V��#�M�~T&���L����јLq��Y���ҁ'�ÝZxB�p���
QP.d\����M%&$�,a�
ՎZQ�U'��u�pu1�Po�Ѱ�C�N?�͊kTH#Y�C��=�/�ON��F�XZ����s��6��^�@���'�ٹ�U����2�f�&PX�'�X �d*3�RJ���ґ�H���|qM���8��IT*��)�+�2ePRM&�38��i�i�0����Â��x%�3������sÓ���$��5�Qi̘A��^�(6�	]|�u�d�������d4�ũ�(�3!.|�t�Dj.W!�q%�N8m	��b@�RFii-ۖ�%O�ucA�_��
Ẅ,pfzLݻ�!�Tk1 RҸ��>��1�����h�����=N��k�Bi!�����c��2�I<:xE�r�H����qNQ2^I�Q`+�o���rSc���č�π�lRG�4�VcA%�Z	�h��~����� ����u��I�R�k��v�&Sv��Г�!��
C��f6Ł�3)��T� est�yP*i���|���gYu(k6`���m�	�T�~,"OB��l(��j !d�0�N�h��
�KC�6��mQwn5eMCu��b==0SYqd�fc"k">���Sh#��1-��G�Q��Hez��t�{��󎼕�?�Y��xXl�jMP<�u�T�n����\s.;db���>.�C@�,mF[�<�!f*г���]D��=�ۂ����E�O�:"������#����R,;��Y��y��5dؒ���/�;������bՂ]�A�,�
���ͫ'R���34��<�����';"@t�=>�Q�B�R���;&E�P�}מX��]7E�.��Z��Mr�fsM� �S�޼>$3s�)Ƞ*�a��r�9�k2J�x���wV�b��)�j ��>A�k�Ed��t$���=]Lz�=���ͣ�j �0�f�2�9s�⤘c�Sg��m<���i���G�H���NA��߷v�w�v@&�9��,y`��?=�����}�CW7��,�-G�?.���8����#�z���4��!1�f��h$�a»�@���&�.L���(��p�Љ�-��4�Jk��.H��3�z�����"��JM ��;э�<�ԉ!��Ts�C{?�ы�����BTWӻ�Z}�$�Ea7]DC,�,��:f :�^;Ws2E���Z�ޔ��RZD_����oa��Ii ����� F�oB���CB����/& �RK��D�B�^��x��l�<��rx8�;H�?t�x����2Sd���������X�������;<(�!��n�c���xZN(,�F�g��s,J3���Ӊ�gH����L���&���/�+��H8��r�ӥ9�I��ra
��!0U2;�P�U�P1�FW2G'*28��JE,-,��=�T�� A,�v/^"&���d�~��l�X�*��'��^�;����7q�����6#N�	�R�nC�oZ\�����I��<Q��43"��dy��pZ*S��ی%���`�l2"0�����l��i�A>Aa~���p�P��IY��Z�,(r�<A�TC��OC�XԊ%�BI�I�v2�dT��p2���a�&�я�I��.X�#qV$#��r��V$�z�$"�A�fz�H�Pop�F�)���YP2�Ò� �C�ø��t��x�fHP��Z��z�,�;��ɰ�"<t笲D-c�1��,q����8����*C���0��lpRW7!�uI��b���(�捹�:�e��+�� R"[$S��E��Ƅ�d2^-YY�]D��i�Mҗ��o~�w��4��QȐ�-��6Z��p�K^���@֍�p|D�%N��&��g��l��P�Pi�dl��޲)���1��i~Q��k��(���4 �;�� ���<�h d(�4����d�澜&b��P���z�ӜE��p����od')Q8+�=Q��F߇�kh5h�TցH4��ŉ�h�jI1J3B���;�(ᐐ���C�����5K�n�D�Z�j��-��]u׋H<�������ڂ�p��'"W�A<J�rI�\� j����3��C֌`e�wb����y�]�������^�p�{���Z�۲��ot�!18� ��ظy'
� M'�H4%Yǒ	N'��F�S��XNJA�ًNqfR.����	%҈�i!�����Y�w�.2�����M�u& E���xg�J� s�;v��af�� �5�k�ad��	V��D�uL=*0��n��W��b�9>��_�����_i���+�hB�z��ۯ��.��=����z�߲��[����@�B[e�dCh�)�����N�dB���'$�����@9QZdzR�B�Ң��� -���T&$}�ŢM�7Q*-I  �!#��Չ��H��2ڕI@-N��tQ�$'��e�E��BO�W9-A�)�b�&�����0o���
��}񐏋��Eq�:��(���]�Xf�]9N~�Ω��BG*�CcaaI�9����$�I���V��Z
��Cl�J�D�F>8�<)��g4�á<�������ks�[�l�i�x.��-b�z�К�g���8�ɗ�}8WJ�#��	zK��p<���:W7�[��ڸz�8Ν8ϩ�T3HFzK���E�o���P'�&�Ωdwl�h/Z-U��1�LI��/!�	�T��Ii�b3�RBWbh:���IT;,lJ�x&�8�{ڭ��e1�0���`�8�'�1"�Jf%�}H�Y��o䵓LB�ˮ,�?_�y~�����q�b��.�	Q.1L��ؔk6�	Ss�K�P�Gq~RM�tzK���$;�Xm��آ^��a�L�:�ӱP��U����T&�d:��B>֝5�J�S�8�m��(�;>7䣰���<&���ɥ���=�@�gTl�T�Z	���1uI�S������@:Y6�mى)��c�����9S�x�j��8���{D�96l1��☹t��)�R9,�]	AD4D�A���Y
|��d�P�M���lO^<��,v��W�d���"ڥ��հ!dT���Z,��b��>�Q��I� �D�$�TA�����ފ�U9��#��E� ��B����^�C:׃��^�	�%��p#qx�	|��SdC�o�����m���߅��M�Fu��	ju���UA_ѓ�}ͺx�]�л>�7��������������ڡ��V[^V��I0R�tv��e���,_�~8�K�N�R��`��	�Q��4�[XB����ྏV݆�]�D��fZ(�;���f	�A�*
��9���_�|d�'o�0�j�b>baM z�Kx3Yh=YɭU��rjN|֪М��V�,�z�cˑY[&�H�bG�²8��H$M� g(C��D����]3�+̦�iZ"f@�[��2�~�I\�t
>ٖ��k�c�}����b♒.	|*�sN��H;�V�>���]`3�L*@�;l�F<��Y���@��Q�UzzN<�8}�K�)�ǨX`FQj�� �xj��^���:C�\����"��A��y�,�|q���dP���j"aq!����A�F�:�XW�O�w�F��͏P���dB�}ަ��1�r3�^���X�J�B����	y��A]�^P"�阍t`g�a�)$�*J�`RA��JB����9�:u���}�`r�)P,w�
i������K�kb�'�_&�&LR�h����\rx�eJW�i^���^C:N�u�X� �m���=%��,�!\��={�En��mq�A
c��\�_���%�-U�K6/$�����`�M/��$y����k1��g�R�!�J­39M=C��Z\e��j%��rEY�ru�5�ٗ��庍{WZ%GذR�lFDz�3Q��ux��DV��f1ix39M�tÔf���y�t"A��C4��%$�0e�MD|K���s�1~�B�-��~ۀ�Ȣwx5
UK�sa
tS�-���*0ħ��tJ�Rl�j)�&��aA�I~�%���gҭ��u�XH�O*ֹ�VA�\"���CO�2)�j�&t�o'�P �<�N\2'j���9�h�	]'���])�Xmԥ��Ó\^���I�CLU��鹨y-��P���̹���PI����U�QsL�s��s���I�#��YpQ,W�M��w`�ɷ�K$�
�Ra�.�]#�+
���s�CAR\҈Ȅ��Bt�� �.2Xs|�檨��gS�$�҉�P%��b��]m��,�P3��i(yFoٵ�h~�Ͷ��B=��&g`�䵍�¥X���xD5�bf}H1���CE�s���X�ˎ�_��?.����s�����6m9:/���V��(�=}X�~+��_N~$5y�p2�0r�����[b{׉�4M�4[����"��M!�>���g~��e&���f�rhZ=�ts�8)��%��j ���H�q�4O�+I^6�dR~���E���OQ-�
"�z��{��̤2�'��m	���2�b��͕��a�FiQZ&M�pD��J2�3p��x��'q��	�>v���	|�hŇ�
%d2�*��<@52����&�G q�� ���ۈ�1��1�E�G(q	h��1;qY�-�G�����< <�����Vյ+�h����R����(�N����َ��i$D'_�W�t�=O����d���x�5!LϢʘ���L�-p�p���^Ź:<����ă��ܯ��ū�� ���G�f�^T��q)�b����	����bP��q�E��?�I�/ҥP,X}��9�z��e!Q��-T\N�t���٫IAW6a��C���Ԯ�JC,\J������	贚�@��|�=4sBbԓ��}�0�����"|F��5�I�0 R'ɍ�@F"'S�G���˸�,e��r�0N|a� �����}��ܺE6�-q3FQ�(P��� ����0�U��x�+G:�2��6��`W�#��%�6�G�7@�qL1�}D:&%�F5�@��|��x��I%_�qzZ����� u:�)م&���Z.�Diٛ�b�z&��H�g��" w��e?#	`j6��,N���������=CX{�TZ,���B��QI� B�.r���bA��v����*�DB�7T{�5@h=�M-!]kG��6���qRl{h�+h�kR��j%�N��rʔ';�P�CK8�SIB��ΓZz���ێ��8�
���Ң2K���Dp^ �$N�r�;��=�8�m'�}[Чt&��J��nA;:�����s��%����TH!7���R�*�!��~!��jɮT��OqE��2�#'��B2�Q+@$D�H\oQ*k7Ь�ѨV����hv��jB\0>!gC�K$��G'�;�$dg�Њ�J�~�iar�rڳ��ױa�^�\�z�D��`$yD�����ȫF؃e/��ŏ�$WA�i�B���(������������<����?׽���@�V�	g�Q���)[S�ע�M���'��G$���7���CO&!���S�ҡ�
%ٝTʦr��Fa�a �D�S�������}o=���������3��9�$h8.�����"�jIB槯�q-��#?2��ec�Z.B:%��r�N��^�9�F	Ն���܁=w�/��E��d�jqiW��cf�:��f��780���0<��� l����NʋKbQ�n"������Ƶ'���[.r�c��߂���юS%���G2_rʐ�{"�F&==j
��[m�B��!Kԃ�5q��)�ë¨G*����X�	�Z7���t`�`F]�iBg|�����PX�<�I�}�.�)��g���~J��LX�����]����ʞ���@�rE�@8=����]Sq��uu���p�J�]��m���O�������q��G�f�>,T�Bd breÒeKQ'��*&�=�p
X�Z�HixjU	!Ag�{Ҙ�~�����Ԅ�ǭܼw~�a���Z��B��q��$|BN~b�Av/�*�:<�0e'��U�ϰ9LD|<��`i�<�j 7��}����Ulc��${�+g���RTNd�82�Q)FA8&����k�h�[�P6�˧���ן�Z�A!�F�
��s!��n �[2�ǘf�kT�)-o�
֌ť9b���IX"�(��Q-a��9��%T�����hrEK	GB&*"H�k�e#Ew6�Ӑ��A;M���d�-ty?qn��i�\�m�!{�6����ԥ�U|��u�"m�,B|�H���`JP��PÂnh�x��~�MD�&��ʵ�@�����YX���� ���r��I�;�MS�HFc�1>Ӳ:,m*9�J�[��w�����ȝ���p�D1#���j({g����?�v�+Ji9�/U����	�E�׼�MO5M�yW
�:H�N:�*���J\��qГu)��r�*��r��D�*�ڳ�g �>�T�14�/z��;�s�gaK+������{�,�¤A.��'$	e������Z�x��6�~Kޑt�ɟ�p/~���ٺ�@���[!: � ^��Hz�s󈧔�:��Qb�.\�az��xJ������$9�Uh>l`H�l�*��Od�^���!!ǆc	�D�a�{�rF%�[q`Dl��md�QY#�J7j���~5]�0Iq�	}EOn|����ڽ��}R�?����=65�7|sB�䁰:"�P�̋�I�l��\/�l�_c�Y���za�j��~x�8�^��ĥK@ˁ�J�΀Z�5�c�ƛ�B`&P#S�/���٣x�_
�ji!|����[P*Y0)	�CR�Ϝ:�+��b��i�"��ĒȤQwZX�e�oہ�뷢Ѡ�����r���ړ�i���m�����`faI�,,J�]�����? ���'�&dFa�I4+@:?���U�}�n�=X,�^�H1�Z5|�W�z�pX�S�|�[�e-_�CC��&x�sї���4��g�07��ɫ��e{r�вeHe��c�j��#�M���?�w�z�f�������%l�R��C���a�(�]���U��:��&�����Q��i��!���v����@π�~��Xf��n����{Q������n�\��"N�8�f��YUf<�C��@��r��\���8�|�dE��^~���_QZ�@.c
pρ�qӮ�1]� .D��F�ͦ�	�Di�naffNr-h��������b���h�+H1 ai/?�+��y�g`ۃ_���{Q��>��ˈ�����R�[f��IOB����ylؼ�D
e�þ��v��^���0{�#hN�A<�7������h5,	l�������5Tˋ�_cǮ��X��flڶS�*��9�0ȣiU�a��q{��)C���"�1q�'����0W�&-F4�Q-� ��ieZ�q�i��d1��aza	n8�L������u���מEP��������JdQ�.���Mv�������j�9O,���-B����%lmj��{�iL���}_�3�i� 'K�Ʌ�I�2���LO�����F�ݑR��h�y���ebHG����`��	
��`�������x��.q���S���}��E��\���:H�F�ʔ�XU��&I�3Q���ȇ]E�("����g��B1��
HВ6�d�5���N3��a�hۂaROϵI^$�9���,�->S&*�:am����@�K�E5�]��\���:�)�[��Գ����B��@�f��Ͳ�j7���q    IDAT�~���bfM�����q���BÏ�� �mj�e��PD��|ޘ�h�=iZ*�U���s�L�XJ�s� Z�F�D��`;>J-0�p��4i�E�;M��`�vq"v"�,�j:���ų�
�xE[g�E�)���f9��6��!Y���*��9�c�r,A�(����(j�-�,Д � 6J�#^4�g��1q�����d�}YAP9�r<�Lx$bGCrOW�f��[��;�/��6˽�n���_�'�g���F�At�d�N� �������L#��Ŧ�����aل��������(�������W`իش�&�[.�޵�+8v�CF/��{������M!����p�^��/e���8}�/�^%,_���J	G��+?Bcq���l"*�'M�K�*"�8ʶ�����������P��Ѝ$�aO|�P/-��ֱi�n)�զzA�Fo��,����U��P��ɺe�y(�ģ>[(�ll�m/����0Ri!�tebA��?�0��H�����h� 1@ο([mģa8��� )����Ʃ�6;)�0B�j���K���1�f�lލ�Qu���<o>�$LCGvhv�y/R�A�SiT
:qu�:���fν�c���ˇ1!��X�O�@��݋��Ѥ!L���Za��oP�����{�ǎ�b�{�g��^��Co`b��	ia�ƅ�g�8�=��>lٱ{���%�(=��l<�Ŀ�:{�tT�v��0��sUBk)I�24I4�5}�&q�������ѴB�rL��Zd�WBK�E�m8b�w��ӿ�W��y�[v?���e/ꔦ�d�����ƹ��Q������)d�-�H˂��a���ؽ�.y�\��9聇ן�殜A�^B��2���GN���HM�!���˘;{a3������p���7[�p�*f����>��q/��5'�#������8��k��Uh�+�U��}�{��o�l�j�<�&�Z-�Z��Ν<��kcr�"�''��f����5lRb),[�I��Y��"ߋ�k����UY�ŊMqϧ?K3P�i6�F��4;����(�q��Ey��}ɠ������rtuY��m�f��۟c��IQh�,>��_���IsJ�LT�Dɕ���g����iAN��
�Fz�78�M;v��P
��Q��l�Y�� �8��k�|�]^M��L�ӳ�x�K�F(=�F���:�W<a�W+%$�m�/���%���_zF"��W\�I�\>y��x!C���o#�D;0E6K����hs�	�&��0�x��M����4*rF�WQ�٨@������Z�Ajd7�܃L���ΜRY��Պ�͢�&�>a�\�B7��&B�mDd�K	��n ۶��/~���8�1����m8�зa#G`Ѹ�<)�V<����!D�D~̂)���@�!�F<�DiiW�`q��s�ɚ�0�b-�D
���h�S���1a��+�\��)]6 ��@�"��o"��xKp��tn��b�%��v4.�%�� =.�	#�@�����$zC�����1�
!hհf0�������Il�e+�lۄP4�#�N���uԚ�d��\�=��f���[���QA�������n��[�A�cA�]����4"�z<�F�z��<]dTt�I�\;�������z�ظavܼ�V�ęS'���1[��FR����	w���@�~����8�{����R�����%R=����je�;}�|�DT
"w��hR�n�q����l���E8��-{�­��G*ʨ^��wQ����Eq��}x��_���$���6.�� ����C9T��"�b���dzݰv�4\�^@jl9�|�a����T� �@��[��
g���(Ǥ������F5�C�
D����7����;8��K�F#Ț:�f�$�"���ΥI�իSX�i������n1Ԫb����K��]"=x��#$ B��v�MO��O>	T�ѳ<�8��xF4��DBH�7��J���r�f,۸f.)+n�����=XB!�t������`�XEoO3�q��!̜9���^�u#�ٵ��Y���8wy��2\�^�>l��Al��V!�5=Ob	I�5O��_PgAϐic�]a��{0_�"I���*Ƞ��g��{���8�\������LNa��ی��~
=���j8�}nsZ~V�^��{zk�ߎrKq�QG ��G������$Ϥ)�%�O��X��#c�2�h�!�Z�[n݉�9J8�ï?��'�C$ ���3�w������x���Q���p_V�V���kW������bG��x~�$��-w>���E��A����¥��@�+�������G���JA���ud��z�0}�
N>��+�q���
�,��Ξ�����<"�l�w7FW!bf�x�M,L\���<!�v���m��GE�	�Q��jbi�2&/}���N�]X��`s��"�ZD�@*�u7����[12�����D���G��t�o!�7��|��Di�b@s-8�Y�?q��{Gɱ��PTAN4n��H���|�뷣h9p<���z+�7p��;���+Hj�VS�E��+��W�
-#�F<��7�I����J�"f�0?7#;n�蚗��E���?,��*�X
A؄c�q���8���6n��W�榝hYʁQ������"��J�U�@���#������[V�5�4��O_�S?��Z�������~n����T���Qd���49���l.// ��Dff�)��T�۲��Z6rA/��(M_@��ZX��V��ɿ�R�3���.-$�FSp�U������ȹ����0uA����jsObu\������ן�����}���{@<? ��,���U��j"�)�<�p(��ª����M3�\�M�~���^8��t���E��*�
� ����96׿�$lJ�%�'$Ѹ���2A2@���1��E��x��1:ЃG>�)|x�8B���+���pibR
�	#bh��2�ό߾n�w�v`��m�����_:1;���KAr'k�$��`���N<�������t3<�}�gN��]�у����oɔ02����x����?�E�V���q����,ar��X�7��'�`*ƹSG����DN����K��G�s��	��֫�+E�Rqe!�9�m��_�N˖	mrj��N#ˢPo!��c��� �ӏ���?�P��E�H�{p�C��@���>�{o���SA>�#��ޑ�Z;w���+� Oa劍��Ñ�.��a9!�����Ь6`z�p���)�K��|�k��cB��e�v���q}�M��	I]A���$�v�ۑ��a�X�;����Ea����/|a=��S�����W���0���_��� �^����W���)d{Sȥ]l߸C�4.��(�X�m��P�փ�EK���	ܼo'�VYv�/��'�Pky������q}n�L�=�;�|t������W>� V��1���W_Ǚ+W1]wQm'�N�bq���{�c�w�E��"�:0/��G2�g�1ay��!���.L�I${ۅ4a͞�kO��9�3�Г�Sn$v�-d�)�p-K�&�k���G�͡�Zp�x����X�"p;�2V�r|#���X���c�p䍗�%�F�8�vY�+(�!�F���՛�ۀ�O]"ۧ>�e\��G_>���{W��3�@8����%�L2q/��IL]:�Cy��2�Jw�M�:۷o���<.^G�n�Rn���pa���<��7oG�VA&ŵ��p��K�Zeh!�T�����美�[�c�L/��e�\�po���� ���o���ۓ�h�7�|���M$z�Q$���-�߃�{�B�RG����i����"���l�� n��AX��:j�����`'a8j�͘�Z�%����)O�08<�O>���^4B�L�o>�\?wR����(���O�D��lTù�@cv��ۉGc��5A����|�@�ր��E=0����G�������f3|�}�z�E��l4j�QaA�O��p��t1_�t��l����e:tH���<��I��8BX�n��%��W"��¦M����Ի���~�T�-��{����i'<WG�P�P>�ReW�_���g�4qIHWh�ҋ6z��Mؼs?2��(׹���N� J�8��s(�M�q�=�b����i�U�|� ��®W11~��)c!����`����r��|3V�� V*fZB,��C�z6����Q�:����v�b���ɿ��N�EdϪ��)J7�h��¥�h�r��d$F�ЛMc��e����AͲ�lh K�Wp��gp���<��ȍ���<�T�� �,~Cm���h�fa�q ��g=��l��9q���$��ĵ�'��o�P�v����-�߱�#dT�k!��U��#�A%9���5"�DY��������!ľ5)L�=!h�C܃�?�$&�_���UԚ�8��*�\�Do�}kV������ek��v�~��_>>7����{��%���*T@�)$
Sɗ-_
�ƭ;v�O/��&Ν�񃯠8=������{RH%����;�c�v�z��u�^�[!����8uv�����ݻ��gp��a|�E��9�x��?G��0�'���p��1���p�����a�a;F�!ƥs1�/K��I�>F�n����	�]8�w��
��hil޹w��)k��]|t��غ�v�$���U,_9&�~�AK֪�ؔ���b�D��e�X�}�ф���s��'p��aģ�����<��o��'�I(��bi��{�g�=�o݌���5�B�!�vx�FW,G�Y[@��/a����n�v�L=�C/�V�ȉ��x��� 9��w^}O�8��a�ͫ�K�Hxf'�Ĩg庍�+�p��U�c9�zB��("ɨH���_����H�ӏ}}k�c�\��#Gq���O0aap �O}�N�z�&.��AX�l�ǩ+�X��Qo��&v�u72#�����U��KO�%)�x���!�ۮ
z8C�k��p�����4�ؼJ��+��e�� C�����b��5Ĳ�x��y�[aD����/~m�G}�2�����kh�|l��Q��y7fJM�R	h�I<��"�4&1k��E6Ff��͛q��Y	��Y	/>���
��~��ѕҨ������3�}x��Fv`�=�U��\����C�<��#}�el]��n� ��B�6n���4-"�/>�
R}�(�!������9j.MB���N��p�a�� ���>�����|����p6���I���/`j��������Oc�M�~��1�����
��E�Z\���ßÆ��96�r	/>���?���SX�}�������OѮNa8B*�aê1$�8~��K���E�O`�0�R��ͷb�������<���BDo#�7�_�+h�z�	<��c��^|��=(L^@�����Ә��;!055#�����pu��%���^<�w�7����ȳ�5p�����Ы�G)��J����z�?�N#��������9�#o�3�b$�F�a*ղ���-,�P)5q��b�]�@��	�����{���
o�"��>��ȗpӶ��䦓�V����N]��8=�\�T�4TLsl���5�u�ܼ�v�L"Bݲӄ3?�����%�}ش��?� ��&{�\>��k��;1{邘/������#��4x!"�;��?�y$s}R��pT�8��
��g�=&�!�`�ŪM�a߁o�dE���#��K��a�L���R?���5��$�*�Gh��}`ho���C#�D�fa�?����W���?�)(����[�wp�&&����7�Fia
Vq��{��yQ,�j�iy�ãشs��CH&�X*W�j>҉�]�s?�!�e�Q-���c�ν(p��6��F�䮺�ٙ똟f�}A�.l�7n܈D6��ec���wV����N��HX�l���)Ͼ�;Tk5|����R�{�hL����<��طn�w�~���vA?5�N|��?�ʩ���j�C7
:�\�U|t��[.�Fưn��p\�s$cI��ʫ8���h�
�y�j��%l۶��-ǩ���Z6�'^���~���A�G1����ks03Yl�}+.\8��}Zv�Q#�/��H�3�~����Sb��1��q�.�G:���r�̰�Z�&�ʖ[v�Թ+(�m\/��y�m�����15~~8����?��kW��+/bif_�Ӹ}�f)P�s����/����"RLQ�[ĚU۰��=�ٳ/a�P��[w"K"��������0��	�ڈG��-8�����,�x�^}����C��Y\�pa~NqD���zxl�8`]�x��۸���b�@��%�����I�[�"u��
x�?D6�f>��oY�d��6m���zP�ԐL�`��J/_�����q�S	D�3��)��E����7���<���Ϡ�u��'��{��Л���,®�ɯ�la��;�����ӟ?�sWgq��l�s��������8=���27�t:�j��wq�Nȝ�&�f���O��
nZ�Ǫ�<�/[��?8���A�oߺS�p��q�-��b�/Oc|���_|��#h,���'~��UA��`ӽ�ź�wc�fc��>�L]<���F��/�-cC����,J��%����K�tjh=�����w�b������^{��8w�=!�����'���H���۟�P�3�eM��~��.�<q�����������׿�G���W_����W�a��ز�6AeN�����E����y�ܡ�q�a��{/��@��F����?Aua�ɘ�߷���P�X��<�%�&�L���Yy�̗�e���=*�d�m/>�4�|�|��Al�}��	;���A��jXџ�M�"l$��^(�05W�#�B�$����"n�ħ�a����p��ui�c}˰�O�ff�?:�Ӈ^��������K��JB�{��w��)T��A��ʫ8r�$�d�_��+8�+M�|�g"3�Hx�=G�ފ�D��*��wO��ݍ����ىؙ����MwW�J*y��(zR��H�@z���{w/�p����}��<Kn&f����-�E3�`D߾$�����gZk��D��2k#�">��#���fx��}n98����.�������>&���,ɽ��Mn��l���&w��A_��ӣ���)�.U���~�5s3�XR�df�QF}�y�i�"Ic`yi��/k-��**�7Ҳy���������?"�u��ݱ����Z�f5c��Ǡ��w�y��р��`Q$D#�!�˂� �
�� �[m[w��[��""B�+�B̧�����>t�AU����=��6�F��QID�ܾz���7(�K��<'��� ^��ӭ�N��ݽƒI^u#um{dR�-��5�:�-]���BOzv.o��B�͡3���@o7���'��mz\���%���i����jJ뚨�]#WrQG�$pLq����WHO�e��Ô�]�\8({��O12����8��j�*	z=���`_\�+5���_�JNQ91�X��xc��ܤV����<���o�HzN&�M�\�y���=�#�9�7U��]�������_��<;�?y�k��C���]�	�ž������ �d`+�rd���M}�Z�QQ�1Ƹr�,�c�X�	�R�dg$K%�Z�"�J��D�&��fB�cY�*�����Q�td���5�L�q��Y	nI�(��Wߑ��ٙ!:;�SU�OU^VK
���DWB�߉�|d��ȕA�/z߰���6ZpE\{�ɞ�/�$��K��2Ѵa[v�����7��e�q��V*3(�ˤ��!��L	�	=d���\�*y��Z���YUCEC3� �$�q�+F�< Y���^X��#/��0)hu&�a�Ξ �����W�`5h��czrT�9�:��ދ_xL	�/^���}r6�o��z�6��U���y�_=#o*k>���"��;��<�5u�R,Ilڴ���IV����	�7���R���u+�@���Jl2��w�����MjA/����nݹŽ��)�I%)�dҐ���-���    IDAT?�ƠL���BB z4:�$�jH5��%��݋��m�RҲ�C��ō�o�Ś���rӸi?���Z$�T�q������d�<���	ov�N���������~���/ŜY����'�6B�tv��KԽ�Փߠv�p��]�)kق/�C�p�ˏ)˴��FX][D�EK<$��~���6���&��"�^��䌍Ew��������񭋴߸�V&ɚžw�
�����c�Ϟ�f��2x�I~A.z�!l�&rG74�Ϯ��)/.������d�$�Kf���eҾ��m�o_��}�� ⏲F�;q� �\�`�c;/�0�x�ki����wc�Zj35�l�	�/�pB���gٹ� EUո�v��>���!�Q���݇^frv����Q��#0���uul\��`� 3KN
�J��|f,S�Yt9�^������9<��_�T|��s<��*�!+�/��5��|�&�H���{/��ӧOJ�G\����N4�"{���K𠫏��E�8�������������޺�E��1���7KT�F@t��Z����$:�O�I����N��u-�%�t>��ɘDII�<�g]|��9�*�^~�̂J�Ifݾ��@��cHֳ��7)(Y�����]���PY���'/W|~\$k���u:�xX�;(�oe�ex�C�V��*1��������)������1���h1
3X�D_��� �O��W)HNA_'=��LV9�tG�~�C�lޱO&�E@R��"�����T]��rE���k���n�� Y)PSZ�w�������2՚L����b��i5��)��B�Q6<�*y��҆��z�s�}�7Qj�dd����o�2&�lGoo/��fϖ6��;x�q���A���*)%]RI��0�R�f3�7�0	�x���'���y����Q�f5�xH�܃�ܺp
�"��>Ϯ����[o�4;�͛7�p�
*���'�MԷl��rZC���*�N+:�~�{Q����5�$W��v269I{�"�5�8��E�}CU�_�d�<��礸������䭧6���NU��[�x���4��R\�$ _P��aRӳhln!�>��\=^��Ł�����������IOS(cd�Zd�R��6�$+9EU���tU}�ܹu��I~q����W/ۦ|r��M��m\G�5�ѩ��G��N�?p!�HO6���t���/�a�aQ��2e���g1?;GT�g�]��w����\;�=�T#��4TQS���P�$Ref��t���J%��ڵ�l�S*O��R�l\�G������<��Š���R\��s/��(�z��9~<}��w��뛩*ͧ���[7����-��IҢ��q�=�E�&�}r.�]�B��Ζ�-<�w��7����Z�O���~�ۯ1��I��HOK������~�-f�G�q��g1ݨ.)'����y��ާz]I3���Y�[@c�����^XS��z*R��d[��7�0��.	Gb���K�YP-�*�bzҴ��os��[�%=7O&S�����xH�&��pҴa7��]I�HӉ�v:.��"�H]Y.;���y:8�%�*;���%B����PY�ȓ�)�]��/��O�#�Y��w_������=��\�M&����q���$��2ر���RL&Х�3Ye�d��)��GF5�\�)�tv�s�����R^}�%yC�sI�F�����,��8�-ř&�<�KR�\������rհ(����3��/���<�����XK*ɯ�&35����t߽�J؁F#�;q"�-��P�v;N����N~�	q���:Y�)����Z�b�J|�}
:����e�bIɠ��{N�Ͳ�M�W�����͋gy�id��y�gƝ������\Rq��Kx��!�Kv,9�r
�e1a_rW
k,���GW�L/�ܛ?'//���?���.�X@��7{�%���~D�&º�T���Bu308(s��9QXZ�cҩIOK�����O�?���a�ٮ�_X$3-�ގ�<�q�,óM\�G�V���KL��W��:��i?��
�h�(�鴓��)�۶�iKs�>æ�t��`�F�X�6gr����p��5ܼ�j�%�]��޿!-����1n^�HZ���k�Q*C$$�>'#5G�IQ
����q���� Sv7�k[)��#l���7_�]^$MP�n={_x��?ʍ�g��V���:�� S�C� ���lR,V�;:e����A���iL,/{�{�5�|s���Eɪ\���	��Ԛ8�Z�j#��OP�����McYk��eF�������WV^��
	���,��$�\��	�Kf�r�hl�Liy�:%w����u�o�Up�����k��������u��_����lB�e���ʔ��s?^b�攻t!?Yv�1g����Q�K��4L=}��O?� 0�dv��6YUD�	���8�-�X@�4�J�/~�K�mh��3g�q��-���8#�%#�n5[�&;���TI:;��F�p�#lS�`M7��`��
���)�C�m�]E��Ѷ�ҿ|wϦs�@u$,�Ǉ���8���Lщ7�HTF�EUK-(:"���]�D^��5=��խ��.�'j#��^e��	ue�ڻU���G��ɲ��j����������Ie�f��K}
qSWۻ�߸�ѩ	n\<#o U5u�����`�����y���HyE	9y�tvv�p�inl���U\��@������oIy�����������X���ջ�����\�~��䎤������K���n�rs��V�� W�1N�XH�䜃���Lb)���z�rѬ��v�3>�4 Bvq=�^�Ψ���<9Ѹz�{8��,�����yRRS��͒�s��W{=df�J>����6l%�4��~�EPkd��tܽJ��sr��[��˯�����ˏ�Ʒ@KC9��8����f1'���Go�H���T+bJ��.IPJ�+����������7�O��o%a.��W�~���JN�<��`7�5%�5W26҇V�D��L�Y�R0�#>9ʷd�16>#����k�x��k�C�޶���|�}�.Ω/~��6Fr�
����[к�0s�ii�ܻƓ;Wi�)���P�TD &//G��2�se\#z�J5��=���ޢ�����E�M�m�r�Z����� ~_�u��Ӱaa��مY��������O3��W�03����A�j�����L�^%ȥ<������q��#<|JjV�����}��+gI;1��}o�
�?H�tq?�~��wY$3ҭRO)��.D)�dlL����W�b\��?�2=��[�cQh�����A#8�^����¬޲����FR4f�^<I�>�΍Ͳs���1�����z���ܜ�7Dc�:�����5f.���_J�_�A��H����������[̎�� ��-&ų�nVa)N��N�2�F'nξ8�`���tY��9ݜ�v���մ�n���y������`b��?���+��RSĎ�2�l[�>�����^������S(��"��d[`nq���z�>y�)���zv:���E����4��WIW���D�b�*e���%nȐ;�$\:�G��a�W瑚�aζ _��yK��4
!r�-#C#c����(��?6�|�Mm[�s�"�O��p������^y��Y�&?EICu!i))f�b��pbRf"@B�RU�q���9�x�.aU�*B�6�~�5A��@,N�V^z�]:{���e��q��/�ejr���Ȱ�I*�k�N��"!,�5O�?>%ء�!7�e�^\
��fh\���'��*�W��Ѳ�5\A��V�Y� 87����4��?^`rjV��Z��%R��23��2Q����y�iھ���k�����<}�@��b����*���N:�^Ǽd���ҝ�����q`JJb���dr��M�;�%tivΎ��f�Fj�o�� ���۲ae�1���Gߢ��I�<E�{��M��Ҩ�,��W�135�����%���/㏁'�S��Ũ\����V��
	F�:�1	:�]Cq��	˳��@4.��"X)R�± ������4�ZW�?۽�B ��g#�nW��_>���.F�k�/d��52mD,a%��D왭L�b�0���]F��&�7!Qݸ}�2��)�uj�{�e2,��"բ��x�|���cHJ�G'h^��Iw�Αi�7n����g�'�wQZ^��W_!ɒ���8����T3UuE���1蓘��� ?���t�%4�z�Ƅ�iڰ��Z����og�i7���#Ks���n�ͦ�����ύ$�Ӻ�����TW���}	��()������Q���?~�KFN��͝�Ӊ2� ��,C��s��'L<F����G�*n��kﳒ�.iSa�<�?�G�S�4V�Ѳ����֨HI�`�$������)Ib�D�H�����<h�n��[Z�y̙��Qv��m{�}�It�������;G]i.�9�����1$i1[�"1B@��)���� �5M`H�k��r8���۰/��~������4��Ȯ�/��'_0;��K�w��zN�������cIR2?;,�WƤ�$�<<Ӵ~#7�'y4:O���T6���e�S_�#~�,f��^�l���-�w'�$[�u���n֬���<���b�^�Q�s+**$��`N�oٶe;A_���z�|���9/�زs/����Cԡn����{iܸ�1���1	�Y�����4�:v��w[$ow�4(j|A�Kn�{�/����ڭ�L���U���ܺq���.aV]@2���%S
g����t���Q�>��� ��O�ɐ0 
4������+k�wr��SZ=;v��M03:��߃J����:c��(h�Eh%	�ZǽK�	���۟����`ttXNl�IB�SH��.�K�p���Bfm�?q�eo����#$���X�F�Z��~5G^{���a2�z�J�	L=aqj@�C3�J!����)j��1�fvlQf^�Ks��(���������u�m����g��j'���W�ޣ������=����(���uD�QT$�f�q10����,!J��L��ʌ�'�b�_B۶�x�LOn^����Q�|��h�PZ
����I�,&��`P�p��W��Q_���S�ٰi�K2023�D|n��q:�ٴy+ɩ��y���R���#TԷp��K\;w��7.KI�H����_�K�r��y� %��+Y"������l�}�nu��2e��N��G]dV7r��QV�.N~�)�S>g�[6q�ţ<�igb��K3ȳ&�r�$$LE�T�e��F`���$�M���f��"#���-;ɮi��tc��9����N?�ӐPLG��m��zD��u�(�#}(�6*s,d�'�q��m�`2�O� �d����IɤXt�����P���ƶVɎ�y�K���2̼幗� ��3�s������ܿ~E��V�Q�'�YY���-�F:�>x�̂����ֶ��c����=�DCr
[�%'O�r��7���tx7���������K�oD}��i�:n=���0esJZfy�l���4�@���j4Q:�o�8��!���/I ��(p����b�j�3?ϒ4�ZS�o~�o����a.i����^�;�����?������$kb���5Q_ш]��E$�_��
��"jW5ʃ�d4b_X����,̣��y��(�����+2�R�J&(�NQ�O!��{X�~�xQ����;7�{�<����y������@� g��J�7��Y]Ozj���	�`uy���ɷ�Χ=d�S��ߊ��ʌ;��U�;�}�������<ȺM;�-:�v��3�l]�H�EGUy�#�赂٬'+%�J<����$�2hn݆����>��7XQ�Qi%���O�H�Z��]����~�yK:l�8{B�{V�QQ�+�C�}2p�b�J��� ��e���iIGo�忟��֚���[����� )V;�º;p�]ܺr����lY�H��5�&s��C����`�5/;��s�BYa%uS6׺���杻�����W��ߋ�og��/Q���G폸w�"m�k8��fƆ��?-�Hn�	����T�N������NNiC~T�s�M�F!�L���������,D��wҲ��LǛ��<�zA��74�b]c9W���q�c��U��MM�����̼��-/.=Cuj�����g�]���Jp��%�J0�۶�y�f4f���O~����$����t߻)o&Ii98}�CoMB&��*�A�j����	]�#�WӶa׮�f���D��R��޷��5��kW䨽(�̫G�Q^��ן~$w��? �ڢ>$�]=O�ij^#Ii�:{h�"��������L�s��		$�rϷQ���k��� �У^Q�~�<)1;�64K����$��6$���㔕����-�e������%����'g��#��$�͇�LA4�����_&
����tm������^��Sk���P���A�e�g%��ә[^�L�Gc�-y�?p�������Va�9}��8�!Ν������13�}���5r"�0�cJ�̟�<�``h���r���m��Q��B�ƭ#�`&O�^���eL1��Ȅ�/ސ��w�
�Q��-8f�xr�,�Z�-Ie��1����rt¤#��������ts���X�
�T��r�Q�eu:t��np��w�e���;�Aa0q��MB��W��黯>�jb�Q�t�-�QE���>��5Zs�����"�ݕ�������%�uv�e�^��ƻ4žu�lX]˕K�eCB�$Ӭ�$��13� W,�P���ZF��?�GmL�e�.�kq��_"��/~�w�[�o�k����[x�3����4���/�z���	{�)�$3?Q_�ɩ9�IIK���38���<)E%lص���.|���;$Ȫ�~-������ܩ4U��}M����O��a%	axc�+T�q���K�9u�2��<���Ϧ�Ǩm�c~�1_|���A�:#���GUM��F�S�m�g���`򋞹`�����dUC3�./O����dlz�?���m�ʚ[�E�](�#t?�C�c��[���A��piQ�t�<�$�Ք���{�]����Ǔ�����X�D��J��q���P�	X��+�ψ>b+��"`�zm_P��b��܋��tK�@uI����X����h�GOw'�D���,��~�~���y'�e����q�K_.G�����ٿA������Ξ�$��,��9�W�J�rO�V�3[�i�cht���"*���dS�j�D�?�;�G	��X�e/m��K}���<i�OEa6р����27=��>Os}-^�Sr��-��&S:���T�nc��c`\�`D�O��O}��@'uw("�ï�����̬\��d-G��j��)�I�)ș�qj�*��ɑ�b� E�<>Y�ٿw/a��a�M�������x�ִm��r��q|�1~����ڝ�	�>}B�n
��Y^v;5��l
r�X�w���@�z�Siٰ���Ǚ�?��^"���=��{�����_QY��/�63����m��e��[�`�kuFTIh�2�
opTI��<=����Oqx�$'k�ࣿ�t
=J�����l�������������S��B}E��Erok2���̐#+��+�e��#�"+`_\���OW�{�(i�_~�������hٶ�������~�?��*DE���kWu,�Q��7�֜�Ơ��sc2���U�+y��G��(m;�����������U2-I,�ü��GfA�/_dij���t�2-���Aݿ���YY,,.I`�ťff�u�^�?u���y����(((@��˗OA\��:�W] ��{����0���7���g��3S���"��t+)&�\�%,�`hx�E����J��(C�S8�!�����i���3
��T�Zǎ�^fz~�ʒ<67W����)��2r�p�R���lN<�I��#%#���]Ե�`����=}�;�/c�0F����5q��s�}Ky~*;�V�0�Kv����B�]��=5=��j��w�r��X� YWt�dt�U��Y�as�v23R�uQ�)J?ѐ�e*K>G���DU���4>��Kgh��a��&|�9�?�u]~�0����@��z��PVUC릝��|��9:��)�Y͡Çyt���    IDAT�7.���s�Fǋ���PB��+i�)e�*��#7��NM�&#��}r�	�H�(�oh�΁q��f�����+|��	��C+�o���M[�w�1��67ɬ���.�*ʤ���pRVR,w�?^��%5����y�;J�ج��<�<��|���:%�D}⑴*bzj�mg����W�����,��׿|�ɡnzK���w�S�I�X�/��;ĪCIN^��78A��4+:ۏ����s�|���{RPSR^�����$������J�&JO�MҬ�X�z�5Ue|~�-V�i���Ѻ}���˒+F۞#���ej��|��2��lͤe�K�U6���!�M�$+�-�|��x15�*s*��f|j���y>�IPV�Ď��I�J/��Qz:�r�I
��Ԉ���@H��j���7� ��ān1���*��_��q�O���r>����u.�Y`EiT	ǅ�����{�@C\�U(��!� %������!xXZ��ε+2<P[V(���ZV��;��%��&��Y�7�dz�Òp� @濧f�UX$�Oo\������LD�Z��&9���۝t�ߧ��m�5d�)�˓�H���l"�R]]-�Ss6٫=tQO۶��%���<���Hۚ�MԷncׁ�.vr�gN��i�/Ǩ�¼4)�_Z�Ǣ�SQ[M��9#,s��s���z�6Y�Z�d�Nv�o��	�C���Qr�)o��7�Ǎ�`Y+�>�˕_������4��S�y�dXS��N������Ԭ����#8�
q#w::�8P���?���k6�u�!�	a�
��g�gۆ��߳[ڎB��D?�üm��y���x�$���bp����ַm�>;��/>���@L���<��|#���>�bT���g[kM�p�f��k���@�V�1f\ѱ�Ya�����F�k��U����9N}�{���E��R�n�<З���i`ŵ�7�{�
�)�H��0���I^F�|�.--ɀ�9Ŋ�㡬�L��22����qi�hX�	�2�7���c��ϪM�hݺS>\E���sL�=�.���U����FW�c�C"�v㈄�\�R�2ʸq����~�=;�{s��'����eA�L��o��m[����?�=��$�Lz�E�����f�e�=��H�x�\>&f�q�"�5���E�TbJD������~Q�$����}�m2��W���^�{��a��U�i\ENfC��=���B�е*�sU�)���%w�i�]���x�k�S�Hv|:3��ʹ�>���'I�"�%)<KA����n��SR���g{jbe<���jfYt��y�_^��o�����w���ف�j�I���7�:�n\Ż<�[/�&=	�'�$�L@���[-x�QIe�y�{(���{>Oai9s�Kd�'����\¢���^��2�~�� �2	E0 C��9F��V�X��f�ɗnZp!�	�����e7�u,���{�L.y�*�e��-ܹ|����tF�v=��������U��8튟�w���L��Ċ�5-#��=�2\[�����X���^9���KD�K����]�R�ٴ��v��I�kʳX�藓���l�6�D�J�Fì�!(U2a��p��C����LiY���Ip�����viU��LԷ�e�+8�!I�` }���5u�<�GJ����RVa�г�/,+e"��_X��]��08�(�;��@Mm9�N~A���h\���G��a�I�����L�#���%r�733�ŘD�%E��*(%5��������L�)iXϾ�;�Mur���\�V�b��c�d13>.[(���T���I����μ�,�_\"�P��[������Ꮢ]Ŕ^$�4 �EB���u_�����p,�B��Z���]�r�9VC������j����@�^����?��3����Ơ�k|��8�c"'���@�hqC����2�O;Z����]�޿'?l�dZ�H�c5iI�)��"٤������fzGf���}E�h�p�Z,Y�rg�{�&W��L����#Ǩ߼���e�)��`��ŹbLh�R���:��)<���z:�R�$��W��LAq��W{'�}�w�m��bZ��c��Ä���etp�s'�C���xaa&EY��'Mj#öEF�m���hZ�Β*�v~����D�8����h�1<�0y��y��$��,9^PKؽ̉���>�*�;v�c��87+�Ci�,,��s�!�I�Wʝ�#���o���z����_b2�I�.��_����q�?�0=���{%l!�Z����k���/,�_PA�!��2�Ǹ���b�9,�@3S�>�=Ks3R��q�*j[0Z��y�+g��~U%+� �%e��f�!�]��(�����L��{�=�apf��?OE��
�@H2��Stx��$aLLw�-S*u�@�}���R��*�3���1?9L]i;��ʗ��bᐤM�]N����q�fX^^�c�I����t&��tq��/�/���z(_�����[���[u:>�o��mͼ�ws�}T�� �Vt������Mfv�#�O0�us��W	%�X��8�8�3t�����s���a�2����lU�gɪc�ICc]��;8].z���]��)qㄢj7lB��N8�']�fnb�O}�:�Cs�U
;��M�^&�~��V�~���@�6AQN6�W���'H�k��JgqnkZ�之���N�܌�̳��#T��efb�[�N�]tp��nl��k?g��亠9�f��\�ލ��?�/s
�Q�A����5a[��;2ƜÎ���\�@/�N|���8N�eR*����a�d22<�ݛi,���M�f�<r��8���df%%�j�+���y�{��E��ūo���xD�F������^$i�%��:c�� �|�=�,�����~�/�Fba�lʈ a����=���F�B�#Fݦ�"�$n<�g�梩m�֬���3<�}Y}D�m�4�k�ҥ���	��ވ}~T��E(��\&+'w@8�b8=KR	[Z\σ{��}<�&���C/���̉��:	{C�my�m;�1�m������-=�|�ZL��.��l�s�d#��(�oF+1��މzFg�5���O�-DC!,�8��?X퐗���H��]���"�@�^�q��Aq����>�jKQ��b:!�Leiم/�/�´���d�@��ɖ����͵���|W����}/280F��`�6F:oS�c�p��Q+��T����1E����O8{���<�i�s�~�7���s�}z�S�|�"�Ü�Ǯ�� %����Nvmj�3׃&$#+Sf\��2%�^L��$5%%�E��Ԍ&<y���װ���]�K���Ƿ��ߣ0�iT��u�gji1EU����|3�bx�Z]��_��z�O��������D_�)��DHPឡ_�U�"(!t��D��̼J**뤎N�O�sX�ù�L���\��V)w�j�'�QR�Cey۶o�xF_X����)�TvL��0Өd��m.}�������{�-���-b���rD6��%�eE�dX��"3SH��C����BJʫ(���,�H$�Q���+G�ͻ�v�N\���d�Ozx��o�nj�������,ؙ�yyC��+��a(+����R��\��1DWd'���/x(S��p�ܪF����\JR2󈅽h�q��Ƹ|��z5):-��r��l0�t�$B0 ���(�KK,�<4��@��-�Wnժ�y�ۗΐ�l"�3��O�ǜ*��a�>��g,�Γa5�eRȷ��t�r��F�d^f��f|��2%�/���FX<,C����"���-{PײY�'D7������<���@Z�2L&L�5�l�Ԃ�b�U��'�|��i�j^G�V1>��fRq�8��GئG1'��Mp�7�9�=��c�4����!N|�y���ZMT���i_�����E���5j��M��U3<<�̒��D�G��0'O|���8�H����l�E|�H���dl#���c})��F^�xANN�*�����T�Ƨ������T�Ӳy���&�!��C�?��Ќ�덟�]R�mn^�)�c~bmL��B�m�f��mx|n�?|�ݮn��m_TIm}��kY�	ǂd�TL��p��q4	?�[Bzbq5��_���03��&�D���vƞtȟW�)IB�B�e��ҩ,+�63'�9b<9������c�+��^�����7_�<3��=�5��a�Q"J5sK��w�GY ?UK^zz����Yrre�]���a-�c3�茌�͑��z��o�CL*^c���^���;ƴ^��_��U �n�/�eb�!���� �p�{�.�{I5�h�������+-{��O��3�`��c���or��2B��Kt�>�I��q�CW�sy�Ϳ M�d�{E��ecr���u���r ��"��������!�(��Fo�d��܍$�Z��!73��;�d�S���ky��Ȍ�Z5Քa��dW[X�D��X@g0�>}B���
y{�4Lϸ�c��y�v�o^��t7�N}I@@UBq�6`��#����]�li�47���\N�P�$��0��ݸ՚&U��#3ؼ1��tNPմ�֭��*�Ģ��?|�,N<��0IT������ /��D���^
3R$�ܤ���I�s/J��&L�,P߸���R���|�����.��)�m��:�����Ǭ(�4�Yώ/�����bk[���ɞ�y�CR�)�Z)�ءP�M�v`����嫌�;������;��i�g�HI�F�����oP��F��Ԗd��,��a�o{�Ӂ�d�0���

�$��~uws��[�լn�e�N<��v��+<zp]R�	a�r��AK�8��5����*VD��{]u��lϖ;z�>�(�o��g��J�.H�1�H��#a4+�5,4"])t�����"�����hyF�3�	<�>���k��B���V���Kj֯���K���ҽ~�_K<��� �f���=���35!z���>�%�Ҿc��p���IOg#�=x��R@ R�^��5�9���\Z�l�`J�j:��� ��I.��D���qk�표w���23 ��i�{����!I�Z-E%e��X���T�"�,+B�'��Z��`},���_1:��*�;$������5�x*��J*_g'p�8=�����M�b4Q��-ӧ�&\��x�ߏ��nmcM�f�#�b�	C�̌�>cFIv�Ř��ќD�픙��9�}l CR���,fgg��-Ҡ$��Ѩ�?Fq]#u�Z�,.���T�u$�?�_��<�WPH[��G�*D(u%Ϝ��.�JCq^q��Y�k/�@AQ!�X��O���a�Ϭo^ˬm^�t�4�����}~rDu�Һ�{c�����Nzr�����8!��L%'3]��n�BX���zQ^~>e�e$��ݠ�@&Ȳj���?0>1DB�����{_��@Q�4��rG��~�AC}u9W/��>3+�5"=�5%��
xMZ��6�[Q�'��2d��M�xsX�����_�0�Ȫ�X(W�����V"^�۵���v��Wǿ�4��㪺��ԯ&�� �J�$�$���S�W�(�.��װq�K4�~�1GXn�0٢��÷��M��J6�����uT�
����ǽ�<!��j8���>z��{�J��ǿ�'~�q5�[�R�~;��
��v���*a���>�V2�����2"Ms;���a����g�>�k���d[����k����h6I����o`�-!�b_��I�-<�9�RH1��֋I���=�����%��W��?P�~m[��h1�W'�϶p��q:��%ͤ��a�F�����K�Ɯg�(�^�_=IMa-M�d�g����ё!*J�X^Z��q�(��ev�íGOXp�QݴF���/��A<���EB���oH�/��0a��)̠(;����dNԣ�gf���SR]ΊB����{���y���}�(i��xG9���x�Y�$�ް�}�_&���c�?{������n
r�Y���ϕx����������_�ǽ�a�*���)�Exc1�;N�*8�����#���W׶��{_e��b�K+�\_I�ZVKժf\f���y�����c�r�K����Ǜw21�f���(���D�K�}��P7*���uml�{�pLɽ[7�M7QW��oi��j�Vk�J�^�xUb	��L��,{#L-��_����������ç�C��2f����S������D=4��{(o�i�zfg�%�J|�,�@��Vq�v;c�N�jٺ�����0f�I��;�]F��c�F�B��c�gV������n����'뫊���[������D�?|u�?�b��B)VIRX<�\�1��X<N8!�,�QR�˩_�*Gd�@������*��|.O�gjb�F(X#���Դ���|�����!M��⦑��ؓ���2٭�+��w�ǔY S�ꨂ��L�����ׁmvJ��D�B���/X��Cx��.�J�!P����c|.;!����;ٱ� 1� �:�
�J�ky�H8��������	x��!	o�N�B�sD�%�hU0�i%ʵs��~t���FP싷z�`"UR*�
z�K8%I+��c�L��X���qm���F��b&%'���RJ�j�37U��3U����\;y\�xM%z�U�i�Dc14J��� �si��� l�I��N���"<�$+�H���>�?� ,S	i��FB|��?ɟ�H��m�������Q��r���X��e����a�SV�^|� Yy�8!ٛ5��]PƌMt����4̪�\��}�&�b�,�@ �� 			Єd�c�N��Ǝ�N�o?}�t��77�?ם���v�xvlk� ��$H!�y�*��ԙ��w�oo(+���y���ꜽ��}�����n���:�"��s�����訴���0߸kn�gL;		�y�z4�hV�ĭ컀��0
��:;1Z�i3���&M��k�,ƴ�31�:o�A߹���O���,";��+n�d�Q/�L��V�)E�J�� ��o�������Uޑ\S:�b{	3f�ü��5i
FZ�n41��Gc<���۱��A��0w��W�;U?e���mE��?%�ʬ��
Z�1��õz&�Ĕ�0a�T��l׉!��z������c�ӛ��G9K���w���1u�z�6mx6u�-L(���0�|u��F��W��_��/b��Ś���K[���� ���\�T�Z����Q���Sx��? �M p�5i��/���@�\D�q��8��>�?��(�c�R�����,�O��m�t�]�Q�h�Qo)��C[��[[^F{�xMf|���������b9���>®׷���qt�W�^�k`�5\|�s���H��9�|�$�_~3��MDY��H��r���{�᭝/�T�j9e�g���*\���o�����^T/Ǭqi,�5E�`��o��ٳ�ݍFmgϞG�ՂZ���#'�bʜ����f�ȦR���f~k*�'t�M�Ƣe7��m\8s
�N~�K}瑣�@������.��?q�<>>~�OS�&��+Wc�M7!��}������w�a�����{Qo���:���oc޴n\�p>ҩHj��A|���X0>�����g���/�|�,��{B��*d�M�S!��71t�����&!�kWߧs-T�)������}h+�a�*x�g�>�\���ƒ�׋DCr��o����Sfc��c������ǹc��GV�Y�>��z���㽷��53'�ԫ���#��l+5�>�#�B�,~x#Hc�M�b��K��Y��[��?}m%d;'`��_�C?q�c�}�>�Ok����8u�#塌/K,��w��W#��a��]�����8��P7	�l؄��3Pm�����dZ8��UiOp\k��[��d�
5e��7�L]y����|�o�����N��������$~؂�Ja���k�b	|�Ȇ�Z(wM�+נJ���;���/&���Ud�l+P�D��R����Q��$���ɶ���ƭ�|�����/����X}��6�j���]��9��MC�8��ӞX`6�ZPn���Z����8�2-�    IDAT)aK�1�k���'d��Si,[���-�gE,�҆|��j����3��FrN;��9U�#��J!d�K+���m�3p�5�z�Y|�M��i��k���~-g�&��r�3�(�%��RI���"1�ϟ?��7C�vW'�m(2ke��,�<�R)Lnk��׶�������v��?�J�ƣ�b�Z��,��-��fs ��*�� ���{��9g��͙B6���t�-���<��Ґ����r��y�����g�3HFr�O��&}��G����j��:S5j�D��q�H������~�o"�N�����]������p\�D�)�.M6�c#�8j:��8��Ã�oJ%��i�f͙��Ӧ��K��l����>��٬��v��+�b��w��u�|� &���l:�|N�jk�`xh �ϊx��T���-6~�҉R�ã�<8�A�o!�wv��}O>�.���6���!�=I���JE����/�������I l"e�SQ1��Ub��D*�B���l?�Ҋ���f8ih)����羊��V��n��HC[>���gD��Zؙ��b�uK�`�LJ(��?�қV��7c��T�%�A%mɡ���/1z�l���Y����$\}M�b�g��,�N����ža���I�J�q�8�_��ӧap���WC��1��ǫ?�	N�H�3垉X��G��3.3�(��C���B�?�6.�>��1�\�ُ�a��	�4m��Y��߈��!��&"V�Հ4�Yrp��-����(s�l�'SF�k�����K�a`��|���!'ӕ�*�Z9'�C����3�U�q�*�64<��q���)3p�c���)������
�ڎ�vv.���џi
۵f͘��ǰ��g1p�3�L�|�p��Q�I�@�M��1}��X�lJ�{�{_������Å�Ø{��X�����������w�7k��T�
��Â��g�{xyۛ�
]
*�`�6
����P������S�	E�
V�~/�X?��z#�8t�38��G8��ADn� ]�a��|�$?���p��E����,wŪ�1q�,Ԫ�������S��-�,nX� F��3�9��>:��Ձ�mI�w��kQ��DJ�{�}��u�V��C5�^z=��p�����4>��P�L�4q*����*�z�N�w ١3�7��,���s��ѣG5A��g�C�P¡���Fh�����K�X}�øv�DN^��<��=��5M�tВHe��ه.ݘ�-�I� *���7Ο��ݵ�����_��������_�p�:)�i:?�����B3!:�f�z҄�s�58�͕F`eD��(�J��#���!�����>��p>�}V�A�������>�N�%[�R�E۸	���9��k���o�8�&|�!��mGze���щt,鬈P#������@Xw�u�"3��ŃҠS�����B>��ᣔ/�w�x��iO!��i4�#W�I+��>��|�T���_ߎ��C�Q`1o�b���a4�.4BR�1���f*����>iY3ۤ�n�>j-W�:ۘ8_���`-+�ő����ۑ�ea�KXw���완�zM=ؔK$̙ͱ��"*dryE��炵~�h�C�҉����<��4N��oyY�H��E��d�jp�5g\۩R�i��آ��]M�jUGQ��qqd�b#uT:��� ��	��ĭQe��<���~ �Y\{�J�\s\����}!7��� u��)�"L�V���v�2[��	_�v�ZM�d�2� ]�rh����-��b��Xv�\5���pN&�ёa��D�뿤@���]�g���=�����z
�̀*�s`+`Ǝp��||h?�S)��,ݺy�B�P.��{�{�4*4�l����i�:�Hu#���QǸ22����J�#���/�tXG�	Y��">�{�r�b��4l�Ot)�R_/�錂PN+�Lo}dmm2T�r"'�cg����D��G��9����}��>o�8c6����a�糭��Qd�@�]�������6uN��Q��]=��~ʑ���,G��N���'?±];��n<��_�D*�5S�S!�m�m]���sg�N����!�O�,��3��P����h�LJ��Ԭ�Ж��on��/>�vp�u�x�x�{>��@aFZ�Z�`�ʘ�ꐐ!���n��
rt����?����+V�٫k�$�:{�f����7��W�C�BTX}׃�2g!�lQkӕ����3ػ{N� ��@[��z��}W��0�?���YX}�]�9wj~ Ȗ�x��Y<��DTF���U���Oa��QC=���؋-/=��'>F�&�'@w[�.�i"�����яO�‬�	8�; '�E&g�%�bG���}��QcI��u�c��0�R�>D!r�%��c�>��}o�j2X���YRY��XC���C�0i�UX|�rtO�JR�>"t�<�O����FT����h(Tʈ�:�߽�����\Y�(q��y�J�<�>>����8s�f.�+ׯCy�4}�R>��<���"
���p�����W�m4UB���� �ڴ�n�A����;b�O�;�{�T\��ϼ�:\w�t�LV��O�1ZBƩ�=:�Q
�p=��s�Hɼ�=rR�I����EO1��_����v�F����3s�������8֡ӨD~Yz��}��Œ2֬�����2�*Ԛ
�64�H��C.���ՁZ�*�s�{�A�C��Q�h��P~^+@&��F�1"L�N��f1���L�A�d�ȳK�Nxh�M��0��\͡�"el��c��j��B)�l�N�:P%��[sZh��>�t`��z5^K^3���y�>
� V�ɈUZD2��q\���v�؊#GH��Ѫ���ᎻD�*"p�������[P�a|��8j��L�$�d��0%�<�v�IYȄ>�fSƞ-hd�r�E._F����X�hU�Ii���e���{�L�vr��&�%�-��_Խq�y�~��u:��$�!�1��� -��o�hԆ����X�!�Zf����sp2i�|�v�J�Za�V���� ��knŲe+0a�U�7}�>�/H�5U�2�D�24�5e�$-j��P�r�~b��"��c�U�zH�{1m���:�6<fm�eM|��Hf��1\F��F�YA�����T�BGf�������ή�/�7"�&r�2��"�P���֬��H�2B�8����V����FƦC�~�k�[�01����*Ξ8�W�~B�\6��<;�G�ρ�4��A�2�,.\�G�R����
Zd^�'Ć}�t��.T���d4&������^|j3�C�<W��VI�^F���=a3h��Ô�xA ���gIs��u���4ڵ��;8��-�F�4<��g�l9�t�%��pxȦm��������r�B/&͚�̩E[�� p�(8>N��/?�3�8Rw��l���3��/�.�NF�[�4�Ď��i����'�S1��N6W@Ǹ.uutO�$9S��Y�s��D�ٶ���h��E!n��1c���e�t�J����ܩ�������^,���>c�հ��<w��3��Z�'�����sgTJ��j��4#/ڐ��B�(�~N�	�Q=TJ%H:i�\}��s��Ց�FL�laN�`Hq�P�9��2V޹	����j�t�I���uT
E��ӧq��I��=�̑���#�'g�Ϲv!�͚�B��UD�rG'l�}'>�X�rVl|�>Pm�1������'�^IfϺj֬Y��gN����8~��̾7��=WMA��󃣘�=����3���&V��26��@i�4�2��Ն��q��m�����_�S��ػw/�y�9�<sV�	�5�.j���Ѵ5v'�<ˑ�\�\��{�¯�����}�]� 4�2OY��d�it��)g߾i�������з;;�~�����cc+L�R��i����!!cӶ6����֒1�����R�7�fT�y�y�hdC/T� ��4�c��������"'e�P���ﳡ��E�"�>k�
����6c�j"r��3�%+Вv���6[r<|��f~3FzJN�	���dZ$��-�����\:#�v��1V-6J��yJ�р�QV*ka�:H�QB�.3�R/oy��51Z�b��Ÿ��O:Y�$Z�`���Ѭ�����u밙�"4jJ~������������DB��x���)�vZ6Q�PA�~u�M�9)z��F�(��Hy�+�1K�С���E�\�lAAS&Hi 
>����*`d9z���CG����뻒|�h�J!4�^C(5뽖Q���w�I�����P(TtH�4�h�8~�
ۅ�YA���Ȩ�Ữ4���B�	1r�Bk��<<<1h a&�B�����(��2�]�v){$�wΜYH�|i*0�d�ƣ�l�2��'X��
eS#�ύ٠���B��	^e��}�u���~%�]h
K1�#�N�G�Y����0�~ �aq�[&�R��w��́ˎ��)��/���^���*C�*�4���=�<XJqp0�j��J%2�����,eW���9�Y�dOxr-���,����"/�� �e#��˔�����\KC��\����b�F�VY� NBT�HӜ�^�r�3Zk�#d�3��I\bF����!p�9!�4��+����9�O�ˏ��<�:etM��~Q��Ȗ
BEx�I���Z�c2� Ҝ5/����U*�/^7	��:=�w��o��Ӡ��]_�#�̘��&d�{#5%l&A�4n��u�9��|�H+�"*Y�"������3��!`��7o��@�Y�^���ti�|NH��pkJ=�lR��0�WhgPkE�p�=��EZ�_G�kh8����P.���X��~L�v5Z�,��<C�-������)��QP�_�N��Ӊ���H)PK�ղ`�s
�r��m?�>N����������Rü/��Z#�,g4�B�Ν>��gOi�iڻ'b�܅�8a.�(ww��e��m[��3O	��tOƊ�?�r�x>��R!:�i\꿀�K��=k.�q���5tL����˚nZu-Y��5��+#Ŗ4�6�G6����_D0ҫR����=�L�����T�>@W����쾛�O��m\��7f�[�����=�������T=��k��-����ޘm0��}+Z~��ޕ�6mZ�Xnӆ�a���#�Q-��8��=�а�?o�C�]�ƭj(���!��M�j��p2�J��+(�	k�Id"��7dOn����0C#c�"�1X$�^�X�s�y��:�7l(c��!��J8/Gr�(���2 �,�thÊX�M��+<��t��es�"v�ى�;^��j51{�<<��g�F��x�ti�-8�Y/k��.�!i�>�Ç�a#\Ӛ�*3�<���p���ؚ!g�ё����&3;*�,8>̴���9�1�Z�>�QX�Т�t�ju#JS'��d@���C��
i�-n^޼c��(�FH��1�jZ2~�ff�t�.���DZ\��@�N#�,����Ͽ����`p����q�t�8hj�\9�Qf�Hg��R2� $+���^K�ά�P(�'Y�j_���3�u�**QD)���R�ÈF�Yg�^@�c�(�J��Eԩ����զ6
Nn}TF�HI*� J���Y���Xl)�BG|��2���b@�`�Z-�V����s���q��;*x�������bɦ;��|�˰�.�AZ�JGhxM!(�J=F��L��7��)�ɛ����!i��pM���2�	f5�i4\N���jC�����%�,�4�u��ATܚ��@�y��R�):[]!P�l8�,��0�[2M��u�a
�zK�$t4J&�,����/����G�!���p��,qx��R���#��ғ�@&�=�Po�0n�l���s�K]h��ϒ�)�U�
�6������mlD��1�s��	�Z-�Y����A�j`�:�l�4ؕ ]TwE%W t�`��0
]��\���$9M�Lz�f*{��@%4�O�}���Is�`���:��c��8�@�(Z�(�S����!�/W��}�A�bȦ�~i����	�tV��X��A�X����6��W�4P�/��'�ٺ?�Т�nN�IU�^WٗsM���	O-����Yt�j�����4ʕ6�ý��P�ܶ"TJE�wD�hC�-�.U�����s�0R�!�1=�������~Ee�ոa�"4�r��?�����)�jT�l6p��yi?��9ƻ[��\����%ڈIYȀ���Y��R9��מ�C�N���z�ٖ��9k,�Җu�ѸRz���3��[�������O��K�}�T�@�ܬ��E���k��s&F�y;;������`�̫��9c����B�Ԫ:�Ɋ����s��!F$c1�d�
���@Dk��N3��I9$�e�l���P0�1�C:;����v3Yr�����][�(�;#w�&!�G+���Y��4Ƅb2��)��cVC�DGaA�� �//�a�0Є9+L#f`E-˺2Gβ����� �h �<�$���P�FG�>��`@D�?���Orבھt*2�^�����3��"��[4fd���BBo��7����ҽ�K��10q�,<PDhv*z¬-��(���p�^��\�A�w5����u�^N�� ���frR��R��1A^�~iHd ^'�
;���&���f�S�ry�ۏ���O��3f��5kq�Ï�s0i��E���D^�Z�#�/c�@���b^�d6^�)�F}>#�2f�i���f3D�ߧF3[p�:��D��(SL��7��Ty�R����"���(�'jeq���r�!��T�����|&�
^5�:���&�A@�9�.݆��h �b	��U:
V�a\8�?�s؜:֐.e8Y<�� �L�e�صЂ�3C"Zn���:�t^��x�z
�,��}_�.��Y����r��ܺ�1C4Z�L^@����(�PȧE$e�@h����&�ȤLi�F��k��Ut<�=��2%4��g�f��;�)�A�,�}��"Z9�4� ^]��\S:u�4is39������yL,l�u-����O����U�'�5k�������b�� �����T^��zr���J	�}�'%kT\�.�w4��r�
��ut�;u�1��������%:*�σ�m̒�[c��5Q�]�1yg	��5U�p�u���Z�,x�	��3Z��I[�{"gr<��|e�$pr@:���.���wq��h'����!�Z��F��F� �6�F���D!S�Ic���i��0��B�΢>���t���4��2R�|�}���zhԫ�� ,�7-�BWG��E����<h�`|W'�v�CR$����������Xi�ܥ��2�GA��{b�,Q��F�|A�Ą� ��O��Ј�/��i2$ێ�L�_�j�ٶ��z9ǵ0�s",!�f��A����6z�S����������on[;zt��~��7.��m�ȱ�V���W縺�;�w�#_ر|ō[��L�0qܤ��r�?04�u���#��n��Mv6�Æz^0��qf˔D"ec$RQ��F)������`T���]���	1�{�[|EYH�T�u�pQ�X��Úߛ���|39S��(�C(��z�HCC�)q�c�9 tFn����ZL�����.�R6�0�
z��-���
ZR�X�m���_>�={�T-ī�ش�^\wU��6�,�5�(j��`ZB��nK}�^�7�� ��b�F��aV`��V��/��D'K¥KH���D��vd�ȌW�&K�[�4�3B��	��IK�Wg3�����ėUVɺ)�7���An2���p#_��t����.n숅z;��x$�#�F'?\��?��Kh�����^�>��G�kʑ�a9��fB^R4��4U~�����9q�(x!��C.�E�YQ['k5�s�3]DAS� ���ѐs6qVh�L���dnK��ʐ� pi�j��3����3t֡�2Wv�|='�0|
"gY�X    IDAT,O�ɝc��7e*1��-Rw�,���=3Y֦G���G�A5��rG�l�<���8�����?��Y���
�n`�5�x.hy��8T.�z.q�"P-���"��ҵp_x>�,�2�S�9�>s^;k�%X۫K4�+�ȒM*�G#E�@
m���-�M�W?l����FD�iة,l�� jG��'�E2�� �N
�2U�Åz�I��m����V[b�N�Qk��Tp�셸��Mh�ܧ�!����k�YN�#���X�x���&:�B	�zݠ���H�@{9��'�A�o�����,��~e�m�$,S�g�/�e�H�P�9w|��ly�|�n����	aI����<�fz�I`�s��Gt�)rYTG�����n��	Q,WԮ�Nr�
�+X�ƍ~���2t�X��S�������+0u�0E�SJ�_�9�D����v~?����t���f��T,W
���(�TQ�u�\,rpRhUt�����2˪�g�^wqi�g�Mϯ�h�4�����2�c��V�y��6�1a @俆�F��ua���&d�Q,bx��g��2��k<�����C�z���{��B1ˮ��ۍR�cX�ArT՜|'�K����]��^9o����[��F�����������e���Y�ʩ�mG��h��뿵��[�.�r�3X�(ʾ���~���|
���0��ך<plac(z2�g��h��
���2
"��`m�J�VY7��^���}�0�j�)e�R�1�f�Gj?��0e���6S�b�ô<d�k�G��ś�䟸�L}CH!�,�3p���Y��I��D__
�6p2����OLX>�z����/~�QZ~6�������h��Ẹ��	� �L����f�;3G<:+!$:R��N�BN��.4���1�sHjk�g�A���cX��#t��Ӏp���~R9���h�2~�@+����9�d����@T�'���x��ױ��*�tv2Si�w�K�0a�A/��P.�c��7ABD~@C�]��k����|Aм���!���1��=��d�)W�p!,>�x�0P\O�b�p�1���{e��Qk����ڛܷ�Ĉ�ߓ�Œ���c��Ek�r�1lEUjI��B�!�uX�5��0/�B_�����z��,�X.#���{����Ъ�����Ð5��{-nZf��dˑ�����qO�煾�cPq^$��=�<�Ð���	�Uf�J��H���#�;L홐�yS�J>ߴP�ܓ�d@ɚKg��&?����4��7��?$�i}��,1?��^���oV�4ti@��y��/�#�yT��d[���VY��!��l���̮HZ��zP�Jg��0GM�	;Mt��ܙ]��A>�Y�=-��PuH�K'E�g�"M�>���Xw�T`�P(Ă���h���3�w�><�!׏�����ۜ�˶�%�x��x�k*m%��]l����0�f�b����_C�4);/�B�����bN�l�Tά�Μ9#��؆�u��7 �:����/`6+R5�7�K�5Z>'�RIMA>	��AzM���F�'g����:�VӖ�\2Q��s���y���Ʋ�L��=��P%"#1[6�	5r*���)g��dE?q�ܵC��*)KƧrN�Ør��MԨ=��&u��~�������F��¾}K���o�7�,�TO-�v迾�yu�M�w-l�:��7H�E���旯;_Z�J�Z�n�aupcn�-o�ƒNw��9�z����	�Ԯe�M��@{	��l,a؃�CKz�y�r,&�נ�J��Η���h�)��Z��˛�$Cj�{~�IN��{�Mg�>n�sk�)��:���r��QF�<��d�9�9�h�=�K�ɗ����$rk6�B�]M>C�9�cge�7�}�ӧ��T�>v��L%/S�YG�A�x�s��in3� h�cڜ�"G������;j�c��٩�A]x��xx�
T��6J���ƭ��r�y�Q�d\�8 H�3�Ԛ�Y���ǎ;02lڛ��w�uf͘���Ƈ�����ԶB8"%d��P����M�J�92�cP�^l��5F��6���O� ���!����Q�!Ο��CG�k�4U�c���؞)������:d�h OZ�9�dؒ�G�l�w�MYA���8��{��������S�9��$s޽a#��Y �_dUǆ�
�FF�}�Q�p_����'�]N�g��o�l�16�o�k03����Y��>���H�D!�:��&���g�l(H��g`J%ɟ�Y����d\���[�9G����������5;u�~���y2�����H(�[ך�MU�HϘ��!��$�ҩS�I��7���<f{�a �mV�1*��˵����1�����@��D��~&��ٵ�]�I����:r��j�"&9�V��4����&�J�ۋ�g�g����y�Q�3{��󵗱uۋ(W��_�p	��aX( ���0q���� ����W�=�O�ЍϠ�M�+	�\9�)��u]|r⤂Ζ�Z�;p��$`Qp��D��6O!W4���/hkdI>v��$��,���,�_�q�<6B6Ͻe㵲t��n[�]3%��m|�ё&'"�"�Q�GX�,��\*I��g:��;���{�_���u�C��+o�|��7�����pr�
{W.��_���/lk���|�S�������oz���_kx��Z�%�Z�8r��EV���K�1m�n�ԙ��8�X���q������HpcFkx��:tnf�rאR���ѩ�[d�S��u}2ԯ8t^�7G�(����G�q����J�7�7k%�9~Fr��ߎ�.eo4��!nX�L";�a�R�����h��l�����꒣�c�Z����0���3z���8;�������0�mk�Ra� ����>[��8iv+�8�����u1���t�q�E)`�p���;h��$�uc(A���Hlj�69r�|����֐��)?;��Ƞ�K`;l�@mdX΁�H�NH�����6e��S�1'�@C��;��ΟF�Ւ��1CWT�{�y0��CT�eܝA��=JG���2�4��,� �,���Ҡ���j�1�h6Z��1!�8���N�G�>VĔ)SP�p��k0窹���U��H���$?�h
�?���	z��N�>�Y����q�"}��B��y֞[h/�+�3E��pXҊ�+�ob�$%�'i+�=���x����\3�g����A�HF4�6FY�Ʊcǰy�f���v,��;��ҥK�f��̓,XJ�>Y�7�	�r:}�4icD>3A�ʁ�C�5p�g��'��,9C��Và�Bø�`��8���i�(��;�>�W�3Ƹr�&a��"G�{S�{c#��e�L� ȼg�e6�ַUZqO=�8>��}T*E��u������؛Z���-{Ӕ
�������֯��7�ĸ$j����ɡb0��a���lDԖݜ[��p�Y;����4$Hh"�b@�gA���Yz#��u�,i����\��&�x�s��$��ÔTx�u�R)���|QD�ju��Y9x����j��������T�����&�e+
`�M�ʥ����%���ɟ�}ǡ+����I����nٵ�o='�@�{t�K����]�n�����?�Fc��u灅�����zc�P�U�fV�-8"^`F_!U�:q����Þ���Y͇ǚ*.��D_f[�HQ\���Q��_e�+d����k�_|�y�@E�	�}�j��B���A&�3�"�I	Ɂ5�]b4蘮�17�p>�w�yG��$��e�V%&/��:Q���Al��m2B�rT$�b�C�VS
�c�ڵ��_۹SF��P&P��&�k�΀`�+FQ�vqФ��a�
ATĐ��N偏��\�i��$za�=�1�A����q�1c���p8.�r�Eb�3&F�4��l^���vٲe"�����R��$��IƦ̊�}�����{�Kk��y��i�lf6�C��M���A�!�'�o�ˁ�؟c����/;W�R���K�O*;t�/y?�9C�!�A�n�`֬p1;�s����!D�ρ�CV$Q��Ae ���Sf�Rj���seL��{M#,�6���x-l�b���2�7�<�y����I_V�_6�sl�z.:�Ke\��!��:$��
��z�wR&��Ñ�B}~���혀;qҚ�(�)��a	5�:C�{� ���!����w�U��u��Ӿ�wy���:�|ou�С��Tj��+���:�,	��K.�!�@��KOL2dpN�$���<6�%���� 3n�7qw�L�%���`�|�'�{Rrк��K�݌�,��\��"=��0"^��%ɓܻ������я~��Lm�%�]��>L�4�5C#�̀�����?rS�ަE޽b�.G�W�J���A�q�q@q��� E7(N��h��,$dXS�	�ǒ�}d83v����]d�Y���:�}���NA*�Mָ��.w!�alm$N�;9`�B�B1:�©E���d�u���94h]����;r��}n�úu��u���lX�P!/��>�dDwb9�{ŢY_���{�����п���wn߽�oj�?���ΌU�~����z�u�X8{�G��������ۿ��o��cg�����A:��]g���^��+n��S'���W�+ʍ���Z�J�<�P�p$g��yP����+�[o���s/<���gd�@��j�j���Cg'���X���𵹭�O���֮Łw�Q�2{�%p��.Ae2d��`�@��Yo�C�a"47��r�FOal�x�n�u�Ѷm�����}��7w��Y�:]I�~�ؒk��2-d���yD���-[�j�2d��+��<ˤ���Z}h�9�a��L,�R1̘2w�y'�}�!��xU��%=c}��5a�u��Տ�R �d�Re�ZX����&�!��Q�
��ZdF����+Ūs�n�S&�t�}�q�>�dbg>֩�g����=��$b�����˦E�mf"+��[�NA�������
w����z����1��X����B9B8�A� �d��N��ٳ-0	�������5�	�(7߃��r�ls�x�r�^8tPY�H��
���j�ç��2���2��_�b��^�&k�1�j���	x}b�sK�	Kq�}�Bۑ��=ɢ<'I�MG� K��1gG�3�}&���K�3� ��}p��x�d�S�O�swb-frD��6m�l��)�N�X,+�R�0����y�wX� %��АYsTT����q�鰑�qp����"r:Tլ+[�>�,c� �Ac�m���.��6(��ˏ����������O�P�Ω��u�l<���$�uN�0�]�l&/m����^I�c�B�Vq��2�3�cK���3���*=�b�O��# eB%�!�̙��:yo���C�I�QMgP����Ʀ�g $�ƾ�FK��+�c�����S�� ���i�4�i��$zR���ԱR�Y�.��}��{6~}֬���e"�7��y�]˶����rפ�#A��$2�	x�P�z�+�7�.]��/�r��O���G�����{卽S��[��B�oݲk���׬��I��������FQd������;����([��R{K�Fv�z�	0���W���'����f�89�d�	4�L�N�7��*R��d񬍭�i��}�Dj`�$��f��:1(�%�[�xw��{�4�U����s�)s|�����;��>+7{B>�fqضEp&%�nnrgc���2s\n�8f;����6l��Nm�g�#U�JIE������7�Y�A'56���o-�!=��#r���/]�$N�K$#��qF�sBL� ZWr��Y��� M7|j�>�m;^5jSq	&y&ӓ��Aa�z�]�'�l8n�8�9s���6'�<=�8*��G����b�?���UY���#�����Of��Φ����lb���Y�y��֋F�g�5�g1Ǡ�V���$;3�(��s��``��ɧ��A�Lb߬�30���kx��;���{�~-� u�{sO3&R�#��ϘL��� c����@��Μf5Xh/Wp��M8w����2Ae�Dqh�[�M&�!'b�Cמ���K9T�E(��Չ����y�g$QJT������$�q���3O���8��]�`�,Y�ݻw+2�:/�l\�Y|õ1��q�ϯ���ղEG���Bc��-�9�?��ҥ sxpo��W�Yc�I4e���,��VO2k��C��k�Dc�!DkE����z]ˁ���s��fn$��%�z��]2���H��0i�DL�6MhY/��9��!ʚ =	Դ�,�>2I���f�;sV2�n���,��O	�tR����3�Mť��8{�<r����ffg[n>W����J}~z�P�WDnMl����[�|��::T>$�Ab2-!e�}>c;�,=�f`j8O�\"D-�ːa;qZ	�h�.d��6h�rL4G�k�%�D��mZ��rN�5�q�k�������=+W��5�+� ���s���;�,}u����R�_]��JT"��B�j5gt�_�g���i���h_v��ym��Ͽ����Z�����ԭ�����]����Ee����������W��.���/7�ft)X#��ZufL��U7�$�N��*�Y+T}E}xW2��W����&�7��H4
�I�q�]w+�~�3��V02IAbA��2�kLE0�Ɠ@$��lŲ�qݵ����Cؽo�T�Q��z)��@}{���H�s��םZ�f#�	P�h�����*��zCm1��{��7?nZN�ܜ52���cG�Dډ!LH���Zj���:]���x��gUwN^�cG�Z\��� 9m������c���I�����qj��胣xu�����8�-/
�6���L�Fmΰ�y����U�
�6Ϥ��t/3��|�ITGɟ ��F���Ds>�'��ϻ��B.bL�Fg�(aч~X��Ϳ�~�F�N�N��S��/�	��a�;��j|@$'�8��/Ǎ7.��8t�}����Ψ\���R���s+'�jz��)�Ct�c����r	�?ŃjOˡ\,⡇�0�W_}ϕ�Qf��fc�]��ӆ�ab>�]�L(�:���勒ŭ�c�*�<�ܳ�FZ<ۼcN�"�cr����5˸�N\lxr&�o�J{.ĭ�ުkg�ِ͠�t9�O�o��|,��{TE�#U$Q#x�}��ԫ��3s6�_���x晧�%aF��kE֓ӎ���+C�D����^>;�O=����Jd��Q%%�V�`�H�*@�Г3w��:���˗.�«���ȡ��r'���A2/�~�w�� S��H��M��6h�~�������&������ٳؾc�h��cʱIr����= ݇8N)�8W�� �Y���ŋ�y�޻GϜ��;g��6��{��;Y���hZ��šI�!h<�$����ٍ������8}�e!���5${IC���Qq�9�o�����:���R�xp����\2��o�~x��[�=q����l��A)�Tơ$z��i��Э����9��|��/;���ު�/o�f��`f{���_��V����	քڿ͝���������=���I�WY�9�_��9WM�M7.�C߹s��fi�b�/���y�M@����f�!�#]{�-�;{�� o��¸qg�pr�h�����X/[hG��j��/��+��o�=���ʺ)�"Con��x-dM2� ��xj��P[)2��x��+����=���$����OK|%��d�t������'��>#6�t
4X��|�AL완-[��໇t�c�(��|8��cF��ڴАT(�ϖ:���G1u�lڴ	�[�m��ߧ�z�i������q2TG��K�1�D��z�^����Q$��R��Zv��n�ݟy�aa"%�09W`���r��k��c�"7n�c�%��(�$�*)1�#x���Γ�߬�i+��Nµ�e�X��ܹ�Nl۾o�~�BNuVQ�    IDATY�,��H8����[���8AW�!�x&2��`	��>{����|2�g?��8}�4�}�ye����L��M�(��9$�W����ƙ�Z,{1��u��($�hb\���w�Cڲ�����Jy-�����1ҩ(������t�l�&�J&; ��E�aժUx����uL}U{>����T�O��[��&�D�������0R��{�fL�����ϞS \f��k���k�`f�	Z�pP����5�g|�����c���:?/����3t���A�7ᮓLɶVM{I/.&T)����8�oa��X~�2���.���!K%��ɺ�K�9�+��_L��$Dm��</B>GUJӦ�6E�'�B�«71�����������hP���58��$�]܎'�o|IBe�Ҕ����^^Q�5kVi��<����j�ZC��Ô�T�������.+ ٬���i`��pٽ�Z�O��Uk�(X|���:�l�%�/I!�J#��n�� <5o�����g�.����vwW}Fc����o}=�m�ͯl�������|�DQ��92�d�Կ}`�__7e�����������/��s�B����*�fv���;n�����އ���s����GO?��������&ե�׆��D�pFUk�ӱf��x����ē�p��h>�R�8�M�ńX6ց	�Rk�i��eD}�M+��ٳ{���{���0�5���M��;gi�(�����Y�ˮ]��׬Ʈ7���ݻ��ƨ��m8Jњ�)pk�%�N�|�Lc����137Bv��c�w�	�/�;���߉�Y�:$�7iˋ%hǔg���ԕ˘u1�Y{˭r;v��#G��]����:��Or�bB d-�mw��	��144(G�C�����s��M�bߞ�xy�v�fp��`C|�0p�$obr���v�%,iIb�����A)��C>�kx���{�
Ų������B"��=%���]&/�Y��a����ʯ7�|3�/���^|��J{��3*!%�s&0ֱ'�l|N�K�����2���t�M��[�ҖW���}�hvl��5э��U�}|�4n�����+��2�8{�SF8���u+Cg�������dVHQ&^;��j�̔������a���Y5U���t�AE�<��Ğ{�8�ۏt!'�������|ǌ�o�Ω��4kt7M�e��o7ވ_~o���!w	�K���a1�7��L�bzk�+q�Y�����A�(�LŊ4�󶵷`t����zJ�?�!M�8��Y#��Hދ�2��	s^g^�ҶIR0��g���V>��3zo�t����6�1����қ��xfK�<uL�32�Lܸ|�?r�{W	�\O�or.�=�7	4Na.�"�����O-�`R�C�XF����C�?������6S{$$�ݴ���A�yb���/'Z�{���,G�ȧ���R 5<<��l��t���(
e��zB~��/��(%,�<��q�#�'pJ�d㖧�'�9s�L�v�:���~(�D���$�B-X^ȧ�jت���U��/���/�[|(�бc=O>��o�:�?���S[꧷�.�1����/<�өC���r��������'�>���)���7T_8mܓ�-�����W���vqo�n�_~�1�4ҙb�5������R]c�.�1k�4�]{��.���Gu��>f����FS5#����k�ӑ�F��v|�WذH���NN�!��ܲS�NǞ}��o�ۨ�u�����R��,G5��KB��&ɈF�sт�q�u�a�޷����p	��lA�̾���~��1�\�ț���RI�����*���a��Ix��Oapp[^zAb-�\[M�
y%�JO�j�W �*ք*а��gF&��4�D4Ȧ��f����C2�<�|o�m�ӟ23]F�$U�}(�P��=&?2��_�M�߫��7v���|q�4���V~bxQ���&H �>ד�a��C[��/~�w0:2����~
Nc)�V�3vTW�8Í[̒�@,�����y�ϳY�_w����o��W_ۡ���	=�O�������ʐ�hH����a�D;��wm�����ʔ95LN!�:gR&�aj�I�4�z��J>l IK�JT���h��{<�������O=e�Ŝ�Ƒ�:��������!=c�+��ɢ�Re��DK��p��;q�5����sx��7q���<q��D�Mz���MA�,Ŋ��hYE.�[*��>nX�L����wȡ����d$�doQX�r�G�ߔT��8��#Y2#�@���/�;��6a��3}��S��ꅑ	��u�RѾҠ(�&h�X�1���D��^�)&#o��ƍ�V}���>�+A}$���e4#x��|\O]7b�G��%K�캥x}�x��!Sv����2��(fQƒ���M�V1�"K��xerꔩ-�;#tq������?���xy�V�FFaQ$�L#�Xm-V*T>~@17N?����X٩��Zps�93����/�Ѻ��F"y;�W�D͜S>�K=���i$�Q���,G�̙36l��{��Dr�ދ�0B._P�)�s9�:l��Cw��z���&�k���+m޲c�k�~�W{N��58�����?�v�s��_޺��:������KM�+-�ّ���1���-���%�n�0�v?E��~�G�v8��R�*g�K���l`V��� s��k��^O7ke��.*U_��ɮe����D���Y�;3�1�
�"D��Ą�ݨ1k��p����T)⥗_��#�"��eV6�xW�J8�4|���bV\�W͘%b�Q�᳇�F���^�[�ˉs,(�Ȍt	�2n�S9 ~�X�L���3V��*�-���فO?��ǎ�&)��\C##*)||�88,�p#3jBٺ�DIo�W�V�~�6��3�h����&ty��傕6?�>:v�&W5�C�CgLCD��(��p�����L��6J]�\L�:�������W�K�U�������\_�����g@2�şU(���"~�w�����޵���(������WM��I��2�!Al�4ӥ��.׉Ϟ{k���[�W]u���?���;�n�Г��<[�"�N$�;��e}I���v��xm�xe�v��mhp���_�]��(CG$
�㠒�ΐ���eH�Ɵ�EA�'O⅗^R@�/�55��H�ސ�(����Q\2h1��s��#	=�:��JE\�t����3g��֭"0�s��`�E�����<�}�8T�h>h?�M��V8:R^��7�V�֭�%H� !q�[%L	���p�^�+��M���Xj�+����X��������N�<���1j�(2���:`|I��n)�]�0C�lӳ���+<#/���5�WcѢ�:���
��^P���@&�~�h�qJ\�$B����k:t���0ʹ�,\�U+Wc۫����B��+���q˱C���7yR��?�=NW�_�_T-s1s}L� ����3x��geS���VF-v>3�R���	�]D�b[ʌ��5��eI�(i�]]�ƾ)�I��1@�*KC
���_C"�9�-�J]k(�W�}޼�r贳;w��B�]<���&	�EN������ln�������m�}���o�^E�>��ݯ�=��g��r�x��/<|�n�?i�ou��Ͽ����:v�"`��:�tt���36�tݢ�_>s���^/zE�S��/����7��-V��5��O��`��������3~�L�K�h��'75��#�%ͳ�]����8�M�1e�	�''@q�V�!&$<{�<M�9~�T�����8�$á$�I��5\>ԥ�.����eL�J���c����8�}��4�Dr�Ee�{�P$��R��y�?��/k9$i�9�~�-�2i�4�	��ň�3TD~��)Je��M$q��[���p�$F�5iR�b�/����g���44P��L�S�3�ӌ��ONϲ�a�z��ҏB)�a�ƹ��w�3�hr�cI|cu���=���OJf}�w !O#4=����+���p��p�#}�{�'�	��'�h6g\��d�w��,�P�Ys�tS��I�T��}�?����2��_A�5^�2`���#l��,�7�g�h:I8�`0#{�����m�p�S�9u�d�+k��+���kќd��֧Np	녘<a"��K�gv��	���)iѡ���&[&�N�Ř'g<f_�q�M�S�9�����>tw���ߎ��-F��%e�gΝU	�Ap��o��b��Zk��O_���1����%r�(�i�(Mڏ(m�4J�HU�R��UՏ~�_m�(j�))�j	y R��<j�+$`���ql���~�j�9�>�^l����Q��=��s�^{�5ǚs�1T!;� ��k3�^:��s�Zo���Aq۶�̔�����|P�T��=	��X!�a�/���87�G@��^�������}�#���#�?���9t�v��6��i��%%���5u�F`i�:��R� ��@.��������α��N��xN�#B=�Oz-�B��7�B���w���{����k=�����F9��ʟ�U<����ĊUS�R�ŗ�-��!Yavl�fnۿ������}�t�K,M�
�8=!�b�x?�.C@��A!YNٕ�܂RR��A�{��5ڰa=��/9�n ��އχ��� �dF�z��!��?p�By
e[���)���L�1e2�jl�o��P�k83h���'n���?��[�. ��k�T�ʝw~���~�ׯw�y6o5���磷����׽�e�����}�s��w��ڍ�n;u��:,�3��{���K�_��o/�_��&�o~ ����.��]w��R��nn6fQ�
8��7D�V�]�tG� �u����""&.��$#e&@��՟���k1��`E�9$4� @=
��5�G	�+�eBKQ�=�Z� -i'b��@��;YLr�/LLO�����.p4�A����n<�Њ�ra��d�SsEw(�%fn�.`@���	�2nX�Ȩ@�/\�R�:H+Jm���� ��&%[�;�IXhYF�
VmG��AJ��A���Ĝ}��RaN��!!+;j���Ea���!�&�:z��-8�Ib�|�� ���ŢÕ�H ��R�g���i�
h��k�#O>nN.-�Y{��y�I
�(R��ًKJ�I��7Ͼ�<��ˀQqA�%$̗43׾�}f�����)��1��bD@x��'�3�>o�H�J=��g�Ι��q�L��ѫ+�����1/���Y��������R��H��s	s�V�}��@����0�З��9�li�Z!�^�u�=r��߃K�<��*�����y��Lo�Gn��\���ļcϿz"���6U�P�_� �d����V޳:���� �\ ��បRB�\��|s����=��q�vnN:g`��]6߸�[B2C��U�v){Ŕ���MA�x&�Xo��{]rQ.�B�: T�?�#�Y�u+���"����\t����sT�)�-�l6 z}�?�`�mj����FpP�υjk^3&%Qb�U#�V	����9B'��έ[�-���;��Ǉ�0�j^���/N�4����%�iMLp#���&Wt��ܲ� �#B�,@ȫ�7N�4ӓm�� �� ��h�� �`ά�Z)"��C*s����4���⒉�g��5p"���kXι��frrΤ :��8;�t,�=_SsO_���?��?��ݿj@��������G�fa�mܰ�d��C7_��/~r��_�C�����������f����Bcjr����ܺ��w_y�]n���΍�����a��G�=���p�C������|��M���ߔ��h^#�!x %���H ��b�V��	^"' ˱�QYDB-=�qa��
�EֈA�Vs2\U����d@H9h/��ۣo/�m`��+(@��`0��'�XPy�b���x���3�v�
ΐ�
�s,h[����us��baW�c��D��3�9`;N�M��� ��`'�g��굀����"	G,} ��p"=�4���u;�,��&�~�@�>R��Ϩ�7*	T'�[t	N�V)3��J?�����#� �/-��O�l`k�,$E����s�v�`�4F��_��aFS�&��|�u�?�⸌֗Pc�T������rG����"Vo03�� ��Mٽ���+:�u�"-?���74�q�ff�����J3�t���BV��V��ɕ^+� �.h`��J���fnvƬ;k-���^?�k������!�]����z��^l��N�ڲ���r"����W�_�{� [N ���{�׽�z*�̀�ӌ���������U�]J1t����[d����w�A3@�^��:���
RF�G�C�hX=�.�a/w�X������P\	\�k?8![Ɍ���۴�.wLo�g~���0�����dL�&b�����:K-�P�Px]-�p]F@G):�](�����у�B뀳f��s��7�h��N���0�&�U���ys�w�cN..�e�d��"�.��O�t�%�����86Kfӆ�̇>����͘{�!3���i}�<�m�J[��H(M~Ԗ���]@Y@�P�v��C���N��H�D;�/6��4��ȎMk���?���^�s��JP��ѝ_��<����k�F۴}��uW��§n~��tܹ����G_YZ�����F����V �F�j����?�v����-����]�I�|�Г;�Av��c�.w�����ِڨ��陙�u�y3��^�Х�Zlq`1d�[g�U�Db������S����-i{�O{{�~������7@� ���p�W��x��u�6" e0�a�<� ΅�
-X�F%p�zn�1U��2���Tv��|ƮT/5�iZv��!8�	�E���Eo�Q'q	��H�K��A�*t��e�D�B5��wl��.�YA�&���X��ٖ�T nl�*qa-i^Wp2����q�j����'���Zc�ڳMv8Y�j1Jv�# (���H���Ҽ����+X�(kf	v��Y1���l-S�,L��ǀ��*8f�TPc��Ė�V�uNΥ��Uv���'���f���HK&C8�u���$	�P�#g5��j�A��&�F���i;��h�ˮK$DA��0gAPN�=@���%���;	�"��4|�/��}&!�+%�N�׶:���]c��E��)/+���CWyS�R�0� ��yyl~ޜ�i��u�`Am��e|>}�cI5����UB%Q�)蕠.l�P
�t���/��;K,�@	��fC
�H���0��/�
�J�;ΐ������������ob���2�"`��v��A�ss*8u���f�ٛ	f��9a���f{z�$H 6|�d���4Q��05�)��r���҈�9� ��n6����D��uS�1;�P��?q��!�0,�馩�Fn�&G-�=�0��+�}�y��6?�P���67�t�ym���֮?����Y��0w� ���߸�l�|6����d�n�i��桧~l�k�=v���C˞;t����v��&&��߼�o?sˍ���u��^ye��?����M���E��a��<պ��}��ɇ�^yZ��7t|��y���}�s�޺y��������i5�c��͇Ó�OZ� �P�7�����tVD5�_NMϙ��t�T�����g\�FK�� V[I��&��$m��I�dt%=�x�,�TJ���� љK�ӱ����������6�ա��?*�?L�H�xA$�3�vK�/�1��	æ��U�V\f���M�uK�Krb! ���r7���1������v\��'5X��A�Cg�L^
��H��}��M��K0a��P���)
�<>jz�
Q ����&=��b!(�w�(��V!�>���&u �I&CQ�c���&
� �A4d��'kl�^ VI�h��D�  �IDAT�&�ꇓ���sL�#��ʝ*��9u�b�,�_u����c|ж���<w�B��7�;�F��1�Վ��� ���}��� �`y�����+[UЪʆa�J>A���Pg��լ��q.p�B��-�IP�S�i� �{"���C�^�
�Q5��q`7K9յs�A_<0 ��=�����9�	�;�3Q���9jga�}�r�!5-�+l��6:���m��+�
!8Xt�6H�w`���y#�xF`�����w �9fgX0�� p ��D�\0`��qC@�gBa�sA�DHr���;v�(C�{p/�̆�:'f�֘���F �^O�KO٥��@����·�y�ey�.�B�$Q�;t	�40Ruò;B5^�8!D\4���K s/� �\�lh��;��� d�q��g��q�(��� al��MS	�$�����?Ef-1h/x����v����e[^���K�� �nM����	�S����X�.qs�-�;t��c�b>O���{ʘ��'�x���}�s�{_��~n��x��u�,�8qb����}w?z�/�z���5�n��&Y�޳����{��w��OO��_���=��m��n���ě56���=��#g�sv�\a}Dm�cd3�����0S4#�'��ћ����B@��/�I��Z'���.�*��R ��d���\�B�R�{��$Si���i�G�P }�4cؽ� ��h�tc�=���v�B�e*@�B�m��j�����`e<�u/�m�ާ�j��;�9� jm����*%W�(ִm�UP�u����r��H�9
f�:`�`��h�1��34k�gVL�����P~ER�#�=�wU���u�/l[T�Ӡ�� ����l�Y5Ǫ�\=�0�4؞#��e�$���aw���:#��*����S�}�yDv�D�N�C�RȀ��A���?+Q
+�}8)¬|��Ȝ�B���`�����;v�4�}Bv+�q����%�=V��C�~��W/�`�����<BF,�C�3����\5	��v pW��\@����n�YE&�i0J{�V@>5�U�|"$�Gٍ�~(a0ݯV����B:-V�L�?��OKbt=,A�h�)h���վ�ԉ1��|5�Jm=�I�x���)o"�Z��Łc	WSלp݂PVu�ʵ��|��^]�/}�+s������s��4-Y`#�n�g�5�Մ&E���Y�d�1!=FM���tش�O/<o�w�����_r�綟A}6�~~l�=?��?z����Թ |���Қ��{/��/>}��3���1��z晹��������X��ά�PoO��Z\O�"�i���|���TC��
��|�]�gQ���g��|�{[�Rr�`�L�w9�9�&�٨� ��������Q��(�����<wy��-U�x�(z��`�e%�,�@���905;�sqB~�A�L����ʝ"��!��I�^۪��`�VG ��a(�yx/HφE��4�]����(���]3�\ �{�.���u��<��>S����F�$���P�80�k�s$f���[�1��0><�+Z��@0*t���j��G����Uo:ί0 �����W�^��꠫c�&����M����\���ъ�rI%�З.�� ����̔,U�0�W=k]V���0�F?��uת�L�d���J�T>�aV�X��@J*��p�"\�PrA;�-�Ȋ���'8OP��@��ɠ�@�\�Q��yK�E�5q,,�{A���$�#��[1O��"j�\�������h��
���A�+z$�I�S�
�̛?��p;��*��+���Lڽ��>�f�%k� �_J,�>�I Ae`\ug���ѿ<Ax	�i)}��W8����o�a�{ϡ�Q�}�k5C�Z�	(��]��^�N��*P.{��L��_P��p�Ko���-�#�3z�I�����-t~�To�v������E���L9N��29=$ug�Aoã�����_��+.{ס��w�"5fy��ɗ�Y腗/=���W��;wnG��q�Y�״Z�]�}�?�x���ܷ{w������[������K/=3����'N�x���w>�QnҸH�M�9뢼�>�Ӽ泬��lP���Z�y���g�F�:D�3b�:�I(�P�Ҙz��<�(_xǈjrdn��Ȣ$+j�<�1�kHwQ-v��ŵ������"�Y8C0������(
O&;Є�	6�5����ρ48k��C���yd�� i�����}����y'7: ��V)�F�Dl���e�/��³$�ɂbڰ6͆j�̻��B��B�\�� �MJ��򦳅��b������9��Ta�΅�]�Ej.�#�DC�#���8���d�����wv�65��#c3n�(��כ���]�N;.� �p�-�ȅ�v+AN��縍 /�'/�_��N!���E�N��5�k$$��Ӑ�ňI@b��B��P9��$+	�o1k�P�������� F��6�.��2n�S8Z>��	x��"������@I$�;�U� L��;ĜS�h�D�� 0�Q��`2Z���V�8IqTmEsqK��~�e`�|��W/�!���.�U`������ #��Q鮚(WO�څ��U��vi����5O�{佡@�����c� �H�b��+�pr��'sz��#��_���;pXF�Bex��$n�+�(�������"#!BK����J2��~��j2���C�$|���rY���o ��X�N�{X�W0T�A�de���J�8O:[VTY(�FH�g�YS^���ę��o�ˋ&���5��m�tp�֭�l��}���5�{��G��~��׏�ʜ;��j�;�Jx�d���ɉ;n�����W9S0_}����~��Ԟ}�D��a7ǶD��"��~S�<z�w&N�ܩ�_����F�m�c��pࢨo��\��6]3F6v{��qiY4����i�N�܉~/��n4�	�M����#��=ٮ�"�"��כ��]��H
Dq���V�,�m�?g[��B��ٌWvh�\XvE�9��%���4�K2�Z��/NAб6����(b_ą����!��CL�?"<���%&5.�6�g�;�3���tX[3跔� �9�x%)^��@_���s��rNi�
��/��mDuȯ�V���|��i�D)9C!�a���\��1`�����2�E�I���Ys�g�T��BT)�321|8��#E��P8J��� s B�"FQ��՜z����!t��kFظ1lay�i{�Y.�mx��9T���b,X��D4�0lE�ͣq �0".���DF�ko��z)�h�ȑ� ��)�=�'�������@�� ���aQ���c���K�$�Y�QdAܑ��Z�>'�b��?ɽ	,����B�ZhvֹB@������P��𜧀kr���	#��/��
,A�\9��a�)2�N1��Ȥ!�r��������$Չl9F����� o�Th�3&n�<d�9�p��o�=��J��>�QrE� �� �r�gR¢ˌ�X0HhB�g�f����ןk�s�Drm��F�Ϲ�� �@J&N3"�#��R�!�,�8~�ș�0TA�%�&b����b�����y��QV܃���n��c@ԩ2�z��n���My����J@�r�J�����t �2�e4����ȵ$@cjΏ�$�C/��$p= Jc�8��&�O��ugNN6�4Mk�^w��k'����� FIrzr"1y���m[�}���_��[o}q��������}��������!o�i��y:���'ȟ��o���j�>���Es�����U�$��o����o�Y�`�$��"���.b�۳�N0b� !�\�V�L�� A��U���}�4���I�>�,���Ȋ���(�`���8��(q6uI�Z
v�rʟ	S([���0 �Y��aG��`C#f�a��E�s�9[�qE����S��6Ϣ��8w���l?G���<*��ߋZ�)��]\7��=��ȭMS���yƻa��
[ �g= ����H�v9"�f���kL��O�M���3�Cf,�h�K �rx���|́�9 _��ki;�q�ω0o�&����5^�h̙��pP����I� �~s'zdT���A�Y�<��涰��,��(xip��|v�0�Tc���=�@� 2$�P��e@:�C�L�mpM����HEB~_K�B�\M&'K ���t"ɜ�鬘T��h�+HGFS�b�5�%�T�� R�X���̽������m¯
�Ho���p0®`����6b�q���+ؖ�_��5�8��̋E p�c��s�@�"_�>���j&Q�Tf� r>�-w�8��f�YK����ljj��n5N��Ooۼ��}���O��{Fg��t慶�;��G`<�����* (�t��"��1�u�� B�Ѽ��@�l������Ѽ�)���C��. sd-�������.����s��hPG��L&q�Zzt0%h:�q��$��lv�,� ��#�j��\�Km�"���,r �|�'
��8���ˬ˜�v:��3B�Y~�d�2X�Ke�zG?'��QA,�%mT�mASf�md�l�dm�A����s��EĚ�wQ�fS��k�Ǒ/ QY�D~��x0L�
L���E���XW>�!H���*B�9
���) o����˛�!X)21�޺�pqL�rS� �R�ԲZ�L��XX�ۢ��H���;��(#���|fo0���Țy_�ٮO O�dH��n���E�V���5wn;��}�굽[��Ʉ�L7�x��kY��_2���G��7JV��ug�X��1�M�9c��3X �C�h���e��H@T���^�w�+bT��# �@e�����x0RYr�`� �wE
� :�,�e���{��wiV��u
�[{~�>��d����Ҩ7�$��h�xhӡ�q���f��8����(�C���xT"���.ק�ut��E���s������}wΤ��V�h��~�����#0���G�8�����S��x�#0�������h<���xށ#0����>>���G`<�x���8��������#0���G�8�����S��x�#0���������Z�    IEND�B`�PK   繆X.h�G� � /   images/f072ed7c-bdca-4b42-938b-e27227333132.pngtzC�.��ضm��3�m۶m�����gl㾛��M��J�R]���R�������H�)���BA�������vQ������!�	�z�_�j՚�������>Nq[$g(��ĥS��e�����1LK|N�d0��_A|��bQ[�@l28vvM�Y���TQE�RE�P�L�&s3�e��b�:�7�P�F�jm£݁Lľ�ow�n����\��2��]��@�/���~�s*����.i�? �����Sa�y�. �~������5`�^�m�n�gu�p��;�~�I�4 �~/ێ��~����
��4/�@�����ckp��:�um�%EI�Uv�Ow�i��u���+@�����-��uW� �U�yd�WF5��\i��(�jb۔%I���3	�k�*��)ķ�1�9Z�l������Ժ�7�k2�y34�TG����4f��W��:��/k��h�9��=�D~��['�������2��ع�t�������;�?�˿�?9�������|���k9U:��u�?[������qEX��likCX�ę{1Z���rq�q\g��T���"Y���y����Ȣ�6DZ��k�
��DU�Dv��pBc���Y-ĸ�м̍1�mY�
�_.���ۋ]*��e�Pjؚ���;�M.G^U���a<�����H�X��A}�'�÷F]�KٔH��`iw3M5��`�h��Xs�S&�3� �YN<zT6N�$�#;�)�\����c9�B��D��)�'��YI�#Ր�gH�[T-#��E�d����<�>͓_<�.��;C�����>7�.�5�E\u$1��C¬�4ZK�K�!f�߾����C�>Ø
̞n�"kF�ѓ�攞Amk���HU�P?Q2��<#O�*^ZQ3;�q�����H"[���1�ʍ#-R�F�L�z�-��w�pS�r��LY�k���bq��\��S���R2=h�Q�cE���8���&Q�)ga_{�~�m�	X[�^�p�	�m�Lg7<�N����+�dw��G~�NnK�b~��4������?���:?N	�*O�p��Oow���Q��h�/t� [각p2����N���,��Y�������Z^�7�&9������p�*�:��j���ۍ��Ń�E�G�@v1}�U�dШ�D�jfu5�⬆��d�̕|{�{��wر�n �3<����!�x*�� �OUK��W�éf��M�L����}K���a��љ�kW^�՘���p@����K��Y��޴$�@a���Sk���mN���A�cmR���dC�'t�[|�d������ݱ��fw6�˩{�w��tٛ���P�d�I
����mY+=�*��}���Y:N��z�t�
��'����y�i:�4� �k.�����$ǂ_�2�ۂ�����7���D�Lc�7G�����z����<h�̹!��]Aֆqu�q���m���T|�Θs���ށ�pM`De����T.�"�x�
���O��s�����)tpl��!8 K\��O4$�6�QyA��ǵ�I@��9P���fzh�,��f����W�,Nj�E8)�U1��f 6{R0�{�p�`���0pR�3��q���c,>l���8<�Cs�B�0`Th
��7pHJ�Q� 6�{�\a�q�`.����x |)k�a�Cp��%����K�9g\amx6��& ���<Tq��S��g*PJ�r���u���8����!ͥ=�:&��|ǜg�.�=,���L�ٗ��v��(>E(�;��6�<d(���2Yߊ�"�#<ꈭ&.f�K=az�zzdc��))�D(�4~�X
�{����xz��]"�.��,�qUL)/[j�F���(T%�#<���ƽ�NQ�Hґ ��S)W#ג>j��%�؟�� j�([e��)F״�١g��w� ��N�;�(�,����&�*��˟!a�Nv���
Jڔ������S,�"5�Dv�&	V��el7�}9�3D���3
r m"�u�.�4	���LZ�1�/La�=�d�J�3An�]��LᄓvBTuѬ������JKl��Py�.�s/�:���RBǭa�.g1�3>*�r@2f����I��h]Z
�ـ�08��gL����?��2�ڪ��>��1�D�<AiY�������Wr�l�Irs[������8��+$���h�{M��:#)CM���e�Qf�������]]���i�<v&ӛb�
��F�Y#R�&�x6�T�Q��Y���1	��y�d�ɮ!�L=mMQ�d�fp��:v�Z��Q�]�,OI�r�n(���V�V�����ԴJŕ��6��7�ta�)���h��Au$VS犓[Nw���%�F�	s:0+��ibc�wD�ȹi��(Hk�bQu����m�cx�<`����d�{�j�WL�dZȣ_xQ`���~w�GS���
4��#�E��o�f��B<����Qަ߄:��T��ԡ��w�� ��C	�.�X�A!~�x���,d0��F����\��PHs3bU�C�Im�Hpc�+�tP��B�d�����=|��iih��c�P�� �a�	�n �hN���Q֐Ib;��t6���VE�n�US'j�/�M���2���?� d��FdM=�('3EI�C��YС�%���a0up�4$�
T��R� ??����7�@)����:��^
Z��������F�2C�v]��a�[5$�}?��s�3s�O5x���f�Ύ�<D���-a?�1;��2~�����a�B�98�	�2���HV4��[�W�0z��[�V��@Y��z��~�M��xi@���jz<�x~���w�����a��-q�eG�b�2?���I�=c�F@�XM�K)WCG.�B�N�@�X����7��Z�H��/׌/O7�;�n���'�����������[���D���L������SI� e����Q]6�G$o)��=B�/C�+x C���3_N{��ni����p�)1"��=�;�Z�G���[.�v[w���(��6���U#m3�]C8��-�3Y��jU\I�����f�bb��ZH'�7�t�9H^H��qG����fiCyEz�rgSB!�bq��R�*>Ǧ�˔��:`OY�c�V6Y����rC!PO�lH��T�E%|�#�\�u��[*]qd�s�*��Mi��<����	�u���5)'�=��?x�b�]�&�*uT������ousZ���4���d���'�Y��VҚ��S�n��ճȶc?��-t,+&�j�sqh�yurI����8�u���r)�����y������f������#��q�R(�DW�"<��,I�7�k0�U���/�� �8**��}Uhwb�tSb��>K}���/{\�SK�_�\N��?��r!���*�Q��A�bRЬx�bpnd#=���gg�s�9�Wg������Dٞ���;�u��L	B�N���r͐�lj��N/�ڭ�cP�]0-O�
i�O�="���[F,�*���9�V<5��ut����qrO�ݎ�΢_�Ye��'��+f���M�lC�(�9���@M�ePң���Lw���Tt��ʠp�͈����K��/�D����9�}��ev�t�?ٔ��S�V��
�Q"���-ư�heFZ!�.P̘
���Ħ���i�mةJ��%;�� �%k	��1/��ݛ������$r�8D�p��Y�T�����o����#XZ{���7�5�}e �;��m.80�e��K���
Mfdt��r��/�,dۆfL�VD��_����h�hI��4���$���҂"IS�kS��F���"�p�2�j~E�1�j��a$o����7w�o�lv�TzO��}���)'�1{I�e#u����c���^MCq�\+"34{XP����PeA8v��
�J2�d����U�Zc��HB�V�Ku���A֠�I�j��Y��C������Kȍ�o�ծg�oR:���Y�33�qѕx�b�|%_]�(��Nol�=�:Ԍ\�MLQɸļ$�͸s��f�*L6	�1)�s���`�l6�w�U�����eQI�Y�mN4��<̼�ǒ��aR2K�餪/&�k᫣S�+s���ԡ{�s�7>{��x&����$n���fRϝVP�mq���e��A��GMG+��rJk!O	w�Ç���V3����:\g#�ie�ƣ�A$.p���d��U��e1��ዷc�N<�2�lX������%Â�s�tH+�W��(�S���VtQ�$���i����ȓ����PUn��ļЍzM��QBDg�Hl��t�T�
����aI��h����6��T����PPO���-�HH��$zR�e��Hy����9J�><�&�%����·��䱺����,ƪd�ɋ�Y�y3��^�I���.�I���t,��O,Ϊ��3$bB�'�7F�Pt!?�
�4���P:�E;�v�]^�:�o�ҥ�V��s&j�tFa�����$Fb�Q���n�]`{�*>��Cw�;����TF_b27�A����ڨ|_���P8��#��{�߭�J�\I�C+u�OڠS��Ԋ<��x
�Za���%�0��;��&��� k��|��DʅѕĊ�E�h��V<�6���wh�_�ă���2u�#��5 0�G���1��
/��q����aL����l&<�=�_�e̔���K��Lw���P�M�J�	a���|N����R��+Q�-����+B���u��]�&���$@C�q�	g�W���^�����!6�$��4�z3Ǚ�M
�k����V�̺��w1Ux�x�(����ͻdI��Ig�fm����dfg�����mͰ ���!R�K�c���vi&�cz��T����'5��z�o�C�r�� ����Jo�Q�N��\i�ܓg@����N�H����G��ePe_<JR�`?�s���Dk|�3�Bu(z<�f�����g��H_Ho1/gr@�D�,|d%����P����sF_��.��p�پ��b��=����p���:�o-$F,p���*�@Z_ߒޖ�֬I߽�{�?����I������w���35��GB��	���ijDΊ��������FoV���I�#�?�vVs����#߷���D��׭���@���\.Pa@�6��$�R��S�ښ���<5����;�5�@�R�=C�d�GηP 3m�N��l�a�$��NUh�b�7�ƪ�9��3���8_d7�daǃ����
�]������A�n|,)(&���yd��Iܨ�"��D�Һ�58X�4�"�dQ*M�3�H�� 
����yrf����>�:u�C.�*
n�8ka�������[ǫ�.�8"S�T����Yǟ��t%�������wR�É��R����Γ�Io'o�Rf�O�]Kr|ϤTj��]��X)l[g�;	7���{��d��J�b?�FOP���	�����ʯO<�#L��E�w���1'o���ɛ��ӯ�i����a��VHP�'�U))B���}ER[�� 3�&�l�A�U��SO�z�>��D�XDLw%(q� �zР����WH�\�*�J�����Tڸ�Q�b.쵬]��2�N�e~�'B��J,@��J�*��	U��,Ӄg!��Ee�{��V/���	����vS"�7'��zV` xI�	�����&�E�W]ڪp�o����)8��3�g�py��(�ƶ	[~{�mNzx��㬓��B��x'{�>��1֯Tw�	����V�����㯄�l�"�����G�P^kD�]߾��=�֗&��Zq��B�(��t�ʱpn�@�b99�����9�9�6�)%Ji%ϫ0�6y�X��PQ3a��Q����x�g��2`�D?f���[��ZX���<�`󍸊D��]�m�2�����p��,���M�����T�6��ۂ��2�Ð�◭���y��Fp�gC�s�|�l��#9{N� {� �"�$�wm� �p��t`�JI8�G�C��F�F1[�}�����|�56N�����jٖ-�Z��Ս���́r�s
����6���Y+M
h��B� �٘����32;a��ӑt�L���CWraD	/^�A��w��=��L��k��ܝ�_�X
RP�/Z9-F-�(Cׂ]%zŠ�����t�)-%KDA`>!��Y �Rj��͕*�28xuDxI@�����{���AJr�D�B��%ib�?ޚ%�"�1
PP���%J{g>�Gk�YF�
U2�TV��
�
�8��ح2c��Z;�C�S#�п�)3��qC�I����_�7�5 �W���N��G<�J�RW�ഩK�1?����V�*�!Z)�'�� ���Z��t�Y/��@6h��9A+��9�/�)�T^����ʯ�'j`xm.�_ӘBD7O��g��}��`�ْ�����P��%�f��&�Z0Q���x��� UpW�7�W�@Q_'i�D�V`E��CY��+A�Ғ˒E>���J��E�xg":��6�@8�E�w1+2��uҵ�3|?�v�ך���JN�P�j<N�>�J�?�����3MI�~���'�\|Y�O9P���g%!��f�
�	a\�W@7�@N'7%�T�g���亝;��D��|�0F�ÿ���1}��u"��`�;�J��I��7�)��ħ��ҙ,��=���^�H��[	��% �yyI������ߙ��>Cl�	�)#�g�^{�����>���䵜����wɼ̭��l_VQ�w�Q��2H�# *�����D���r����d�u����!���5|��ʭO�@]^I�gą�JT�w��\�׌�Q-�A��T�p ��Z�  �p�C�M��+��?���;�[=%L�̔o]�VK��3�ц�e�#�r��+�t$-*�L��4L(�r��~4�_�2�5фچռ�-�
)�G�3�����ұ+e�E�p��~"�1��3;��p��3�#p/I��z�)�u�߹C���j�D�@�#��9S�o��p^�� 3�N�	͈$�9�����s�a5�z��A�qy)�P3%5w�I==%V�%�,,��R`�0�l� Ց	\�R��3,>4E,�w7�h�P�	>O�7�2��Ԁ4��g����[?̿�U�q´ r�D5�V.�O�-�䨳q��xZ���"��*H�Aw��l�`�W������,����o�C�i(Q�#/��z��E�MƄ����U�t��}`k�����c�n2�z���,K��+������j]4s
N�>5��γu�»�bAX^a��qS|U�Zw����$�{tN:�)�6`��%��Q��~�wkd]�ZA8��P0�_���[��A=������J�� �0��q�I�6���������������ne�C�1;Q,��x^t�l���	JG1V~�ص#��S����J�[H�/�K�h�VJ�H��Ӳ�<��7����é���@뱚�|�b�	��L!��P��^�r�'~y~����'m���T�M��<��"���Ի�	��i/�0���m� �zPҾ�j��}&0�a�-_�b�=lIl΂x��y5a��x�/���_E���x�Zb��@q�,"�/ �a؎t��@@�����[j��^�_�H���OQ+�J0lY�8�V:12��r�F$�i�&�l�ʃ{���Xӹ���ɻ��/s�]1Sep�>��v�bF7�H\>&��$�,Y��u�|����o
��q�LV�
8	�
M�d��"_3���+Y9Y��/�O�C�K/U"eU����0�w���
D�M�-93Wfnwۼw5[��,�
&^�)������*b�A�0����aRd�B�$&`�I�~�����-q����	X\+�X°W��Ʀ���V�F��� �o�WZ��U��ҷ�̬'R�=r��Q�m>���Km0bwv����z�s^D�J��ڌ:�8���+�@F!w̄2�$M;S�zX��v�Cf�E,�:�&���~V��&�Iŗ�G.�	z>a��R�ϹBH��r6�-�>aQ�W/����F�Z*�J���߉BM�*�q�(�لY�1�ĸϡ��\�y�^�b�(���\ �j'- ���S�H�'�r��.!���B��=�����(�R�����:](N-����f���djs�*��3�w�l���<��,5mE~i�()���?-x'�H�̭ϤX��L{���>+��h,ï,��z�Au�Fy!x�ՠOE�Q��BL9R�<�M�T�X5����Ɏu�e�D�HeȰ��f[��p<�{��L���G��ٟ�@x&�%~y�?Cn��~/�V����!�$�~�0��{b����1�����vW��M��Yz�E���.����$FMR%��O���A�ͱ��Zm�xH�Í��W'��
g��[�W�&��p�+GV/k{�u�#�!RR�ͳWl�jgA}eQ���l�q��vzqc�t%+�����%���.@Af%���9M�����s"8zH��<��ߘ���{lF��굗Ǜ�A�]cgI�"����@���wJju�177O.������Ɯ5���)�'Ɋ�Z���2G[2��t�G�^����̷>��������1��TC��ǚ`?��*Ψ�d�v%r/���`�聜5�l�1~LAlҥ��X��҄�6�x�Δh���r0�w����՚�4��ct�#��nT�� {^n�.��5[�!o.±L�LS7T�O���8cj0���I#J`��a���w���g_�L��ǐ˸���\���.�!
�e[��R[Jf�@���_~���@/�K��v@���%+����
�>�=#΀T���c�0�ϐ��
ȷ����ٲ@�G&��9k��2�����z�����"�l�|���
N��,⺫!�4>�cK�#��u����}�8������I���O	x�Q��d��O���? 5�<Ik��m����`'�G�ot@�`�������"�SA�OV/b��N$�T��7�*7ӻ���Ż�B�դ���p`�b9����M��w*�H[��/���n�$�~x����y���bXF�&��������� �T�4K!Q)�S!O�O�Kx�F��䓎Y��_-G�X*G�$�shu��%���������L\�]��V���:M��ٶ!Q���	-�Y|��I�c*:@D��W���F�ӏ�fr�>=��!q/�\L��~��C����������nWi���R6\9����,k4��Z����������%�!�wu<� ߌfx
���GW����/��H�q��0���v>�'hy�0v���u>Y<���.�[s�Fʕi8��Z��hY��@�;�w��O���W� ���M�k	*/�t��׳�[�k�_z�g�!����t7.^֨Xk�CD���9��G�n��U�ݘf¤	��UnJ�$2� ��i�{��]��)5�6��X�.=���x�M�$׸�� !o��x�����*M0~J���j?�]}e�%Tȼ��;\R��9&_I=�Clra:��+�H��u.�� ���"3�(h����n�qw�ٶ�S�˱g�@�~O�6�����+��ٺr�y�i���X0�'���=^%�E���i<��I�W��Y���^w����oT���e�[��Mw�������̀��慎��r�s�-�kX-)�OV�D4�����@3S���9�P������K�H����|��Ec8jD���ϫgcC�ԋ�!i'Z�܂��	V?лl?7X�7���|�,�l`���b��8�(��Cq�K���R��L�f>x��5b��<���
��1�Ba�!�9%� �'w��ppHY�ଏעԿ<(��[QQ0�v�Ѩ��i药ᴷ����dxh���b"
TH�dC���!g���=/|c�1���8��bY�J?x���p��8=;eb�`0�}���u�9LQO1]1C�?7��"��=�O��7!q9��>��O�hhh���y:���I���I}$_&��hV�>j���R�5��2�\
J&����'�,�`�g*��������pz��eA�"= �	�yah�&�X�X��{�!K�x5t��sSS�/R�_T�x7����
�9������x�i����9�����{ɱ)�7�NSr�_Nn%�<0_��\��w���l�R�j��Ȅ"`d�6҄��TaF���D�-�CI.\�
Qe2-	E��9�n<�]�h�.M	���X?#���q��L�yw�V��U�qk�!�[F�4�L`�A�Q����A������@�?��D�7F�������`��qZz����N�\���_Dcg�Ga3�Q!�bk^��Kು�,)aM�\�d�X��qA��6���|Ņm���P���D2�.Nۛ�-tòɴ53쥚8�GDnn�6����xxoU�9��IA�\���r��@7�{>3;?���gk�>*��+p��E�6c�!#� G�	?V�;3?k���b��a�4�<3;c��+2���3<�7�C)gұp�1P�%��ѣa�	V�v�H����g
�[:��>��}EHj�p` ,V9�γ�qW+%O�N[Ӻ��_�\�g&�A�g��ܼ�b��7�=�/���47v��r��9"\����R�pz�Rgh��?mӦ��Q������#�"�oqȸyQ���W�����QE^<#4���:a�D����BϠ�_f9�<�ބe9�K���/Sy�A�.�0�5!`��U7�(pǯ��b�k8p��ۖ�^<X���V�-%,ؾ��^�� �?�o�v�z}�_��*� ��wE�����-<�g��w�c�z��2屏N��.�2��m�.�k�������rB���)|W�?�L�Q��/&N����Zx�`jE+vF�a��w�(�֑[)����U5�|r����C{���r_"^bݸI�KĒ5З)K��K�N踳���:�1v����h	�R3��zJ|60��M7� 6�i����Q�8�pf���a¹.=\���ޗ?Ԏ\O�ۧ��ñ��r�J��4gԝ��K���7p���c;!�:_x�s���\�͹�Ø��5����+���󻳃b�[�Tm`�db�uT�A����M��P������n��֧�� )�H�3#'ʢ��B�7W�.�����O���쌺�ױ��X��X�O!�O��b!��,g���t2Ujk��@�L��;N`ɜ�y�gZ���'q��Ѳ���P����h�G �|� �P�!�;��w�M�~x�썏�h8�lGtx�Ɨ��!���py����6�8ͳ���Ge��k��-�A�=�XꕽDɨŘF8c���dȸ���C#�/�I˟P$?�̉�(�箍�8Z<��ׇL3R��9)ɬ�e|/G-�����4:�u8�O�l@�'C�g�o���f��f�q��8 j�
w�f�Tr���w��I�k��\d��ٱZ2-K����`Y�me�#d7����:�-�/� �9��3c?�0N͙��;�� ��+�8��<4օ���&���°��ϭ\9ԝnz_>2�
F&��
UV;\1��F7?0趮d2D0@�
�[ՅQoU2s�i�6���U��O�5k���(���Oy�
n22�����!��h��ﴆó�f��(�8��I�C��A� ��XW�R�<��3���Q>�@p�3T��o���,N-=�+K��m'��Q#������/Q٪�����Dc�oM�L��.I��]󁠲����_��ޱ�^羂"������r,>���9b�B�F"/,�3ʶ	��0�hf���#�&��	6��k6���vh����A�Q�	ij�&��#��2T�Y�a���8�_��,����Y�莮��hn%�˃�񺵰舯�h�{md�2��.�)�<�:�����!����"�r���/���IO�J>�Y�U�!�8AR%x�D�X���b_�zuv:#��W ܽ6ZHڸg@�-T�( �o5Hx�1�yQ�b�K�;u]\�2�i�Z��D�=I�{%v���E/(b�m$"c@�2`���\�u��̴5h��if�q!�����������B��uׇ���4��,�H�ĉ��vFe�P��B�h��J�d�F���Q���'o������#�y�2j�eS��O+�D�
x�&U�:�r���w�*�덩����G�V�����
���.PD[M��aoo���x�ߪGD�yL,dO�P�W�{�ѻ�K��5���G5�Up�m��q�����Q0^�zn����NJ��i��H�����~i���sG�������7�-��qSO4��]��Ō'�	��`0����i����yp�����R�D<����>���U�-fc,��rS{�Dl�Z�|+�6��0eղĆ�����>���^C�ߡ�D?h��K1I3%"}��X,����~�&
5�(�O���r��_V��2'�#Шn`6��y�%�4�00�'ݣo���{s�$�e�lC0��Z�,D�eB�l�7�o���c�}����xP ����� ����C;��oZ��`���-_t�������ш@��_����f�b������u1�q-5Ŕ���,�%/��]d���� xN��b��`.F"��,�O����w�6��l���!;Z�Q:P��Q�q�<?!����|y#}K
)u9�~���0\��v�ƣ��E��Gf���%��"�gJ(�Ӻ�.w����v�����,���������8u}��#���	�n�����t[�lL������[�.�{�פ
�,ؘ���.7���[R)k	���;���[=m1k�}��R�I��0�|�Gx'E��+����eσI�Lk�u��4�5��];`tH�!M8��y�F�?dG7v�N�q{7�}T�=?��{^v!;���x ̆`����Q|�	��]���ޠfX-/ȫ�W¢����I#��9���2H��)��	��$*�/U�̬CF/zѡm��_W{ٷw�KD��?��������gȟ����]���o׊�!�
�O5n@��|y����V��⌘��>T%�lF�.WLaaYY��(eH�rR���6���:�=�R	�&.��?����2΍EJF��LYw�U(�\Ӑ��K;�I'�_�@�X�_���m��3&�?j�M+<��f�3��A� ���"ʺy�Պ��`�c;�7�[\~E�k�5]�-��`��y���ji���ob�Ab��R�k�;�d��8�8�\Y�S�!R�L\
�Ӌ���R�/sٹm.q-9��:<>l�
�xU��g��P=�߈c9�kw;�yd2�-��jݕ��nV��p9]QMS79{���a6�w�ЏV̥gb9:��7ĩP*H���t��{��D�@�k���G<���@���I��m(��Ԓژ�{8�^�n�be��cD�x�j�*����s�����ז��;`*�ތ�%i�uoU��3�huȰjԘ��j#����m��
W9^:�+��X��H=���<V�,�I�Y�����͍Z"YO���������	����r&0�s��а74P�P��em�a��l0�cY�}<k۴<^���2]~\A7&]i@�J�t��2��o�hk��{D/�������m�T�61�����W�����z�c_re>�/���Č/�����W+BS�lQ�3�Ǽq�����fiD2�jⲿ�E��Vź�����q?���oF(u�����g�/�-K�m�_<UE���E��	
 d~��>mI����~���~��t8����ݣ�}�a:���2�47l���s�5����z=a1�~����D���������qL7L�6^�02^��lt��2�8P�?%���kw�eC��MzZ#Vp:m4�C�����00�ĔU�n�v�J�iy�����`�/����\ń��/T�CKi��ooF�a��$$���3�V�u�u��;�&I�}5�h
��'B*ͩ�p"�{����=���U[�~^x(p X�V��)n����}!c���PNC�>�>K^�.�����8��#!�t 2C��=IGI��+)
̫͂�d�4�  ��!U�l`h���	C�G",��J��I���^tЙQG�� ~8Mnʌ���q郜η3>�Pd�CGR߭�=���\�.=V��ϊR2�tj[�#u��'����1v<�@`����\�~U�R�>+(>}�κ}� �H�L���7A%�rYd���ס匿tVđT�1��>cM@�O��.�7���O��9G��ǝ�jJ*3Ů�$<h��:�u�v����m��}`�L�ܞ�~�gp@��92lIF~�E��Z&_�33��O�v�`Qq���Ot4jc���1���������kp��|og]A��ڑ8��=}NމZ�C߮��[o!��N�hDD[pc\s��r�X�s���Jo����Yd�M$JǴ1"Х�3���Ns��2�D?���T�DJ6�X���D����_��2�6G�K���/&��B`b�р�0�1\2�p�Ѣ`D�6�g�#�,�-��UQlQ�Udt��=!�C��3���I�Z(9&ư�Q�R��B(��>����W�4)��+%0םt�����e��h�:Qnv�r`^K*k�/)�b��)|oz@N�\�wƇP��Ul�]|�1�_�ګ�d�BP��"_��Y���j����`���s�{�z^��[�J�;�pW+���[�̟�n��߇(4�۽?�[���[��t���E~>����>��c�����vG�����:�L܋#.
a��&�p����{�}���ܞ��I@.�e<>fx��Q���Ǳ
��Xë�����x�Ai� ��jL���o����y�6ʾ!����92Y����ۇ��=��6�K�cm�������ݢ`�)B�p�f���ѿ��eĒ;>�9�j������v�J^�3��oٞ�]��j̳Ǟ�O�[���y*P"v3�x��\�3�kWPfo׼t]��0�xdD��Qjds�
���?q߻E�V��3c##h�뽐���t�ϱ<����]m�hEqj��
�jgX���[�^����,�:Y�g���6ʊZ)�>��R(�6��_B	H�>+*����F�+��Hu�������m���R3 ["�9>�b�n�9�VfX&*P�r�1��/�7�����J�yF�@�<~_���wyV�ѧ*��'͏�����Z'�C���,�J��ёބrD���Y�.�z(�sM�!'��ߙ���0�Hz��l��J`��m�K��-
�cN´t�<�o�>	��!���t����o��{FƷ���y?���|�\<v��z}oAt;���c�
�<HB��[���}�\Y���E1��
�~���sPd� Y��;V�Q�{�����{h:"xl�a�� 	|�02�/0�	������@��T��6�}���ܲ�>�?�puq��F�8Y��G�Q=�źd�C̦�v�V:^�E��݁��Z�S�%���� ���^g/Ӻ�Ƅ��2� *R;���У	�s����~�g^e��ᚽ���������gF��r��O��OzvW�%�9������˹���2���8�g$�<3X�������yާ;L&�F���ͧ��r�x!ݐ�0g��z��+�d-T#���z���69�1��G��<}�y`·T'�<�	8�q��!%M��Xv�i\9G�������@�qD#��(>PNwT���݌�����uÓ]���\$YT��<W�hIMُ]^���F(:j��Y�8�%(p��Zw�� ��ʊ���`��@��ytӤ,�_�S�,�:_�8�w?[�G}5?���eJ��Q��2�� �G��̬<�PQ{,�=��Bcb*=�����ô���an�~���:�.�6L�j1#�^��8>(�JLU��z�7��Z�K�p�C�Â��C�����˪S�7.�M���z�O�'�0���T���;�F40ㆸ�8��R�W]���B�O�m�(�4�
�hO��~Z�~\��1���P�86A
�zIaɩU��TG�W1��=(v�Cd�1�1�C:$vG�lDn�AK���M�u���h�u��`��SD��� 8@ǿ����_��x�ٳ8��	̌5��G� l}�C�>�_S�lɧ �⅋��{��ڵ2㳳P������1߾S�`��l[��eqd&�����NB�k�=``��ѱ�>����w�sM�a,�����R��^��6r�j�-auXO&��gץmy~�!���p����E�t���c��Ĥ8��Nk[[�x6��i Ҵ#��ء�8z���?y�ܹs�X�g65�XZX��0�k�븽��ݟD�I���8�< b�k���:<v�(66�q��=k�={�K@��lc���� K�-<r� ���=�\l�����=���E3o���+/�����ɱC���;％�^z	���$k677�������c��Oa��oh{��aK`�H_~�.��*���n|&fto�@����@?
�}#���O�()d�I�����o��W�-0�ehMLJA�cǏ��GOalj^�����_���uV.iJfs�	��\- �@z��!�����Z_�St�#�ֲ�}X�����a�@����3@L���Obi�w�JD3�ޚ�
�����x��>�4"Le��*�XY�-�1��F>���Y�Y��[��E���	�^�
�G2&�*n%[Py=M:+�}U+	�p�C\������c�P ;̖��Mk�GɅ���S��;��:\5�k?�1.\8�R�F.��駟���E��ͷDB��_��[���?x	7o� k2Զ�g�}'~��+7na��"�9,���?z�V�(i����<����H����5"#��Rgʇ��.������D��c�Dgʉ_��kx�7D.����5��=�p��a:r9�;A��w�A���i��b� ���o6/��^oO�+�/��P6�a'ޗ ��������������.$�#J11�v���k��~�=T���=fe�P��7��z8߁�5;�����Bf�,&�s���������-���!���_^<�g/��o���t
�z�����Yx��<��,-,���b�{}�8���U���V�*��$�
��n�;��<_i��J�`S(
��ҎǧC�{���E$�Du�u���|�d�c�ip����� *�S�Kݸ���(�ԩjq�p�Qb�"�n�#l:�ȇ���=3`5;��W�� �j��gg������u�h�5�&{���Qc Cf靷��cոi��Q ���'î(|��o3Z|��iz���8�7�D��)����2L`F�cY,ECuo�s���?�g�|��F�2��k]}1�2���y�߻� `u���>��n��������l#�@��fύ�:V�r8�a�/nH匴�L�L�#�{���9uF��:�ئT
��FN�B��Ͼ�����.��Ho$�&���c�m��R��j�wz�Ӏ�vQ��S|������v�b�Bז�D����&�qjљ8�����U>t�;����%�e+p������/>��ꗱ�q�>��ܹ%zh�C]�����7X��W��,˧�\�������>��c\�|yؽ�]�8���i�g��e|��0C%;�J
H�?rJ����n��7�ĭ71;?���%q,Rx5(��tqo}[��.qzfF猣�.=�M��f�{����� 2o~����#�3�B�'#�{r�<�.� ��T�^�
^BA�Hq$�S�Af���\�,�'0-Y����f̌�:)�MhzzXDO�)N����l�ۤw�b�V��#�I���IɊ1~��u߂�s^(�K��ss9:\aa5�-D� �
���B<P��ϲ������1��K���ۅ�4��G���������	��Q���;�1�}���uC?v�vD�u����G�*�>�k_{�=����N�����r��)p���Ӛy��k�Bg��jX��I��>z �墣 ^���<��$�tƱ#� �o�x?�����{�e���Y� ���s��??#�x��gp��m���O��;bG�]�No����C�|�"(>���~�_��a�aP �P��E���_ �o;-,�g����&%�ZC'��41��f��H��]�j�3��`yv\ |�����e�l�{�괅]^XZ��O`�EafM�a�l��]��|o���V.i�E����l�me=qd4��{8y��C�,� �K��Ǒ6���W�]힯=rU�x��	��o~]:>���K�x�S�/���g�>��O������[������_���w�W^Ž�ua�)u����3g���c'p��sX���C�C���/�����ak����)��S�������h�O��;��v��%y�VK���9�.��ա�aX���,K�?��Oq��
��X\؃��y�ǔ����+hooI���V[Xx���u�I�;����7J��`��6�9@�)��0gE���O��3{GRЯS�k>S>+�������Iq���iaC:��u"�@�h#�X2��$����Vb�L�j
���V�?�f�=m�F6<����s����?~�����z���j���(���>�~�a,/-b~zBXh�i���	��l���o
�Z�3��S�a7ư�� L$�Y�n��)�Є��)jA}�0��EAY��E�{����>ٔ��N��q˄�;�*��QRm#������uZ��@�L$��BZJUh��\qS�}��`�CK�t��-G0��vP�@F��:�66�th��`a��XS�m���ʕ+x���ƍ�����4���ޕL����v�muZ��PV=M��xtԯ)ë�E"P��Q���Eb�d��*v�����x�o}��8��)�����lbjbL"�������n�/{�S'��1Zm�qwc�(���� �����n#�'�}�~�#��]���4��@�AN`~麤�E�ԹJ�8�Y���M�>m2��Ӫ��	{v6�l�$�X��$��n���?ȼȼeD?ҥ �h��N��k<�M֋��G��ҋ<G������P>�>�G+�SV�d���[��կ�����������ҧ�%��<dG,p�J[B��x�ӡ�G����=tP�U�o��q�;S�l�Ƀ��]�l����$X��uE �[���x�g������yG��O>���%8�};�L��Ɩ���?��[�n`���8���z�޸�/�ۯ�)�1Q���4���9sTK9X���8���Np*�uW��]����߯Y�����V���6����)c����uzjJ�;���֦\{�k���oI:�s�m�qe�E��P���9�f��^���o�&���OiYK�>�YA-�3��By�,β�bB���,xe+m���P�{Md��g��KO?���=L��h�t���x�4���5�Y?�H�P:��/�t&����Y�l>l�o���T�t��N�ϱ��ow��U�n��1��C�p_���Gj=D��m_C�8�+E|H5�"���~���u�����=ޅy�X�ǋ/~g��*�޹���'�rku���ƿ"��d�+ ^`�j䥈T��PӦmG5��e�(m �e�v�"%a�=��x-2��@��"U �S"�M�*��g���D_}��{�4�gƑ�����&E�'DB�� ���X������S����y���ӛ���[����l�`��X<mq�(N����F&�ͱ8l��\��K֮�̇�3Ȱ�����S�;��GO�[_��tz{��/���&�Hb��/�K/<��=�t�������x��p��%��՟H-�ɴ�l6���gq��a|�޻�s�6�<�=K�q����ǯ`s���"t�%�{������������;eR�֟0[��ޖ�R���>���|�pJO�1��G�����K�_\�l)�/̦�:�N;"�.t��bP�ݥ>^f	��Ɗ���r�n� �0����*�3I�۝���^r�	�$Ť#��R�!��+ rn�2�k��(49���]��RЃdv�7� ����ӎ��PfK��MH$Ӵ��4���t<���eC�}�/���N���o�ᵭ�Wze4N|5ТӉF�>$�߱C�%UX^�ozp(�J��[��E���T�硌�F�Lgy��]N��V�BO���Y��^0�5����� ^5��&���kd�C;+-,�
|4&�-j��6;�X"A���*����h���&t�3�sX����Q�4�Q��֘gʥ�_7����A�-�\�a�)�޽�W_~E��*+�~J��h��p��[c�~���֬d�-��p2eF���Jg�n>��f
��f>؅dD��{(� ��6Q�����{��<v��6"��koj::���qc%���169%�\j�;E����9~���Xo�-د�!@[3_��S�sSy�SR��vP���&�@
��eȺF�PpB�0�tB��%���}��D�b�+L���7��X�N��`���ЎJ�?���6����JԿ��ӷN P�s����P��H�P~�܏n����C�f7l<"���m��*���~�/ⅳO��W_�w��O%��tb����,�ދ����=e�EN�^�����ټ���_�w��]U3�Sʺr�,�*����VM!7�����������x��Ylon��sJA2Pl�z�򳾶*c+5f�Ν;���yϜ}O=���������؆�R�4A! >�o�Ѻ❰h��X��
�w�^��}�}`���S�7Q[�������F#�%Ac��ز��8&�a3'l��D,R4���6o����~vY�-чe)X`��c��A+�-����A�ۂP�
�b�ec9��"�j��
m�t~NӁ��׆-XZZD��ۜȠ(]ʛ�Ҫ�G�~�n[�����x��SظwSc9�'ٓ�Y�D�0\�Գh�]��I�3��4��e_�4�{�tu����W�&!�B�0h۹�y�F2�z��E�z_�`߀��@$�vi�@m�H�Yk\l�w���x���e����3m������ܗ_ĥk�����Y�1�M��Z(���=(�Q]������A��;"�5��e�J�M�'E�����HJX�>,�g/lW�&ZDҤvy�� Q����.��]J����oz_y�q	���M!�z�o�a���{��_���,M�`�C���fЮ#���Kx��wpue�����̩&�g�X�H,������}��U_������uj�Y?ޢ0`�7B��yJ�8��`�ģ'�;��7dw�~�:>���t�i��aiiN�~Dv�}�����＋���~�y|x�#��G�H恲A�]\X�W^�29~?�-ܸv]��:�s�>�?{K|7��M<���8y�1\�~]�y�zf�8��h�/-b��"���dAvI��&�$d�������>Ź�>B�[��N�YS����1>t@{͏5�冓B.��'!*L|D�.�����Z���fYl�o�&vST��s��vu���"J�1�)'5��1�
����;�.���L�Mw0&?���>w��0?����`�:x�����&v$��-[��KL�/{'�=l7�>�X��������Í����"����K�fd	r��������ʲ������齷df�%�E�lOu���%@@��>�{��?i0�0�� a����b�X�6�齋4��}<o���9/nY5� �ឹ��}�^{�6���ıC��ʉ��	%��Z��Z�m1�ݵ�n����q���O�r��XH�0�4��3��ʞΛn�ޣ�>���Sx���+��D�^M��9����#w��ԉ��+d
U�R�FF�X\Y�
[A��(����#B���D=�xT�����2��g��Y�h�g��g��V��K�q��u]c��r�-f�6#�	L�>�%3��ʥ�ӝG2A��\�44�N�
���kY�:�uJ��9�60��4����*X[�Gym�}=8}���j�^ȻC����ojc�:!�4�	��.�3N�.`�X���\¥�w�\(��w �t��S�*-Փ�$���\�`��G2Y'W;��9%��D�iі����ƍK
��?��01O(�I�E�+�I"��l�G����⴪e��2Zr���P����w ����[��|�Tp�]�j�/-��+]_��u�!RC���v=�~x��y�$>���x��;Q��V�9,$�F:�B)"�3?V�h���G�ñc�4<������j�R݈뉈=�O�²!��$��.��W��1^+�,9D?�яp��!�O�?UK���w��õ��0����s��+B�����̙3رs�:37�>��>=��9�h�����ƷL7����� �����>6&B�)�C�;�z*�|}vN���<��Q��6��!��&&�]�z�HLN�}]ݒ�e{�E���*&��E��F*C��JD��o��Ny=G_���HD^�� ��y�I�.�)�[,��IE��o&/M$��'�rU��<4?��*���Z�)�1
!I�dq�v��:�������zs���JJ��;�><GT���]�����0���y�D���P)VK��Y+��S6�~<;j�1�f[�^�c�x��.v��Q������0ɐv����ϖ��k�+Ҽ�p?����������
�Iee&��>5��YC�/�9�;u��w���_�+o���O��?|���2"�sL�C�^���su}�b ya-���Q�n����p%��,�*����Z�_`C���w�se���΅�Ou��P�ȉA�O����x��q�����΢Q\E�Z0��VSjXvM)����u�CX+W�����փ1|��7�Y�y �C�C�L���	���e
�f����}��O�/�	u)}j���]`�4�=:��$ϖQ�đ�x�ܛ��JK���.�e�����d�)n߾��O'p��9u%�u��5�{��:�>�=�w����bݲe��/���kױk���Xjk�\7�=�zT2�C<��A���T�@�XX�?C�()Z��t�x���8[�������,.��������ڒL��ك=�vk(�L>��^�ucD���̽l��ս g[�3$�=�|�-�R#Q�5��J8�6���)�,�ןg�*�6�SOZc$�ևb�� ��� �$*���	P�Q1���|X��(j�,����F�w�[�OPhƶ��G����b���R{�Xn�Yk�^��bܺu+��ٍ����(MD�!�(N��T�iNW\U9����	�%�V�� ����:$��N�G7U<�6�U��_7��^���SZ��/�9M��	�m(ڋ���Ɠ�e���������E�e-�:�H׌��V�(!e�hǱZ��C֑$��A�]-A�J�@.��@o�����������X��[����xeDI�iVJF!qfU0a���h5�}��ݹM�����e:���f\^^��}�n�\�h��s��m���2gg���1��ep�ȁhD*X���)sn�T2���<�oߡ�&����"V�eܸ� cO'P���EG���q!g�!uy�F�ˇR�\a�f�4ppn��ݖ��-)2IJ��[X�$���\�,^a�F�R���2�"��H� �� J���
��U��D�̡�(�f � ���� �' ��x(*@�����Y�_��!�u�U��Ù�C�֝ ��i�k6���0�I�'％w�x>�D���ͣ
d�ǟ*���U �C�-u&ͼΒ2�e4l���v����N�J�GG6+@Vk%%b�=��$��k���//�M�\+��w��ɣGѬT0�l�����׍o._ąK1;;�b��^ũ�/�y��}�߿�w�F����M���O&�4�׌�Qs�_>(��(�@��G������U��w��I�-�Mڔ�H��t��1wfLM
���D"�$�6�f��h��1��j�2�f1?7������J斖�Z�"�H�Aԝ1� D���������z6Kt�hJaBjW1jf��A��â�i,,,�D)�J�E�.�V���~}yMÇ��ȝ�    IDATt'�Aqq�C��ˋR@�I�t54S��"�e�����qdI�4^\Nؤ5r���H%*N5�h���Ρ��uK�;� dɸ�2au&e:���!�:$�Lx��d��䌩~&���|>us�~�S1����7�����U���A�������+��w�}�Ʌ5��@���P\&�����kg�G�\���e�h3L>�|҅�Ϥ���k�D8�b�6���#�Ω�z�ѻD@g2L�U�kT�q�M�s�5���H�{�4�~�5�dX����ܘi��݀��S�����z���?��w�������Y��T�"%��D<�k���>�|��_�u:�1��y2�8ஐ������d~p�Xw�P{I�2>p6-�8z��9�|:�%J��Ȥs�Ӂ|jf
c*�2�}�s8t�����<4f��,�Zve��q��<�l�� ���Ƥ���a���ۧ���{XY+���#݊2}(ء����O[�z�ו�Yb.f���un��
7��Vē�	Qv(;���C�}�S���.�ܾ�t��씺��� ]'ĉ��[C���1������i�9�.K?Iu��e �Q�n��x?�<�kJ���N]��e�́2�~��4;��[H�T �:����DD�P�b$�������O�����&���z<��O����b�ϗ�M���W�(�^:��3:2��l��D��k'��g�+��\��7��#9:������<��S�E�JGv���O�jI�s-���Uw-d��TTh��
߁*�(�P���p�x����^�w�t�w�@��uf��k���:�w��0^P�'��BՊ4l�fG�A�V/�NI|W&��,R1�PɅ�"G	�w�ի��LN��O?��Ԕ���B�]H[r.6�-r�3�g%�u�(�9��#(.-
)g��87��O��嵔�Qԕ���xԽ������2\I�l�Sr��^�%��>��s3��#$��@.��``V��Z-����u�P�{Ҍ�SCڽ,& M��Ȼ,�C!l۲�N�¦�Q�����hpB9J���GK�t���-����x46��;$ԃf�֙@�У�-%Y��J�ಸ��;DU+��5p�b�����C������W/�lP�E��Wm�v������!�r?�Q"t�q`
�¬YA-���ᛯ�g_��?����t A�ᡄ|eM/�������1=3�B>��`iy�SlyE#�_�ݻ���kg182����e����o ���/o��SS�������|�O��Z��wnbۦQ����ˋ_�ʵ�2�bB�ګgt�9L�w�w�k���}�^<�Y�?��wx29�h*Z������.&�$���G�Ci��
GK�6N1t�x�����И�),��%��
��G'3�*��R���C�� g=c�@��@/Z�:f�'����Bq�x{����,&���);��	���n�ڌ�;�g'�*�㓚����QK%Q)[����]?rYy(� ���H�@�TT�A���p�2�6^=yG�Dai��1:ԫ�1���%�<��U|{�?&)|�+>N�kK��v�5�;�X$�:g�Θ�3F	9���.!�2˲���PDɩ7+��N_ 0!���� v&q։r�F�������D(7"��{��G��V4%�2&������C�����M���>ų�eT����J�MV�V�w%���@��.A�?�mO��~�8��H3����ה�K%m�Ajz0nҶx�0q�8)�IGu4ճ�S�Č����ԍiHn��c��9�so��|���ذX[Y�8�r�hߔm�"ҋR]��ƅk������É�n�TV~v��3@ĿoCS�/g��.���fw2�T&#�Z�R��:R�L2��@R��o������!9q�(�~�,*�5ܽs[�L�(�ڌ��
N��L�Ϟ=�Ç�	�bM�(�,����h���+X^\T�?42,���{088�-�v��g �Z����z��K�җ
*ۑ�n`�'����c��DҐs�}�͚���w��ٹ9�Y�X���r�r$nT�Iۜ��k�x���ݯY���ۋ~t�3g�f&yRR5�T�\ұ:|�/��(�%(,���Z2o�>��U��]<'��<U�@q`:�z>6+V6����~��3k)���	�Pss5`��X�X�fq^HD�A�?���{��!z�q.	T�ߟݹ����_������+���B��F�Z��0��M[�N�Ta')��d���(���H]_uj�/�����yXRӽS�:CDe�Em�)�D�?�	�K4�7�q�����7ΌZlLڥn*�
��}0VU�t�=��E������Ҝm�oGۨ�j(5j(�(4�
e�Z	,-��Vd�`C���b2UF�^D*O��C[q5�Me ����D4m��X^X�@����k��P*�)(0��A֝�a���x��quIf�O���a��Fzu���.�PXU˖���6����pᴹ?���<i��y8 ����LPx]dp)�0�z��|��҅�T��bC��#(��k���|��ә����Ec庈轌axhH���:�k%!��lR�,���ص{/r�^<����o���g@;&�	r�׊E��=����*,b	�
4���er�j�9j�?ԅ�܈m�9~�s���ݟJ���� ��S���Z7Q|v�\B�P�-�����5��M��B�
��Q���1���)\��K�R1����v�%�Ζ������V��9Ο�Tj4T>����ʒԓ�v��G:�F6���ǙSg�e�V��"��?�`�Z .^���~��--���}��w��+gN������%��i�&��?�ͻw0=9���a�t�$v�܉�����L�=���~���x0��dNeSҡ�wg^�L��B��q��5|0�$KN����p�+��s����li,ۀc<��}���2t:�6.�s\����`�b��̴��c��C�/re.����h#��cz~	�k%���7���bn�:l^�ә�9�jE1hX�Q٪T˒�c|`�%�|W:-W����_��T���a�=}�����j	��p/*��r�)&�ΰ�aq�P.�3_;wv����W���Oе����QqJ �;|�bWy]i��?d�w�i'��Z���?�l���g���>��g���J������G�IfO�V����lU1L
�8�obl||���/���!K���I��ĩ�w-�����N0I�q�'���+�K�c�\o�,/�� ܠy^���<�����F�&������'���+c8��s_�,E2�Ub��, H�bGzX,��^Ji؃d<���i��k�|�ZY.�5� ��F����M����h=~���1�Ɵ!��#��K���*�kW�����^⒜�b^�e���L � �{�>%�(
�2"���nq=���*��9/祜כ-tg�8��I�}�4������>��N�&��I8<�@T��|�P���gp��5�mv�)<��X��í�7�?IA�4*����7m����i�V\�q[]�|� T��, ;t�fG������a'���QD���P,�9ZKx=�R���}�j�i ��j����x�����{����Ʊ 	��P�E:�f�>�LV��u�<��R��S@��!z>W�IΘ��_��� �^�8�)M�������Y�ם��-bWB�B܄3d�%PӷhI�f�ߨ~\Òu}������,~��jk�Q�Wן������f���oWJ��r��LZ�$�	<�ќڍ�xH�Vrj��S���^���9S�&�V��(*mS�[�@pU�:5� ���� 7����K�Ӊ������];�h"nH+�B�q�%���1�`⇵T�'��e��mk���n��h�қ��/X^��ъH�Q(@����h���3�',�D�אm��Hf�j�*���p�˯�_����%t���d.�];��ء��::��{wp��טx�P|wZ5�zSϕ��6 ����`~��Z��}��[P�I˅�N��8�c!��f39��Z��0q��d�|��1�L�=�K8:t���(BtP�!V�95 l�3K$J��;3� ��r����Xtt�18<��;w�ȱ�180���%\�rw�>�2�>~�Հ��������`c�d�����
�s�A�Z���������~p֮�m���ׁ����7 �>h&C3��Ȋ�H���KG����z���܇��6��R��������7��@g��l߱U���w0�iX
	<�w�ܣ"bvf^��DWO��lW7�]�RZ-Tq��U|��EL-,J!����+�L~��c�tc��MX����� 35&o�LV���W.�b��޷�y�����gR�{>)���õ�e�E��蛿����C�F��������}��Ȥ�+Xb�B���}�LT��W  ��$�(ゔ��d���o֑ND�o��O��kkE��/"K ��£�I<�]@��p)gHx8j 9�dȏT�$��$��������Æ� ��Ă�C��y���^�HE�(U�r�&j[g�j!��(�?�g�dh����/�ji�D�L���������5k�LޙD�N��y���;��K���9��,i��ҹ��A�N2�+�֓���%��;�� st��{L�MHU��bbrQ]�?��&��i�"��b�b=���~L
��	<c�G�	��Sp��sJ��u��bG�c]�\���5��s�Y�ho/�ۅSǎI��^,Jt�L��X[]�ēǸ��
+h8�%U�TP�#�&��q�)��D)�l�H�{�Y<S�ر)�tFT8a�\�5�=g��y�#�y65�d�듋����Q]���Ax�4���$Z)���<b��a�>�y^~�4v�ۏv8,��t&�h��e��,�.�trR����+�1ޝ>�&�M��>�[{$���q�yL%�����36�3??�'c�,�֪B���ރM�6������o�ڴo�>$�iܼuK3J39`�c�?q�V���h��J�@r�T�<��]fR1$SD�	Q�B�9;E<���
?�E��(�P)3m��J���B��g<B.ޙ%)���(̝���\��Ƚ�g�P(��<��h�ys^/�le��:b�	�����l���Tj�����K�Zn���:���ήb'���	B;�J�z�эj�Ium���������O&�q��O?���b��[�`�	|�Nn{����oA*ѫW6�2\ ���	]Kn�&F5��n4+e%<n*]àܔ���n�
'�&�@�|�OC
N�'���6�š�	bӭ{�I�l���2�W�i��QD)��9��~j&m�QdV��fMC���7�֞���^�Q,��$��PN��g䵛~(%�hW��6-�0� ��y�J��uue	�������\)"�An�Q���Q�ٽ����{>�+�\����`tg3Jޫ��*��	�u��\L���Q6�b���rjn��{�*Q�F<��;�9P+~�kK��\[k�ӊ�+C��U�'�b�������P/�ȹ����I::�/ US� �:�ͣT����;0�g��XX^�pi4Z�O����?������WXXXB�\��Q,^�h�l�&2(��%��#�O���Iş��?�Ld�ݘ��ͯ�(����~p�%��"���Vx��33�tY�QA����|o�8�7^:��_}&��t�=#r�07�+�f������ؿ��\W��8r�n߾���q����r��D���2!Ig���A��F*����p��]LLM��[,���x��	�M=����nڄJ��B��|6�\&+yҫW���Ͽ��I����ع� n=Ç翐�<�ߧ��mL܃�Fp���\!%%�u����
��j3� (�"$Z��cM��Z�:�(�HC�45�㢋T
;���`o��TAb���4��#���so����n����ރ�_+��G���0�E��Q���8MD��>�k�x\q�Oʎ����1ű�ʚΎ�#3�FC�u;wnW'l���KW�`~eYC�&P��Lg�TEymE	|w2����Ƀ�E�Fi�D3��Z�<�g��j�M	,��HڎT)~X�z�����߯`7����n���s�}���x�~�۪�s�E��������Zw���XI��$M w:��!�J��Y����⋋�QmF;��J��5�HF�C�D��ɗ�Z\5	I��hB�ZO�u��x����%�:���L�H	���BMD�ut�8y� ^:vX3Z�o�����P��E����"�Bִ�Z���4��Qm(�'�&���J���g"��M�M�ɖ�fy��2�fFD�}7�������)�CD��i��)��b�f6Ha1�M�B�%$�N�	dDH���
�D�.	V�n�*b&�����]��?����cO��٤t�eX�يvl߮ě�w��rMOd�b�X���4$ݷg/z�rJ��ff����3���ã�)�ś'b�����|:�L�\QE-�SS~hx�L�˔�&������J��Xu�9v�S�O4���+Ϝ0���y�q����\@�=���s���3s��巖0G��Q���_����_���K�8R��}=޳�C/�2c����o�������f��ֹd�k���oH��A��8�1C�}�fK�`�7UQm&�~>��6�vJ��Ve�בv���7_�n���|0���ǟ��l��/֪��j�	"�Z�CCڌtfPֻ���V3n�:6�DK�9g����x�����a� TJQp��U_"��4�L/��ߗ"�S�E]b��d�k��������4]�B1���p�H<o�N�#2�Xf�{�o�D�QJ��C�*L�v�r]L\���͒��$�|/�-#�@>�w��b��d�>�"zQX[���4�J��D�Gn]/�י�;��3�ډ7.]���c/%�!�kfN�Q�2�)B�j�6���OO_a@e�Az�4���g5�@�w��6��jp�'�:��J�{-[�u�ܥjIf"kD��yieE�q&� ��#Ǿ� oR�������CmD��7�t�=����D&�r����Q:t�A6׃Ǐ�5�?����K��s�=��Z��S�Ϊ`cׅ�����lgh�������ۃZ��h��F�M��la�{�{=:��:�k��VXp�[5!�#�4^;q��<��_|�t,�[Gd��Aj���͠T�=� ��zp��=|����v��vK�����%N�yYm�;w����W���'�6۶���o�)����IJ����o�dWo�ƥk��3�L�����'�)�����ght��?���$�zz�4QՇݩ/����Uu
�<��а���ե����!�*U%�<h�%
 ���ƃ��@��Nzuc��O/'�%d���ٍ�S:��|	<�d"���I�������,ܩh1؝WK�]+��+�wΞE�+�եU�=~��c㘜]@�\ECn�N�f-�zE���X�BI��J��L�H�I���oD2)�K>/��DI���۷G��[��Ju���ã�qI��0P�mTV��\L2��OÉC�d-�y�}]�rqq���173���d�fuqx��?�n}`͆��y�C��b|L��>1���}v��	��	Cs�;���>׆G��L�q��a�,$sP�N�pl,�٥5�ï>����H�
Qʔe����k/����~���5�n#S��S�wZ�n��?�����%���xi��8HmV0Л��pp�vt���z�+\�xO�C���)���5�J32�pu�"熨
V3�v�ف���i�T3�cJVf���(Gu�[�p$i�|,sk�΁t^�	bb�AZ�D�
��yՆg|"��9�S,�R7�ǎ��ĭg�w�>�_;�sNg�D�$�$B't�б�lݎ݇"�?��Ղ��)�H�s-����B�����V�G�zKCj0,\�Vh���O��Կ'�W"���m)�����JkE��Q���0j�9)Sj�R�u��t�H\ ��F4��5��0%���PZEOw���^�(�\[jn����ZT�R����0�f^�xӕI�[C�Lr�y_	8O,L���MQ�\j�y�`M���g`�p    IDAT����H����[!�l5�>�ܳS�s���;����ys���}elN���J��[���ܙ<X,���w�f4/㞀�_�%T��Wү��ʿ����ׂ�ԷrK�?���b�_���z�|�6B3G 0@Ͽ�Sғ� 5�@��0�tzƦ^�d������`OG> I�`BbT��� 0;�W����B��F��)eo�4����D��̤ٺ�f�k=����lՔU�T/gY�զ,ܫ�ܙ���j�f@I�#��|\���%��E�[��[�&'%}X�1y����~��%�?~$�X�4����h�E}���n,�����[��G�R��(ۋ�m'uF|-��S��=�Щ��`1EZ�3Q��E_��]�m��$�R��eM�P�5�3�n0)ON�3�� �S�[3D�P=�N�ҡ)�~��<�a�%+�]ŷ�M��3�Ɵ'�Y%�T�sK��s�R�]s2����-ضc78��>��O���_��D���Ro
� :F5�J�$30��N;Z�$��]��brn;k/@�	"��i|�a�<}�G0�� }����WQ�8hVП��������øp�Ct�Sرe
K���tJ�`�0�v�B:��Ns%*0a��������'��>|�o�yN{�h}oO������?�}��{��O�p��5|}�:J�:����O~�I����`��s������kWq��t�z��>�V�J+~rr���}����1���;c�q��ML�/�����Pæ����^���R����{0�����P������玂�%�>E�;�0��ٖ���5]۾��Zi+��˥5oo7p`�.�ٺYv�-�/.���I<���Z��EDR��$�x�L��7��S�t�}g���ݗP(�����݃��,��(Y`�}�}�vuY6o�+��~�{<�xj�-@'6�Pl+-�h�5�I��о�h�W02؅�����N�:5���rydR)Ad�ɸX����`��E��	a�&��k��g�ω�~�G�΋kɛ�N���|���KӊGO@HI-�g��"����j?����t�.�4��d|��$�='�z�K%�
��85�`o����=[��,t1Հ'j��[6�l�{�@2������KGe9~��eܸt�����Y�X���\�lR�6ϤF�����/s(fT�t��"W�
͘6��� �74�G���C�|FT$�<���閉�n	<:��n�fW�g$5�p���* ��*�-����?��lcI�����:N �H#F)�(��<�6a���;<�j����n���S=>Y|�d0��jb�LeQF�QU'�B!<W�+I���td�Xv�4�r���d���t~��a
�?�u��08���>� `"No&���T�ɥ��ާȁ�[��Es���z�n�O��k��/E�E��������n����w��3[��8wMOI�@	3��:
�BGNҹ���;C4�ca��ۉ+��w���[GA�C1n5u�#�K0�|�|.S�z���s�?��y�Y������V/�����P����W�.���J�?��_N�]nD���o7�2�	|*; Q~�D�a��T6ߌ5?, �r�s^M�"���!ƛb6�>�6�ܠ�[���ڂ�K���9�}������n����ȑ�s��p�C�a�ި��&�ٺ�7�F%��K�3ZKF6n�6���%f�y��47!��W@�UW}���!��>4�z����Vq��M�Ur�֐����k�V���i<�����T�R���o����t�"I�_��qU�D���b���;/�u��Q:p��Ŧ��jR���ӂu�Mv��~]�:ۉNk^m&�ę�}�f�G,$m�k���f��h<UNn޼���q%{�"wrvD�d̔H鞙ޯ$ﶨ∕�`Rm�T���@����Xi&K��%μ�6ܝ��q��M<{>�:Ո�qq����傞����?��6��?�Sm�-�	@���̀T�Ɵs}��t�����<�ז`���>Ձ���N��\0�%�p���I�q�$>���"-�|�(�+˸~�q����{p��1d��p_Ƶ�ה�S����tC=|���L:�]:�Y��}��9�`umӓυT����7�o.����@����'S���~���Obaa��ܺ���!nܽ��72<���~�]X[ZV�g�N%��1�^\­{�1��dn��!�u	���y��ڐ��{�N7$�8�8m�H3[�:��-~�~(���&��(\�:��2Ia+|jvi�9��װ���d���M�d�ұCjGS~���T�B�!�N�Y�m�c���G4��p]�R�����T�	�їˠ'�G�^A:��ja�+�B�3��!w������=�kN�y��Y�{�V�%�xԁgOzN�<���2�6�|�$��Eyu��{%�8�ׅ��2&�>������Q�k׹ �H���%�0���١�/A��{̟)�p���ϭu-}����l9kա��Ժ,���Z��6��I�s���A��R��_��C|��e)�E3y)���G_Oo��|�!��5��qP�	�
&��o�"B趎7��l��$��Z�u�����]�Y�0��ph�N9I޼r_�9g�P\ZR�e�4�|Z�7�ⲱPț������yM�%����d�x��{�
�a� ��:kN�7�:ϖع,��|L���?�̐��x�xEe6F��s(�J&�]L_ؙ��F��*�Mq�-�b>';��tN^���T1�������86oݡN�k��t♞/!��zN>T�F������&W�o�}��o�� Dԫf�'�r'�A���܌g2�S�(ٌ��M҅������ ��"L�3V8E�V��~�sIt"Σ�8(�]�tx��k��{#��ZE���l�pl�]ش��hw��l&�p��L�$]�΂YhTҼ&ׅ 7'�����&��7�)�A��Yu{�J�
uHT¨������ϙKp�(��l��A���s��T�#���Z(�ʒ�	<j�R�]{?����?��ʟL���W�|���̖�]�ED�i�ZJ�J08�/>��E��KB�����'�eq�.���>lӵL���ڰF�`����[|�	I���J�C�-�'SՕ�kk;a~���Q��UD�j��fDe�`�*�q|{��y�>��؆���'J��nEd���v*a�LD���J�)G�f3$u�J�l	�YP��'�L�����PY]ƭ�W�l�)w2u��&X���ؽ���~�v��|&��s�e�e�u�J�� �j�]Қ���L�z��g��޽����];�u�6�2I%��Q��(�Y�0,�-��<�phN�)��8�d�^��X9e�Yg�a-R<&����$$���Ç���[YZ6=X���w)�QИ)�m�J��{i�fڡ�&��S:F'��$�~��q8p@4 �3�{:.nZ8�A��P�Q\[��ג��(x�����;�<L�69C
�\n�����y�=&��a����m��ş{䂯M�c��L,�v���L�=�����߾�-�}����<�������>;v�=�z�
>����W�hQ�X,�0$���������9l�2��G�4t�008�=�������/�Z���#�L�?�	��<���Ӹ��7*�̭T+�Y�d%]�H�Sҟ��B(
ȱ��I[�+��5顗ju�b�Nf�wH�BL�jம?p��9�a�H�b�����~����˂!���un��>��"�ӅH8!��PI�߆����6r��:=	H{ںi [G��87-���ܵ�[v��o.����^��8�r�׆��$5��vC�]�Jg1?7��\F�i<l4d��e�6� �jM�O�:s>���#�G	�6���QuV�cl7jrbM�x��سc��9��>��>�&������Y�h	0�QɁ�/Q��2�H+�:�?��+��w� g�0��Wb�v	_g���@�D��M����}�@&��C�(q������U�0+z�b)�(�����G��{��+D�9������OIK�>��G�}��֊)���S������tz���w�2�zQ������0A��gbܿǏ���ͫ�p��ט~�T�¤^ѳ & +�T�t��
B�[�M+�;.�!KT�a2k��]�����������c҃�TƸˢ2S��.�(��Pp	�O3B��\Z[U?5��Ϟ���s9KO�?�z���r�%M6,z�|��H/3Q���{8_B

v��P���|�V4��-[���cvqET���Y�*e)�i��11&�3d��5�u��{��qX�x�*"�������R�P�_�׻�<o��؝�kr���[vHy-��k1^�%ˀ��BI�,���s�u��&J��RtN�4�i�Gg"�@�~'Ԩ�z[Ld�&�DR��N�mi�#�ᩉ����VX��%�]G�s&4�c^W'5�΁�f;����!X�����ß����i�Ԥ1R�
:=�ޣ�E���d�����ե0�1ʔ�Tw2���n*&�M"��X���L��o�:��O'�D��飏�f����b-�W��P�؍��"g&��LblPEÍ�)��델 !�G���"�VP��Z.��D7�2�4/Z�@_����xo��y�>����ȈU�T/�.&��<{�&+^����am<.V��]���Tp`�ݘ�<��Lϝ�Ya@���4\�����AH��U�����<iu����p���~6�L2���,vnA.����3<��S�ě�e���d��ʮ���b�q��1�uk�0��ѣGe�u�6�fRk��J�QkjVM�����V�g���U�D������x�|r��Uй�>�t��z�9���<Dq��s����[J9���
�̸֙.
�ZF*r�9 T�����U��$�VB*�5��-G@���#Gp����L<�/JK��>u��c��0'��ע�c��~�k�'ؖ��>x���]�R�0��D�	Pa�	�K�}��=��$����fK:(`���g;�N ܪ�+�;o�����a����c���m�$�͘����#����lj�}�	��t�֊j�2�#݃0Q.�y s]����h���0���9����4l��ф�[�#�����/��3���*��L��׊1�U��!���p"y�lJk��|<v�(�H
��n��w;m^_ �Sh�g�׬'��$p��r0�7d��>s��4�8]�r���g�9u��-0��u4QqK		[�!��Q�+B@�zЮ�Q-5Lj�?��;w�:���O]���Ύg:Hב�g�&enL�8�>?;#*�uz:p������B]�əiovx;Z[��B���P�zC3BL�%m�hjP�^ZC�]S�w����8�o;{�2bL�UJ���$�R��<ׯ�!^�������0Κ� Dk�*��ɪۗ�����v�:�οğR�hd��N�X~ϞN��;-!�N5i�|���LD���W�o���K<��E8���gr3���q��?x2�ߟ�s�EP��f7�<�MvF��u��]\Ǟ�B׫�	j���m"�|�r�l�0����=8����o_��+������h��&�j!�IK%�w��h�T��]�����Ƴ��@�1���L�v���k��H��!��y���+��P��G@�\z"$��k:��`�BCꭨ.~�5�eѿD{����Ǣ歭���M�R�q���N�{��ȡ7���(P���"�D,����Ц�x��ajf�y�Qb���[T[R�,��2��@v��q�����UV����Z��g׸/˚/��eŶ�7)���F#�[�30,z#]�57&�?����ZP�gW�3M�5�ko����x�؄�ǰ�}���Qb���:a�����C�3Q�9��e��" �,�Z��#�~���w�ހN"|~^�j4��0��!�]��������S�����?�<�7���Q�)�J�V�D��+���b=J�D&Ff���;���P�B�4�Z�k��)���'7��9�����R��R��W��ezT)֐M�k�>lټ�xF�B��EMטH������:GK.��(�D�"��L<�g��]zv��H���&�sI�P�H��O���y�M�ߔ���S���8�%��t��]��P.�ۑ�w��:�ifU�^�6���G����vCkq��y3��2���Z)���f������Oc�P7�l�,ԃ����cX��F�^�k� �77���q��li�EU�d$��FiP��>}F<wnLIh�l@���� j|t���=���>��E�L����^p5�:*�0�ɥՒ~koR�
��-�5�(����q��U\�t	�>���}K�C#Q��$�H�Ғ�Z��k�����\9�L�y~O�M�b�:�#G���OH�0��d_.c����X�h�M7K�4��l`��/� ���d��)0Z����j���=�u��{�w�!�!M�Vul���S�q�#����ͯ�I�#�G�WqS۔��Sc���c�5�y�f��wPmnRjn߽���g��49a�k�vl�:$���7�Y�F4ʡ�6�UR�(��BWo~��?Ñ�'0�l_sc��D��'�+�p�vȶ��t��WS	�=0;v>:aނ�G�ec?���k��`���[-֎r�����'�6PI
�)[)q2.���Art�\���:��{����id�zѡ�:CZ5Q�L��fFx�s��-r�m�zq�N���$�l!�8b'�bÁ��.�\���bID��D4Y�,V��Lʔ�8.�]{C%YK� ���KR�y땓�:�G����;6!�I��;�;wnHC�fU䓲[�āϣ���IӣwN�B���ޕ����D֑6��`��rQH����4�fH��\��N���qC���g��K�0[�Z��;$�C���c��}|��Op���0��32j��;���~o��6n�=ŧ�HF�q��^0��'�:?y��ɮKT�C��H`���I��J��r�V��&�x��	9�k+˸{�&n\��gO�(���qm�e<���dc�; ,��U�:7��\�Z����/=:���b	}�}���2�x�5��85��e-˓��`��C�r�&��(���_�ܟ9�������S����C1��Wi�Ks �b���6ZTxKe%���&��A��D*���-��w�Al۱K�˸|��q��4-%�F�'C�m0��,"(2�{�aV��pp��%Qd�����Zo��nXW�����}�T�����(�����l[�j�I���0�,v��A�>,�uT��q�Pn���v)���P�s�H�8�T��������<<+#��f��пh�,~l��SJ���p� ����vP�y�f�ؠ��������[,z*5�T+օb���*ˁ�,g4�*dY�P����4��f�p�tL�4�(D��B��e������#�t}�u�o����=[l�U�^�#�%Y�Z�M
c�ν(I#!����h���Mj�k7�M��N�?�����vJ�cyB�{�D�u�8���·��tR5��f 7/���"՚R�APw�4H�r�����T�4�C�=������L���u�&Rr}���`�ZI��d.�d���-�F��TG@)1�&��&Vg�q�§�6���"kcv�&��aq~M�spW� q��"��	egq���εU�ْ�ΙW��+�c�޽����8�ڐ���X[�j�9�*w_TI.J�Cb����,��$��t�2��&r�*���������������_KՄt��#:��GI��B�4٠	D�D��l؈N����D	mr?����у�:=~� 7�ܖ+)%�f歓���O$y�;d�w����P��e�Qv�:I�;i}���������������=b����B�D�&����G��[�c|����SVM�"�un ��< �@X���A����?�	F�F�����Τ���b^ӽ�v�\^���g��������I�Dl��؎�^?�m;wa|�9>BD��    IDAT��ܾ}Gj@m�a�{���j2��%��u!�����J��W^�X���������xB��	����p��������x� ��"D���KH��8�1��%�y��\�r��B�h�D7cj`s�n:�T�`�D��T�hZ�v���͍�j�3q�B ԝg��C�*LY�YB�d�I2�lq��x�
:~�0h��?X4T'$)���¢�E�S5J0�6*��x����G����<m��!�U���*�{{�?Ы;��!7�CO��[���߿G�t1��?h���`A�)�<�Z]2'H��x�F����{��<d?T���5��D#��4._�)����Y�9�D����k����o��׿�}�{�O.\���8��y���?�d�8�M�u5�L:�kAh�˭=9��T�h��%-�,"
a���ށSG��\X���q�����, F�W�3MRv���A2β3��m��<�b1�3�z��g����_���%�  I<s[Y:�j5P���ԟ^!�֬�b7��`��������{��՜��#Ǭ����3��<�#��������k�ƖYq�7X�q�>O �٭Le�MQ�-&d�g̡�G�?8�R���Wo`��D8�*s��螞^�j�vu)&��n�|H�� ��u�9�_��%ꮙ3���Ɂ��0����2L��(�aѺڡ�L�X0�x)J�6Sݫ5�H;)@�V/��g���o��[��0��"*�H��=u@"���Dֻ�~oO<�(!]9@����*����s��F�Z�o���ˤ�#�Ry�[��������Hr�2�b��*��HC��l�U���q��cR�*$��t%�ߓE��v���J�U���D�߿�������_C�}��f��� �_���_�@e.ۃ]�a�ރ(�R��<���"���Q�b˺��� ���>�(<�'�H��- �x�-۱m�׶L�"��a���E��4Ѭ0�O��,�
O�9���}��?��]�fA���K��qJ�^���1N��{�`��%�B��5d���c��-<�q]��X�����70�|B�HV��)au	C�95�CڵhYA39���c�,�>�� ���KU�خ\�iz��ԉ��J�C n����'��Ή��ZUk�DBDpm\'ou��A���������߫�L���+��w���7R5��LJ���'5D��$���1ESj�)���6�����ػo7Ν{SZ�D���]]^�$��xoa���]!�Dp7��u�/�W��_�v�#C?�a�(�w��a|]lY��k׫��J�ı��鏿��6�?���5�} ���"^o���s��"M�h;*�c��}C4�����7���v�ڊH��!)��96P&E/�ΚaO����a����uܺ� ���#)QUh�kEt+�~_��f�������w&�R�R��{e���Ν�!b���R�q����/�E�Q�g�r�@�!o�nx'���AځI��*�oX>�L`�h�Z禔E�{�C%���8rR;B��u�2�4���;U1(��n��C��f������)DMu���d��I����c�7ڬ"N�ہ�#=(�OI
������.�gzz�ؾu��I��A3�5o����7�7���yҾ�f������v�Yg��j����'��By��N��j�;�1&�`�x�46ɉo�D�8��|�᧘[YC,�G�T
����ŹsL���$�Skҋ�+����	_���+�t��\1j�� �J�tK
?D4�5�ۇ�����{ѪTp��E|��瘞|FkR���LR�ȥ�(�0)�L,���ﱈ�8iIň ������R��05����קZ�*����ιs������1����`���A ic�82�q�{�0QD�M<z�X&H�.^���S%v<';�,�qɮn<ibL��9�6���)u�X�C#��0v�ۃ��9|��(9���b�	L�O�>�[��^�uF�$�{��/��%�5�\oD��	�6�!v�ș�5��s��M	<{>-��B��
Q*!Q��I�C�	007���|�i?~+�d\p�1��gڋ��G���i7���X"�������y���v���O�;�,(/5�W�cS�#5I�7�e��wNc��
�5��Q1��k*߳���UR���S|
�:�~
�VX^?��
2I`�?�-����b�󠴺E���KG�������{}!|�!�����B�j�Ku�L���,�mߧ�3��fD����i<D�}_��h��2bg��^�%�VE�Z�b�Ѳ���\��h4iA�4j��[S�R�8/�����t��#��&���G���"W�mk� F��^"Z1�s-{�F&,"4����d�R}la���k[���m	��s?�ڨ#�B��'���ɝ��͢7��ģ��w[OXe"F�5�A��i,����E��64��et^{�^9}F�BnVޕ2'�+�n8a�/i��pĒ����~�嗕�D�6�&ǝͰڮK,���>��>���������?�X�<��4���6��J��9Ay�Q���{�qI�'<%�t�XXECwW?��4��p��y�4�(�cH�M[�\�n�ufB�*�A'`l��ń}co��/w���M��y�I��C�Kw.�=;���^Ew>#� r���.�T:ۡ�����t@D"�q�~��?H��e䐪e�h�p;uꔮc&�D(�F,A�	|;���	m*�Ҽ3Ӯ�n,�05=�����͕kXY-H�¢����H:J�s� ��xʚ7q�4%c,��]���0[��*��%���	���wtBt�&&���R�nm(�1)a��|xtV6h�F,���zy�ä�� X���C�w�מqs����Ig�L �&�cb3��!i<�LV')M�n�/B�����S,7B�*1v��I�]ʃ M:g����̱}��߅٧Q-,�ֵKƥn7�m��m��k�W	�%���@�O���X4 ��o��q��Y!�{�M�3$�����p�m*�m$�`jO��F$�煩��\�4�=���_O���ϫ��e|���x��c�PF<�GC��ԉ��}N	�+o�S���k�Y. ��~����������egkg�zkw��
Ϗ<�m���r�޿s���_}�	n߸��g��7O�c�-f�?I�x:}W+h�(�`h0i9L��Wĩ߲u+�����7�J���������}�M�O^�Y��8x����Z'3�]9�?��z�h�O����΢���F����4gjrR&uW.]�����,@x�]��f�̡�u)��X�p�0�Vǘ3*�̑�7o��#'0�y3<|�'�07?o�PD	�ɓ'��>y��c�4@Y��>���r�
}T�15t��\������br��7{����/�����嵢���D�%���"��cR�T0��n#o��~.�]������@�ߒZ���l�Qyyc��sՉ��k{�D�c=!՛{�I_�rt��u�K*������)��KǢ���5�Lv.�!���Uz�&y8G`>>����I���hU�ם��poav9�W����u�����������kq�{�x�n����_>_(���6�����5��Nc��=J����P�m-���j�l�ҡA<hٶ��ކO����^�O�_8Ib��fCH%�HtZ"2<��>�� /�P%�4-1�E�h�4CMMb�\���O�W"�r���	D�Y�8�
K�+L��>�`�K��FL����r�hU�N�u��mM�.�"-*5,c��-<�uY��|ϟ����q��Q�u4)M�T��Yb�����^q
�?*��y-�h�B^�����Y�0H�綈���CPU;=J���C���CY�/z��E�O�}ԣS����	�x���'�|SÉ*��؅y�L�oݼ���z�v0�!B* ۵t*��ۂL��T�p����`��ē�)o�;����g��Ь�Q�t����N�	&���i����B>�mD�7�׎�B@�.�;�J��]O�mș�̌L2��L
�7�hx�C4z-��6�K$T3)I�:VHC3�&��Z���w��� #ۑ�ȸ����m�VSJS���r���5s��3�i"��F�r�󋘞[Ԁ�\َ�r	�� Aފ�������3d
t�:!�s_}"��LDE�6�fcG-RtPA*�8�g��뱡���b �W�}�#���!^(QS�lg+��@��6;�\g���]��e����L�b���!�ˊVX#5���1~�@��R�_�k+C��iG��hB>qj��H�#]ZEo&���CW,�{�/�Ai��9�*��r)��6t���󖽩׽/&$,����<"�����ɞ�7A�����d~�������P/wl�m�����&���=r2w�4���>����,V�.������UyV$(�6;�c$*�ν�W���>���bz��xf�����:D�u��SJ���%s���h"���Ȟ�x����ܸtW.|���-&:�y�U%���$;|<7���	�O�����8~�N�~E ��Рb��"�*J�)_k�֐X_�i�u<�=7��޳G�7��`AƟyJ�O�}����`����A�b]guu<й@�[��,9�却�4K��I 4�Q����t�dF	`"�����c�e�t��]u6�'�A^&�\�ׯ_��{wt�k���3*�����,T*(�Z�D�G�뚦SB����^�y�{(T�����J���U
@�"|?�X�^W���ۏx:k(�W�Q�
^y7����lH�-m��G�}�}��`_����{����V�Sf$2�5,���F�,�q>�T�NR�Tt��F=VIS�XB` �8�إ��ސB��Q�6�7�Z�`����b#7Ь#�mz@Đb2m��'�M�����p�x_�ks�v���r�/���O&�����̧�~�?L.��ǥRi�T䐇y�Ҹ�	<)4�dUr[���6�D�	��Ni��%�ޠ�S=��r}*����H�e2?3��7*�ĭ./�yi�1i�Dg�����"�Mm�$�)�I�)d�,~�&�I��e��+�z���w!o���x
�^�\@8FZO��"0�C��S���=r��׽�Vy	p��WRl��F0��VfQ)��LB��6�,� �S�a������w�F6k�!ei�w��$�=�Ɛ!
��|�T��.�mex5��]H7p��T$_�Z�f����W��V�S�՛op��r;�%q��_f�,$�w���ݒ���!i]�2�xz"�"ǃ��O�w�E�\�g���YKx�c��`��T7�-���m�d׺`�E<�4�_�?/R�^H7�bRm�>�^�r-V�"��n�Ku�*�����>p<v^��I����C�5(E
 ��wמ`b�V$���s��ʒ�$*��&�ۖ�1+
�^�޵a�r�ңIC߫F/QQ�xKL���U����`2f��y-�gx�8H�m8�3�H��U��ڷ�};ip��s0Y�u���k#G��S��v��5j�ߜ��C�4c:�]�tL�No���ɜƷw�̀PLvu}�kP�f��2��]�42�]��St�PO0��(v^TXh@��:�L
��3����y��]G�\��z������CՊ���g���Ӕ��k����;�5s�,:��ׁVGIJ�Y���}֞�l��9�c"�iTg��,0Юu	:�p!�=�����"S�ž~!��\�2���v��E�6��:��A��ٹLM���"��c�VE�\A�RCww�}�������x���UT��$�FC�n�zx���ס3�z�u�F����@�@OΞ~;�l������~�鉧(�,�@ԗ{��	a��V�����"��� �!�'T�x뭳J�w��cZ�x�mȒ������\iΈמ���3ub\P�$�_l�����甗G-5��uIJ~��jчU բT(��ㇸu㦼0�}T�����M#$v&D��	�x2������l��L���GO��]{��ʵ��u�؁���͛��间Ǯ_��������%�-�s��\gT���4���V�V()	��a$J�?�kDU�b٨I�^}�b��̼$}c�a����"J��-�@f�K@��;TX��B��K��I൏I{��B�y:�����/=��5E�*,/��<�ra	�S�P.�����x�hPI��^t����w E�2�n)��jX]+J)��b��K���P��X��
i��q�P]�(����M#*
M���l��ԕj��SG�=��	�//N�߿���Z�����+�E���e$E�ٵ���x&B�XLT�@�̜=�$�������^�������RA@2��8%LBr��
Ԫ^���"V�_���ɮ�<��)��
@W����lR���ю4���qBZ�F��?�+�D(��V;ZI�H��l�e;4<
ޖ��y��F���E�h�"H �U�^�{�9��_�&�\�T<�b���0�8Y�&c)����;��L�MLk9�J�q��Pf�wh���8�iM���9�M��+<h[�~-�`[�/u*P�� x��6�wX5*@5���wq���{�[GvmA�3^��m���������q�S[x����	ҩA'S�E�I�d<.����<�l�q1�e�6�mSw����eݍ+�ܶ���f1w��W�_��B̀x��Z�������v*�O��H�x�?���>�ܿ'f��G�H���~M��N��I�06�Hdح>qxx�~�7�qk��ݸ�al��,p�>��tc�7mkd��w�%�"F~�?�a:5/~����
M���n3!*~��s�C�je �I��L�p�7u^?^_���!h֗Z���fwL�����K�aH�en�#��k`�J��k�A��?ܱ��I��DU�bz�'��8O���=<���/�`n�:�2G�dm\u ������] � xӖUB��8��w�'0�y�����^�|ޑ��+�t��Óa�������{	fL�'��f,� f��8�N�ӭnk��f�	t˯�D�4`P��*�G4�`�~�!SP�2T�9(�_�׆ּ�H��m��0���3�J��[X/!����=��xv\��hЃlf�H]]��T�3b>wv��fy��Gώ	4�'����`s�2�n&����- $]�)��:Q�S����s� P �ì[��}�y�#b����h��sw���A��YD���P�ձ��c#[D2فK���W�x�'f����m���)sBg�K����6��JĴ/��� �zC=���MEB�y�����X_�G$�C��4Q��ZX)xs�B|^5���\8z�0.^��cǎ�,��rz��L��5cgn�A"M`�'n�_��i��;$[�p;����=[�L�s�vy�<�e~��M�P�pX�*��h��7��,ɩ�֭q���i��I D8�5(��)�!cG2���xB'|��'�^��}�q��C�,������>�k��޾�B>��ΞB*A�AL�<�@��������6iI)c<�H<������Y__�����g����/���<�����̮ �|�fHX�Z�qx���0=X
IR�79[��_��=�&m��~���-k�*���k{�wz��֜��El-Q&�B��*5��3�X[���⌬���ו���W�4(�,W@Z.��2�GW_v�܋���ط�0v���,�lԱ���j�ʬ�d!��c�Y/��J!3�q���J��7���2f'��[�*������=�~��'�n��|+�<��Z[��J�!��w{���x�r�� �i�Xdg��Y�?�x���jw�
�m���)�,�IwF�N'2��_i���9AM���i��i #�Չ��A��E�����+�
�AP���TjD�ŷ^��7�R`ԺXP~Ш�H�07��a��Q��j�K�F�B+�Ja���rx6~W?�)�u�*�*h��2̻a�x���d88�x�;wH�a"��9 ���rᢴ* ԋ�p��Ct���v5���f�������ޛ�T�^��-7
kf����˲R>���wb��Z���    IDAT�㷥��{ 5���G�6g������2�vi5jZc��ﾺ�.��k��B��O�>����]�����]�����6�h��lpۯ�m�l����r�3�8��aV2�V3��}��o�:��xU��ۙ��@ш�gx�*������ 5@ʿ�@�L'��,�bnq���	�Ԇ�_�E`G:)�&z���AiL�RXV�N��s��SJr6
�.��� �PTpb���1�$r�����Y���r+�M�[�������j����� �@�#yA-�ۑ�8����R`����0�����J�� !)y:@���`.1�,��!F��f�$�3L���Jg�\6P�I9����bڻ��W���8	TY0�C�u��ng�[�Vf�!XP��NP+
�A,�Q�Hu�g�'��8�sG����ZD�Uƾ�.$��/�H6X�o�T,�v-ݑD__��m8Į�)-X��:K��mבg�p�0��8���ā{]�{����'���g��5�D��a��n�;;4l�k����lwŤ�:σ#�#�K��uE��8�cl�od�GSړ.�v	��O���X�̠���Y/>��vu�������"�x��W�6(�
:ne�I��������׸v�s�V��ׅ��.TJe�,-H?L �y�t��R�(@�����k��"�2�ܧ���v�Xt[IR%����mˮ�﷕�X	�v������l�}����	
���}>C�W��J��C�1�u|�.���1�gp��/A�՛C��Î�Zc	x�!�����?���Eܽ�@׆�^�_|���M���Su�����m�BW*�V�Q#d�X]]G�L/u��A�#�J#Kc#�D�Ҕ%�gO1;;����[��.2��N�+!�L�V�,���1ԍ��p��ɟ#	}��D�'���.����z ώ��W�uvj83o�uk��&�8�ѓ-%Uk.�\�5���S<~p����O�$����\<w
'�E<h_ZY��xvaQ���̂���f@WGg9��/����=�KX�d�g)gc��C�9@\�L�U��HL)}jՋ��c�`'��- _�/�ſID���������b��?������Q,��K��y�����}@ >��M�d;�<?���l9��f�`n4]h�����1�7:4P2Hҥ�� gȯ6qDH��|vC�"�KȮ-�R0m���� WTV=f �0~t��5P����/�P-a}s�t'N��О]��>M��C��B�'�?"�-�hnkct�B�!@��O8ā���Rt�=�����oX,-�x4ʈ�[�eWp��?�ͯ>D��A2Ԃ�ZԀ�a�����m�a͈{2��0�+ݹ ��~'�d7DU��Ι�R��Ѽ3P���^[Ԭ���o����b�ݛ�1n��eM���Ȧ��3*d���e���ں��W�����o;��M� �Ï?Vk���B���AG���[8p�,�Wׅ���D_�<~�\���*���� �tf�>�m�3��zk�zh���9��p�(r+���z������a-뛫nlA���0�ۍ�'�p��>�8K�aS�8lL�O�� !ޯŅ%|}�*n��W���n��)�;{Zsq'�P�f��pT@��>�1�<�Gci֒O�ç�����19�� �*U��x�F]G�Mi[�b��v���	nZ�O��M*@�dS�('g�Y�Y���1����M̫�P���\k�%a��q�G{��V��E� ���J��LKG���l/��~%*[ o���Ĵ-�ԙr�[e�j�GX�A�R�^���u�8Q�X�����x���LX�'�9"j�bY$Pb�� 	
�|γ�9O������&o�"��C5��8��DXԊY���HP�����n%p������CN~��>躺�&���t��ב��v�o�}v-Y�h;�V�c#�-�kjz�i�0y�
K��g���g���Ѻ/����lN��H�(�X�Eq��\|�5<����71���&��d���ɾw�L+��Gu����G�f�Lב:uX������M��ͷ/!����+���h2���Hg�eM�ò�4���B�bIr��'�hX�A���d^��m�H�H!�u9����-�,���<�'{?���~�vj�{���o�Z;g�%��u�7���.��L}ǀ���;�#c�@��ҍ뷤a�3�^�Iཀྵ�()n�Cymq)����t��I��?�'�'05;+��즟>}�#��q�2*�,��������e+]�l`x�����+,�T��яZӋ��ֲe,����/cuuU�شa�=8|�^��6��*ǒ�����'�?ޣ=����J]sIF��X�:�|v?4�S�B2��^��]�w��`6ڜ*B�L��q���	C"�%a�x8 9Xvm3Ә��Afeu�@��B<�57]�������a�l�č�lNA[|�s\�>���YI�Ɠ8y�<���߰�/bi#�J����\J��Y1��朤:��˳�,x_B*���KBi�Q-d��(�M,���������{��?~�ڟ/f+�1[���^�O��a���� �P�c�i�y����6�x
��m �ʓ�d�;d(T���9��<��m֐�\���$VW�Ѫ�U-�tz�]` Y6B	�1 	���1YvQ�6�Md�Z��C����8}�,��(ך��k�yc������(hP����x(p���&��I���!Of��A�o�i�y�� �=���7M{�QV�x5��?�����&��������M���(��Uz��=|�(>���.Ǖ�hה\�h��!�����͏������|�^�<�5�Di��s`I[�� ��dX�έP�_�ݠ�v���#�n =A���-mm&)�ᵧw;e/��"����˪��G���a�M;�i:թ�.Ҏ���8�DG7<z�O�8�C[ ^��!H�2��0!<����/���x>=�Y&7�f� ��텀M#d����q��A���Ev#��������2��ٱ����"'�{���v1u�l/ i6]v<N�8�=û���Y�k���ܼ��O��r�l�u4�H&������&~���q��]�LT'�����`�)M¢3�����`���A�`P2CX���P�ŤWE�IjfW�$�Xg�Ӱ�[��>��g�{pZ��yq�ĵi;q�M����eIf@ո��������f9�D;�i։�}���{B��W��9@ɚq��9\?���`D@�JC�s0U�z�^ZHr�����W΍xQ�6P�w���P�.��gl	�w <�H���	��Y�E��5�8���q�,q�����i�9%-[@�]��	7����x�î��_o?w`�%w2o{��H��˘Ӊ�`����@��9������,DYTqo_�l`#�32%vE����Cc8��EL�����7���_$*W��Z�$:(�3��VK�@$�a���P�5UE|o�Raf�s(l�cg��!8�~��5<yp�rh��.wex��n�����#��k�����RF���"��rY^�va�X:��ì�INh^{`Ցo��s��^j�������9�����Ld�a̸�Y��W��g]E��L0���������G���\�8_[������1�5�QDi��:�cbjZ�����Q1�Ǐ���ݾ�9�w�zGF�a��C<zxO3L�~��޿_��F��Ս<V7s�Ԭf�XͶ��W��Hrml�kO ��ʥ��i�_\D��hA����&�m�A����Ux��� �q%48�"v������� �̐0� x��=-=���;3/$>E��,�4�3k����Y�NN`ue�bAũ�YѬM2D��D���P��;��x,���sZ*�HLy<��[�ǟ~��}��:���Ŀ��;x����ͻ�Q����E��G�F"/�L��k�C�f/`Qͼ:�Ր�e�;���Ft�*d�|����������!�!���{��|a���F/�4\(�%4F���d[������f	�ͼ�4R�*3	�2�0}�h��jh�QG�~����Z9���g��x���i�;SQ�-$�>D��ww ��!J�y�U�i!+��RG�H9F�|Az�lnC�%'ΞV��J&����c#_G0щp�܄L�
o(�J�6n�f3���1lx�:�Sl���ꔞ�w3����%�=T6�p�a��'�3����r��,�R�򠆆�蠓���ѣ��vp���#qij[-��2�2:$�uW�5���6�C�F����e"��pl�h-e7`�l����:l�!e2~��Ҹ7_�9�洇�6L�P���#�i�\�{�,
7O{x���~�ׯ_�ד��LCAL܈���X�+��X��#Ǔط'ϼ$���=�y��l�.^|��N[�m �j�����Pq�-P�}�3��8I�e�Vh�v����Û,�ewg�N��k�+E��+���D�\t@�ɂ�s�y�iQ�5��n���Z0:Ѫ��v!3l�_'�+7��˄6H/�:N��Bo/��<�Ξ^|������_J��4C�g������,`Ⱛ|MJd�9`�`�v?��AF�PT�)-ޘ�Hf�2�<2-q��.s�Yyw9[p����ζ�-������\&{Epk�y�H8qu�����5�W3�o�QB��d,J<v�d�=�[X��n�����jp���� �q���'SL�����)��E,յ�(����>����Iiys�
��ױ��asC{�ַ}�m�8M�m |�Z��R���G���9x�t2�sx�Ń����hJ�0�(�r
�J����ص��R�����~���^�\[���1:vw����b�ZX���dRe�i��^@�=?���
r�<֪�^q`��cd�N�9�ɹ9\�uK����(��L��$�gW�W�[�@kؘE�ǋR�ȑ��2���4��>Bg<�ScG�y��	r�+�6Q��u�����{�8j�KZ,����W��[�s��#��^�.Yf�2�V�n�'�)Э,��n'�턆{�u�o��k�|�`p����xMڸ�up�q�X���(k,..*���X\Xn/��\`6��ӹ�X�"82v��ǰ���ə9ldrGb����ѣG�i����=,�L��#x�s(2�W.����x��w0�s7
�&g�1�H9h ��&7*Ȗ�^��l�P��W.4g/�G�P�}/��@0*s�|p�%�*39,�0D��5�)��m!g��w�+w��v��z�$�a�Uk���v�8?G|�஢����&�b��=l,-
[��4�#��ˀ	J�Mt&��5ԋsgO�#��x�/�% y�k��������UP(�8�Tq��kobxd?���"	�<�2R݃"�+� Jd���w�`����A�[A2�Į�4v	��n6Pͯ/�P��d�������};��7�lf��'�FS �?� ���{�F��	)lB�a{���>6�U ���� <Zc=gګmȴ��	4} ˳Ӹ}�k�.�!b�w�	$�-��ѕJ"��b���TAvQ��M�Ҵ��6e�ċ��[F�xH���F�:�V�T���S���-�}1t��B$ݏ,��=��|�-�V�c�����$[�aJP4hn�U�j�@���Y����CM��6�_��/?����MD}x�E�H���X�I�F����8x�,�-��dp����ֱ/
;5��P*����7 �,�6VN�k�f�+n��C���!�ey������ϲvsv���&i?g�L��T����U��\� `b7R�{�~���ؙ�\�������k�Xk��u���w?�BH��p��Q��x	OWo�ƍ�� �a���o��up9xH;ݖk�U ~;��̅��\�B��7�XT���5d�DN[;K�Tɶ��P�wF�ɧ��� �+�U���p�j���I�È�N��%�Ґ��ص %>���Ĥ�Crby�RDn3'`�C�d4�֐����p��\�~�}��2A|~�@/:;�%�^����� ƫR.���<Q�����g&����ӧ�J#��|F}<H}���{���\��;�1u�m��ΐ�îJz��P���	B�ư�� @3϶adف�l
����s��isXq���R"Q�?����ji�����+�e��خ�����g8�9L����sO9�܉���"�Z�t:�X��Ą�I�!��o(��L3XY�Hkߏ�Fr�ଣ��:���-d��V)+ ߪdAN���QN'��S��¡���]^+���v�-�䶵��L�*��Z7�o�AG_�^sv>bYa_�^S[(�abg9�z-���烃�-�1��B���U$��G�p��Y<���p}���N�E�#��&���4��5{��fafa��+��2��f���z1��!���#���u�4"�ٔ�,�h�g
%cf g�&YV*�K/�����w4�5��<�OkT'��x��yJ8bK��v�h�f�c�i;mn��-��/n�r���g��a���y�1W��u�L�oxv��e�ԓ��z+���>�o�3K�z*�B����P���c`pv��H'���}tv���ѣhՊbܩ�������.��������>��o���^��`��LcvaU�}�r��&��:6�W���D�X�7����(N�9�l>��%���'�g� ;��f��%�Za�u=�r��KݖA��2gVO�ӑ�m?��Ŗ���6�0�Μ��p:9u+�ۜTf-�XoH:�4�4�n_Cvyр�(� �!�ѐ��� ҩFG�`�@��wf���Oy	&Q��XZY��+�q���)O��L�X��a�}q�����W1z���>��l��1r)��:�<�}>�V�71ܟ®�(B�:­s1���D���7%4b��O?��ٍ�k�>�Ii�\�wf��B'��!8��k�����z�Ál� ބ��Y(IF8�Ʀb*F��=}psSO���t�0;�!��݇��=�=ԏ ��~	���kЯÈ��z���T��ꚆL��W�M_�d�1�<�"Ҽ�l��O���R�A�=�R3�5ƽ��Ƣ:��f��iSq�Q���R�,`5!�Q5U=uPN�Szr!��c�C	�(o�������b��ʳ�̟�6)+cJ�������$_��5����DL�ld7̐���&���QZRH���/�N4s��Y�P�=�f��Q��8��0���o� �>�9�Y�����X{ƖZ��Y��/�� �'�n������c��a�+W.���G�w8j�x�˻�R���{�������λ��ƛ��-9B�^ٍ�aD�1�AN��ɑҴC{��qw����~�:�^ $�����@��EK�!#�k��W�ѐNu��o�vgN�������X���m~�3�����M�����$�1`�m�R��مy�ڡx�̡Pa�G ��9�g�E� ��زT2`��/_�+����჏?A�X�����رc�V�g��S�|./.�u���!�W_zj�K����\ŝ��4�I�s�O��5�1��+�®�N�$;�@�d�h�s��d��\�95�J�3�[�!���K�l�5Է32��g��k������i�	Si�/SGf�׎6��d�x����d�-fv �ʥ������S�(��q#������Fqo����W�NA�;{Ķ�,�bau�RE�ƃk?0�8x���k�ZSk�\D=���f%�g8;;���8BA���x��3�N$��ݗ�E�{̯J�u �)��sh[w��v��2��5,���
ȭ�?K�[�C�I���ؑ��H�D��8	�ZӃ�7,��؉Sx���J(=ᢞ������LyjxZ��z�ku�Ǧ�/}=g�&>?��q��L={���?ɭ�#����$̍�2\&'����_�'>����N�~�p��';�>�ܟ���n;C�`�-؁r�f�-o�E�8���qr��b��>��w����X6�_�Y)�����}fiF��'�Ț3�/����獾�'p�}�����ͬ�*���'ŀ*?|�0�N��SKʇ��� �٫�6����ޤ�!|���p��1$�|��{�� �e}    IDAT�>v��w���عg��az~�B����5�+uln�a3���9�C�Fe5�+����b��P$���%����4嵡(�ɴ�v�t��d/�{�:<^g����J���3�d�����Wa4�f���Y���bJ���#+�T4���'x8~�J{�GЕ��3��@�d蛜��#����JF�ˬ������ �iM=z2��%��\����u,��K]���cfq������p��+�%��Y��ʧ���B��^��p��[��YF:�ľ�.�LE�u�r�^��:����S��^����L�_�|�/l��,S��U+�˖ �.4b��d4�6~�������>�6t���h�q3�J�C��������К*�� ����?�S��Ȑu�LD�~�w� N��î�m,��kr15����Í�JU�7(z�f3��8��ՕB:�r�
��k^<�X��_��b���O ٷ�*C�<j�s�a�M���-� �1[84GŖl�x=�7���lJf#�����Vk�lUP\���/?��ۗ�d�T�z���V�TF(ǎ�{���!�Q���ɔ�JJ�b����6���H4�d�R���
"�XL��tL�a���@K7�����ō�j�ۇ�=�����w���������`�C`iQ��{�Qnndu9��M��/7�rA�����~����ꥍ���5��7ZN�+-,ȕh��>��o��\P�ݺ��o�!��R��9�]��;��}�!3��i������K�`�>,e �*1{|��:��ji*��q���$�x�<N?���n`v�l��K�D7^[�k�6�e��*����|}=�سg��|r�B�DR,���8v�܉�;��ƴ���N�ٍ�ϟ ��ZE���e��|��e�;�Y�Vt#�cs3�(s��]�������S�;\z�U��u틋mp&W����?z�ŕ�P���c�lI	T<�KN��iVKh�JF�A;A,�[��u����9 �S��߹��[w�����BOa[��۳g�=���~I��������*?�taJ�8�J6��Ĥ4�l���Qe��Z�&T+��δ: da��� ��#?������X$��t\LxH�'��i��|�(6rE<���Z�`@�>c�*m��{�>A��)���/����Cys�rN�1m�")_G*�{�g�3D���ނb�~a׃��A��S�c���ۢ���@Q�M�)��(�ﾻpx��ۥ�uhN]�}?����V�!t5OH2�#ǎK�A��)j�i��/� ��^��N~�Ǣ����'"d��T���{���W/a~f������9�2���>Z*f��a<�5�BG���d0�|�mu�;�:#(���Q�o��[�MD��Ծ���#a�M*��ӵ��3�k�*g�Ѧd:30���^�b����OYƜ���~���0$�Y#��-ɜ�`�E):wJ�>z��$�x�ܻ�P��Nө3̵�3
H�\��h���I4|A����z�Uܾ~�KsHD�x�8Ǝ��];�4������C���7��;��8�O�`jaK��X�W��+I�N�;��5<c�9����#W()� W(K>��4p��A�C�T�~N����p��̀&�B���0 ^���^���k�RU{V�Wކ��"�5xN����s�,�����[W�0�a�SQ�"�=��C#�3�+�O�E���m�:���� �6w��_m��v��3���� ��6���3��.brv+�X���)�X=�w����9|XY&�Rk�<�<oD�j������C�("�:�����9���W������ ��?�|��?]�W�,S��U��C[+o�x���h��* ��Mn�\mJ�lo�%5Z����?�Y��7���M�eM�r��ߍ�=;p��vu��� L�rK�xlw�z�cd0�s6SD�@V��X-D�x��%��&�ϣIa�糫��O?Í���=�����u����D��]m�	�}��K� /�,�ظ7	x�n�m��M� ��*#�,#�<��>ē���V�����(���A��Юa$�iD�I����aTjm���f�&�,V"�y�Pȇ}�^�V���C����k����P[o��Y�\p��Ԧ��,څ���7W{X�?�H��)~z� �]ۊ&@�ϧ���Xr�ކ=�����5�aݸv] ��:һ;!VV7��S�6M������*��ʭq������8]ǅi�#c�ל�`�t�������s�_ķw���~ʂ��b%2�>�x�I�!�����K��D5ۼtw$����8q�ݽ�T,�����3��X-�@b� !ʒ*Ţ��ٍM�yD������Ҳ).�n�0n��txdT�.�T��Bj	����'�~���E]Ʊ�5P���C|��b�� 9|���� ���k%����޽{���(L��k��kzq~�sm}1�q�j���Aݑ1x�<��i�G�Գ'��o���T�ϟ`y~Vp�c�r�֎�H��0,z9{L M(,�2=3��Y����w0��	O���QQәJJ����_���&��Y��b�=�W������w���jU��ֶ����P����8������f�`�5�H&ȾǵG�L�p�U�c)�UL�.���,2�Ee�ˡH1$��:�m�X"OWk @浔C%�.	M�S���>5�0U$U��s�3���}X@�}}ؽ��=��fu{A`�%��2 ~k����5 �e��>,Sl�ň��7�WA�2]G���~�4}0&
���FR8ttL�����%9x@2��0���P�H3f
��J��}��U�d��ϕ��J� ���/����y���3�뫚���Z>�E�H��&y��α��B�]�o}�[�p���d�h:4����5�5Dnu�(��4���侮��s
#+�L΋��}�5#��J�}�.��g��e����sYDo{-I�y�X����r9�5v��>ͽ�v�011����19IS�%����2�8�@��.�8Qf�t!�H�ǰM���޺��(����gp��>��t���}��$m{�Bg�.L/l`bf��l*��["477�չ�\O  ���������l� ��Aj	�1N��1DW,Չ�Ǉb]ս!�8���v�\��s���6��݋�$�g��xui9/�tṟҶ�΅�R�W����4��<vt%��7�݃�8u� �F�KNC����qd�#�yA>�FIB@g���3T$*O((;H(�sqbj�s��{3�x>����UdJ5t�7���G� �D����f	�J�r(�އ��%t����ؙ�!�}����8�C����_�<40i��_�A ��O�x9[��l��O��V6.4�{F���/0�ifc2Iv���o���l��i57��L�4�>;���~�bfq�Ct��8~h##�1�ۉH��Rq���3
�`�J�A�V�>����T��OL�SH��b�`8Ɵ�C�o%_j��o��ϯ����v�ș����!�cI��*��{n�์�ׂ��ƒ�8��ۄ2�0|����&f��ru���y�U�Ed����ݽ�h�����f*rI�%�ص{����~Db	i޻{{�q��y�J�����9E,�dZ�4D��-%������l���X�����T>5�`�>���2��H���I�5����e�[���Z��YR�CP�����tv.B��d�(-���������{�=��.�������B��~�Mv�������JӋ��n����JZS���ג���YZVB�"��k��;ï�~�:-aL���Bu��9�?6���VZ��2mv��7
P倎׃�����o���Qܺ��O9��,�W��<pЉ״Z-��ι��ں�S8����u���
��d,�Ξ>��z�;����է.Q<�f��7p��u���?���
�
N�=�Ko������ϾP�.��sg�ʫ�����>�@�]ֶ���[;_o���H�PD.�U1��bbj�Obf~	�BE>��p��"�ϋ�$p��)����������q���&����n1T��p�7C�|�e�Iw#u��o�$�c�H ���'ж�0��Hģ��r��)�|�y�8 K$p��i��@m�۷���!�6}]]^7�@���++z���g��{������~I�E/�S�餀{���
|��c#}hy�X�����I<��G��{��%у���<��+k]h�u_��G&�Ln��&d�}-y5H�H�X�4D0�
�.ɥ�7��#$�ے����ݕ8�����m �޷��KS
� (w ���ra��۠,'���y���W����Й�Y�Ү�у*Dƈ�3_ �D>*0GV�ν{Қ;�'�����S�fqm��a�y��r�2i���¢:E�&�p��A�|�%�/,����}2�"�굲B�E�u���f}�=x�қx���10��h�����k"�T` �^J�l��}����0��s��5�,��a����L�����>��i����q��ϳ-[cS@:,��y����#U3(��]K�.�jZ_SS3x>1��p�+�|f8����IЂ�)�JˏP��}ع����V*���GX��@$��o�����%t�S�{��ed�@��9LRB��#W�a#_Vw��~o���a�X��bm}�ْh�(v:�e�����:��ʻ5�H�M����9S��M�P;R�-I�{��̏Y6�#�2��&���tͱ��Idߙ\�X��?��/;"^�%C8�g^>w��D�:�.H�,,ͣP�a�rI�F���}��-�U��s�.D,:y��d]���+7�tb������:6���^�é�04|�PR�����H���.InTA:��޾�t%j�j�Q̬�{[տ�L�˙c���Z ��O����/���F�?j��Z��Rg7�����>=�`(.ƚ�FNl�E h����F:)j\	[b��n)����T8���&���{w�öG؇dԇ�	�?}T�Ra����<6�WQ.����Ï��6�H��0�g�k�&�ǒ�D�+e�X���7��������F�}�n�~�J͏Rˏ���8�����GPl1�а��?����I!��gO��~ڍD`f���yн�I�.*�F!�����?ǝ˟b��-$<v ;^T�H[�A.����E�	������&�C�l5+<�aEB
(��߇t*!-2I�[���b��8TGo�vQ� x�.Y�	�{Q��f����F�>X���G}��|�5-E���e噞�AI��wkH	hc"��I�Cn��=�{�@��A_�TJ���1���-/v�;���w��ǋ�Wo���'�PsA��=��.[>��#�u],�F���+������&�:�{��@�1Y2�n�@:	���0�~���A2?� �z�D H�\��?��${ЛN⛗^ũ#�xz�6v����N��� ���ֵ�J���Q�Ihř��ē������U��Z���^��vc��������?:���ؿ�z?��O����R�.y�������}���%�ؿ��%�ml�G?�ґ�̰'��Ρ�ֻ����q�uv���0%�9�������5��6�q�M^oɢ�,z}8{b���op���������q 㯎�E���9�T-��5~X3�C�/�X!����Q���ӎg��!oK� 1%��:-Ἶ��ҹ�b�*�n߿�ɩ)��}�����A�,h(C�z㺺(쀜=u^�"�+�0_]_��'�%�  L�� ����t<�D<�h $֋�Z3�x��9fWVQm���%�`Tz]GRAʮ��mq�̱o�gDM ���zq�V:2xZ�r��}0E��N�n��A4F��[2��#�����kNҲ����_�n$?�1��Z���f�Q��o�IIb����q�0v�N��� ku��~�ב�luۅ��-nm��Asf~��T�s�N?u��m�����C������;��-�t
��"��3?P�/��J��&���~�><z����c'�����B^E\�����/m�����q���{��m\�pQ�5�|�֖״>I��ÜkT�mh+Q���v�I]C�k�,c֒ݷ5�ͽ�ɚrv2d��K����e����Ak[ę�+�C�n�i���F�}u�d�&+ryk������[������-u�$ݤ-w���5T���#��A4щ��!�9�f���Oaqn=	�z�4�w�^�#�c�a��-Ԛ<��ÃG���K�4�r��5�fvC�/H0�őcc�k	KK<3�$� *����`�b�a8�V �*X䄇ѢYy!t4�\�m:��Ҁ3�י�*wR�U@� 3�$��$H���w:eLr0�-oMY#�F_��#�<{���z�~���WN�ȁ=���hK��2x�������h%Q�=����"Z��v��U4B�R��G�l�������G���ML�,by3��bI����8t�v�=��7��b9�>N��r!ت�'������!D��������w��y���'�&���}������Ձj�PÇ|6�d�{��b��u��s�;�-ڣ9���� ����ń6�t��Ma"�!#�Z�
&=�Ӈ��(�%����`O����}�NG��6�lf-�P��`�� !����>O ������*v ]�=���D�G�����M\o�x:5��7�aa�VW~,��U�y����"��@�T��3\]jY�R'H���|2q<T0�T�<LԎw�[�52�MY�m,L`��O0�� ��Y@���?�S
؎�#��%��X4�d2�d<&�*��zCP�zgWZs]��]O!�����y/|�JY �=f6@[9+�&iղX��6l�'�X�y�=v�uKm�3�Ŗy��������e�m�EnV�q7�b��e��Z�
`��M�d�v����Ëϯ���t9i�e��2�˨s�P�m����i�[�n�h�ݭu~-:5�E	C"�`4��@�bh'�����i����P�a�����T��V�Is�kѢ*��dgǎaO7��c��>����-C��f0��{GS�^,@2��?�+�A�ϕ�Yn
>�<>�ܻ;��7H���V�5C��K3%\?7���?�ˏ�ljVSG���7��&�<{��?�R����s��~��hp��j��;d���;�����u�<|���U�tw���C�F"�q�.>���P^�τ�Ȓ��
>=v���[��6��g`v�)⑈�b	Ph���ݥ��lF����0��o�j�����C�H�b����}�	�9�B���z��8������!���E���}T$=����,>��#&�۾p��$L|}��d,���|�����ȕ�طgX�
�_��f��K���r��kbum=]��L&4�ÎD���ad
eL�-���	���M���V�I�~�	����hu�J��;�E�!��+�uIi�������(ĴԍG�����5��_c�z��x�fWs\ND����*�!���f�6���2���bJr��"��6�_f��Q���#�Ǻ	�S��S4p����0Ǧ>���ל���;Ã�&�w�b��i��w��"��?�w�����"~�;�b�� j,�4��u�Gv�df�����y��$>��3LNN�u�>���Y�콟�U/#�
�s������Ů�<�f7����9��k�u���j"x���$LT�����<�RG[�}=��u8(�^G#߱E���&C���s˨�\�ЕQ������;9����3���}=7��]/���Ņ�~a�J]�"v=��˗/�ٓǺf��.rև�m�C=a�BQD��G���A����;�e��xqh�n���e�H%��]���Q(�p��=��\��rÃ�݌j�R�T@ Ģۏ�ǎ��h3�!�Ud2̛�!N ���4�3t��(���Qi��o��F|e�ښzV(��b%���4��� =	�F]�3�Q��1��=�Ǿ��f�M�D��>sb-��_��C�j���;@�}g���3B��W�����G�+��g���5�yk��U�;�,<߫0B,7�5    IDAT�T,jd�h(s'���z�n?��~�=����&��W����c�0������_�'�B��X�
&�(�����}�۟�P:Q
�2��|�����H�/.����\�?gJ�~2𼈥B	;v���}G��ՏB�m4�����X>������<��|] ��H�a�ɩ�֖p��e,�M�# =@¿EG"�x��ѽ�x��i��ՋRv�(������3�z��t�;::t�	��C_\��Kk��dNDtú�i��ud39�5̭l`��3<|2�R�U��_ڔ����8v�%�v`��#�%<6`E�:cg���&0Nͱ���s�P5#	�;�?����BN�e2�F�����ՇX�x����F54+�Ģ�܉�]{�L��=ե�K���$�#�69��δ����J'��Sj;V�d/��W)���e�_`"����:V��/po��_~��������[}��PsKn�rx���v����粪&�Ρ?w.R^s�1�]�&/s�,N�����OP`dp�^�O�����"��� �BU�i�1[v(�ju�ߋ]�-s�NR�M�t�%n~�HH��d^��P.�߁Oz$3]	��jXm(72�y�sn��M*�=ht�|�u_�ϡ7�Ʊ��Н�cuvGG�b��A����:Z�2�����4��7̇X���\�K/"3�w�m��a}�=x��t"�ٵ2�h,��-���Xϧg�}��E��ǘ���[��~��elld4�I{�s�.�����?�䤑ИdV��L��ǎFOg�����c���bd�~���%;���o�Ͽ� &��ɽs��sW<M �&Z���~F�GfmU �k%�#_,�߼ֽ}݊���V�%� �L@���+V�ɓ'
Kv�(!�J��It�R�1Ћ��S���;wi�bm=�kv��q��8�٥���?B2����|��ba~W��,���������)�K*�x�]���t��xL_3v򄞡�?�w�c��O�<�[S���"�V�k�.,���$��Q� ���j�p�5a�mۮ[f.�d7>���׫x���|�I��ט�c�k���5۾�楽���:s�)7��W�Vj�e���V��(о���L�k��p��,0�~a�Q��R�n����}�b��`�%o�A[�|�����5��K���o��D�\h��-��g�����7�;㷱87�w����G�I�7�E��Sq��il�(VX����wp��5���?ssSS���I֚��� ���3g�J	�ټ��^{�5|��ߕ��?��ɼ���b� IݯZ]&����ﲡ����XX;G71c� >[3n�g;�n�$7@�k�ʦ�b	#�\�e��Nw�]p�[nC[l��ȯ��+w3�C y��WAPH���ؔ��իW��?�}d��.�#�by�@8�d�>��v��ȑcX_^ãwQ�n`׎>��B��@���="�8%r��;�+�p��}<z6a�<>1�˫+��3��& ?6v'� ?���L�áq�����
b]o��A�#>��'��ٍ�_�Y��~�	�T��t^J�Z�{Q,�\�89� �C�r�	j��@6�֢�9�-�
���>�g�B�����qt�n�����#x����a�9��뙍����������g���)�G�`���sO	�"GB�N�DF��ޞA��!LLn��O���1�h&�1����z��k8{�m�{���ձ^,�D}?�V��� �`*  ϰ�F��P)n�}4���n �����|���l;F���I��P�O�% �,,�4��[ O�%4��gۚ�	�d$�'����_�S��+�@<�Eg4�#��҅��Iauas�OP��
�9�>��y��R���������u��jn:d	)�HG�j��ך���z��L���<��:
�&2��?��w�������Ad��ó���9�x��<��K�����2"�H���T��6,��$I��J�V��6�	o�RN�)�Zzv M!O�#ݣ�2�� ��:��S1�tu����$�O���'�8͘M���M��+�P��*�զp ���ng��Z+>ˈ�g�qqIh,[�.�j��n�m� d+��?���m&���jEV^<\��i)Jk��YI���(���lq��܃���Jf���qxFL����<p��e̜�}��b#�ua��M[�̰�I0Em5�?d1�L��!'�1�L�<����]2~�6��Ƿ6�Ό��Ԋd�<hV*bYό���~�<y����p��~T��MM���[���
��;�ӑ�˯�`����3����ZE���9t{F�m�.�6�Y1��a�h��C���Ǉ�~.K.z��:��_����'q����xoΟ	/�����G} �����ԏ�B픒ģڮ,/�X,`��^��p{FF���������G���%y$΍�w��ʹU<t�i�m�BA�2�: �tʢ0����s8�g������E�����b��B�$�=��@(�F��]=�Hut�#���=����Һ���O>�{}���,:zz��������C���v���k��Oޗ�w4l�������F�� �P����7u�QS������"����ݙ�X̅`�k��inaQ䋫(s#����h�Ѥ-�@� K^�-x����b�Hh(��@ Og,��r�0�lM)���ؤxjn �0�"￑�x;*��b �G�D�萁���4_�#��Y[�;���C0f�{����S��ǟe�<���Z��� �w�Ǽ����azْ���������.4�?{>)�udd�޻���I�9q'��`c�\��̤��I���C�"I5?���_���{��C�Ξ���D���%r��a�s� ��Y�Xƛo���Q��3�$�����!��؎���-�X��Jg���c$B��,�<f�2����=x}mx�`��˖+�p�k�JďK�h���{,sn��sKq/��}�?�ߋ�߂�6�����f�{~v_~������̜�	��J툿|a�:zNv"�ի�������f����wa�`�"��M�x��hf!g�n޺�GO'�lyQ#0İY,arzZ�_r�
�p��	�8}�\	�+�dɖG���g��J�jf(M���� �rf3,�ӏ�#��V�]]���s�Ѡ�Ɣ�%��X"�dg�0��1<3������I�Nfof�Z�d��U"��V�p��l.������=Љ�cq`��F�R���D��ڷ� ����t�
L>W���|I_G�$,����a�@�����'�ڃ�P(�p��m|��U<z>���sx2=O,�C'.�W�E�������ȗ���3W$詵�����[��|�����p�//���T����������_��B��
��@��C�J��
�=��G�j�Q�@ˑ�x9����P��иxi�Af��]Q׮|���o"���3�������$4C}I�2+X\�B��}���/2�}� ���f��ժ**n�Ԏ
�L�w�)�����>~���E�m��ݬ�\�`-[T�����9~R��S��M ߶��� Բ��B�Ӑ�R�ayq�3&R������CHuu@���RڠnlM *����F2�8����"��Ri��;�������it����NE�۝B_w�:�b���4�,(LJ���y�2���{kK��. ρ@{�YɊ�@�>uۦi�*�N���l�ױ��{C�L|�h�M)�mP-0GK�����a��ρ��z���"j^�
@�~�e��ּ�܇��_���H������9�^b\ ^�yl�����G�L'dD��1�z�����Hl��CDE6��xj��Z$�&��4�C��U��c��Ά�� LG"��ƥ�.`��!\��S��řc��򘙞@�F��,��f�ܳ{':qY�fVVp�66�a�����BA��Q���C��[X�d�\(U�Ɉ�ک�GϞ���>��fF ���3���k�uM..����������c�e����J0}��U�P�]��e�a��.�ދ`,�/�\Õ�ױ�/�U�A%�x����WΜ�w�}��E9��X8y�zz$G`�jyqI�p�XM&$���XY�[�eD=젴L+�r�&�R�5x��8�D�K�5���,K����?�
7n݁/���/��3XX^�?~� �w�}�w�Ɲ�q�����FV�3, !K<�P������̂-�v�6��K=s�=�s!�I����П[��_^�DM�,2�~PШn"��V('c^�ƙR�j��:� ��[�!j�����;Y^z�{%� Kkviji[�r�$��+O>#�����9(l~nfj�t?Ʌ��20�W
mXk��Ēa:I�<�P�]�g`���*N�C���l+|���v�o@�#˓���^�ϛ�1������>��8#�H2�O�=W�?�ww��`����A�pYg�%��Î��H�tc=S���q�>�NN�ZQBs���L>��~�n	��Ȟ�Α���t�C;��o�;�P��f�gQg�S{��墙A���%iT|[ݻ���V�b�
+�13Y
��t?�9�-Ķx7@��� ����K)GW��߱���J���e��ےK���
_�s@���~�anz���_��gS�":��%��"�D��t'����!)f3�|��݇�;��kUѬШ�%-aQ~`��, �?x�{��ʫ�����a5�ǃG�5C��Ep��	=q�|s�+�Կ����g.�Iz���1E�@�sX�t6���)�<;����郻X_^D�K�]�Me��`4���A�>�}��o�c)�M�
[z��/xɒY��E�:�70���_C���Ȯ>�;~G�!h�*����x�/� �l��*U�w��.�3������-�x_ٝd�w~a�ӓ"�O?�tG�w���W���͛x<5����({��u�ο��G��,��BeΠpf��3�:�B^����޳9���;�� Hx[@y�ڳ�n�4�C�rvbv��������"��B�����=�Mv�m������@��gJ�����k8�	!���P( �}�{�y�s�s���WK��R~�'����������1�*�M�\�&SL�V�XŁ�G1:�_ë�r�k���[�ޗ�X_0���1���F�N.��d<�d��}�1�wǱ{{/F���� �]���"�9VP5���+-��ZI�u�q,K_�͠6^�m88Z�j��vD�:��_�~�t�i ��N�����=�?r{��7֊;
d�ĘX[3��"~7��:|�2R�����G�07�P��Zb��}ٍ��A�
e�%�]�A���@���gwq���W��T�j�,����=��d&hI����[�g��-A�v$��ݎ�dі����M�!�(��j�j������+e �և�޿)�i�/K`^�(�#�-Po�v��=���}�?�n����;N �
8�!�u��EkD��!����?�3^�ԸP�R�=��o�+�=>\�zw�=�͗����ی�ؠ1hr�sI+�j��˕zqJ��4<<���>���I	�pY\���M�u���;G����fׄ�k�U.��JK��B�
��X4�1N�Œ-/�KϽm����zz��'+я��L�]Y��:!�L�3=��5�֖�6�MՇH�-���M�?�L��v(\ٽ�{�hx����|�JX]ߐ��ȱ�ص� nݻ��>��u��<% �d�.^��i�kj��=���t&��M#�!�cq|��Wx���ɓǎ��3)�%���X���������%����1����J&����'���L=}$�)�� ���:j3ϧ�8�vw�� �d�6���-6L�tS�`΅ׄ+����1����1�m\ZX��<CI�,��,g������/dϹ��!:rK�+��w�Ck{��?��091�����r!���0�g7�9�ё�S�`���-������kH$Z��GbQp)�C�k��ƃ~깺���+-^u	��L�ּ�H渜<�ФẒ�]G=�O<��b��B�J�ƫY�9�ޤߏd�]��@��x*��g�k�N�x6,/���P��񘀭��a=#�sz��� ����-�lt_a�g�׵X1{��H$�ﱺ�n��^�J���9��b���}f��Dk�l&���B��V.]���A�3�9#A�'V���A����ٳ�v���{wp��p�� ��t��Y/�0�vt���k�i\�}�ӳXe�\, �f������T��֘��kՒ �w�}O�i�Ծs�b�k��o�;�,��ͦ��_6N%� ����t�����y�nJ��Lm��D+��v!����M�?��]��K|��c�)��~n���[�/�P���z'|MÐ����4� �48�G�����������ܐ��r
��dݚHvj� ���[�/��M��7^ś�E{""k�|.�bքe%Z��B�T���͌:���\��[�Wg����&ju7�ј��F����%��E�BQ��Х��c�{�� �ܳh#�΁��x\2!ɬ�������l.Σ^*��!�HQ�'�R�+g��G���I���` g�;���Uʚn\�l�*5o��2߽��n�;ő���֩C��^F�[G�O��1�m#���S��?�3u��u=�,�Y���r"ӳ��<���cuu��z�O����,�ݸ�ߝ�w�����<�:Gq��w���	T|��t���C�Nb�-�o��W���Bn�g����������� x�T+ԫ.��{۶�B��!s1���	/�C ���ƍr�������`�>�ҰV��ӏ���:�Z����ŏְ�8ĺw;´�tW13��Ks���Q�5k������3�W7�a#���b�=u2�1�w� kœ�y|q��d3Ţ$��V���[R5<�� �<�p�yg W)�d�)���uW�RAa}	O�����W�83���Mjy_�H+G�bס���vh�6_,�MC=������m<��5ʛ�����l�@{G�t�>&���"��%��ښ@�t��0�݆nV�4�*ٌ34K�N O�f��eJd�@'iն0��
]=,��CL�bA^��^�!���-Ců�~r+�Մe�uv�t�j��P�G�L��6�E���P�����������{j)��t����͟���RC��]�y���J���áo�����ζ�_���&h<������±Ç16�]>�n����L��}��S;eRi1m��Ol�L�j�ϝ;��o߹�RB#A�8ZJ��^oݺ���9�$��7���gϜƶ�^���+��ssq~�sA*݉��a�0�D�=Dfm~z�+���_�9)7jڱ�c���n�2XYY���)�2�2IҲ}d� �gg�bniI �艓x�7���S�;Y]4"�c'1�ٳۇ����a�ٌ.\�Z�	d���dB,>�;�9e�+�N�\荞�g%�q�*8u� >�][���cE��߷��	�*���SlD�V�\���71?=)� 34�����ū;�G����(v�>���i�ɼqx�r�����`+���p�
�V00�Ml����8sZ{ ����A�����~��TI�t$�6�5t��H<Cj}M�"2It��gx6�����dPi�GPI�E��ÄR�I�6=3�$Bv����moӕ���3�+ �N�a���EU�a�|� ���� ��>�"��E�*��+��c@^wg����66���>�[�x>=��M����v��@&��-���[s1�[���k��Q&����߫�m�6t��cyy��Ma꿹WP�şc�7��Y<<���ײĽHN<������ʽ8[��ٔ�A:�^����j�[�8p�v��Q��tҸ}�.�;���D4�HЋ��ҁ�
H��h�����9\�{_ ^TV �B�ȡ���ǹ/��d���t�����U���A|���`!Js���#�Ǎ�R8��a�Ά���fy$�1�%P|}ܯ���0�d���7u�_&��ˠ�ޣ�o��>�a�j�    IDAT���l��y�м|��8pR�-��,�� ^��JA794;�����_�����33�p#��F$�&�J[�[k��K��/������ѻ:�n\a�u�����Q&�{�s���ʱ�z��d��_avaExK��������b-����"6�yx���!C������ԧ/2����0,��,�GX�|�Kg~���pW�`w��0����[�@X���/���cۏᑽz=�pT3��m6�ל ^m�zE����+�sd[Iv}C]�qL�UΡ�K!��b�*�Gj��Hؙ�ͨ�O�խdw�LI�d)�C$Fī\�|�/_�����?�b�$>����ku�L=�z����8��{�w�T�W(��\kb��C�2�(��O-�3�?o���W���s�/7K�-պ)�х������o�t����h$�WUJ�o�И�|��Bc�����6�jI6��0�k+��W�S�#!ٚ@Wk�He�<������z��6���gZ�V�h���Vz�AQd�Ar��.:�����/Y����z�\�,[���g�lzQ:���#8���h��F{7&ٙ�����j���
'��x��W�cf�>j�2=3�?V�C��F[�6<�:�v�O��%���yW3�0q�2*�=�K
 OJw�3 �m�=���xo��́����h�d���?5�.���3�M�k� kan�LY o���=���eJ�ۍV�a7җ��MCD͌��s���M 8���{�>�:����B!(��e��l���CSj��]�rU��f|�rah�~����f�_�.��z�ѧ:Q�ZO�8ŀXg��n�3P%s�4��-�i�,`������C�9<�j�d���%�U�R����5:tH.C�d�y=�_d?��#�2Y�z�U:|X�ifnV�<�֊��$6R��~�n߼.���_]��O>���z��:53eXAZG��T"of}3�&QH��V��� �JM-����رsԸ�K��s�B�t���O�M���I�ii�	�ȱc8~�u�{�g�]P�M郆w=.�3�G:-y�e��\dQ�&�L���w3�dĂ���n�xz����rpb�]*x��|����\Z���{hOD1:��\p�=�/ǖ瓓�5:�0S�K|nxp��O<R!@yK|�%p��D'F�@{� ���%����
	�t�Ԏ�0=3���be}{���#G�������y�w���+ ����V��Y��g`����=�K뛳�=R"�ޱ]�=E��?�5�5��"�[��=>9��hѺ����%��$'�!f���¡6n�ײ �D���ū�^B�I��T�)�8'�f
m���E��q4	��h�����2j��k �G����!�<�?��EkWg�:���Z�\w|���=ؾm��:Tq��Z���֗�z��|����g���`ucM�B߀����$l��D��u�{���@1�\�I�֕���������!���Ҋ:�d�E�Dwq ����!ǆf<x##cJ�����{�soݾ�_�C>�F{���Vt��*M���.dmI�r\�vS20>����p��!<y� g>������sI�x�\u�����Ε�v;)E��Z�V�A)jv�h�	�E�8�����<�+c�_�k�4��3l�t�-[*@���"ܞ1��e�-���S��d������-���� ���LD��ϒW��-t��f�Ʀ�;A�|�$Ȧ������-N����±Z�
��O~eywn�@������|�4�<�}n`3lI����sh��E�%*�I��?��>�,���vѶN<z����f�sXKe�9`ϵ�����Q7O�X2��t͡�$�fC`V1y�&�����tOk��U�MY�p!�O8�H�m���uIFC�����@6���̤ٲ��U{�M���ק�^��{`�0��ۉ���
�kH�/I�`�PX�I6#�!	dl�m'�T0]ۭ���G�~�xHI�_|����џ``p;�7�w�\�u��N`5SC���w�F�2�w�i�k4�;{�0�f <�J��b6���x����=��_`#�����*�M�P��0E1_��®]{��3�Z�:���k�0�l���hn�1t#���xy�7@�*������O>B�X�0-٢h�"�#�b�H�|<��j���4��ٙ-ͯ���l�3w_l5e���t�T<V{{���ۏ�7�'ӳ���U�����!�Q�����/).|x�(������8I��ߟ	��*)$ DO��&��̎�Ca}�R^��v�44����ڻ������NT�A����V����<r��Yx=M@w$�&ӅH<!om2vF�'���H`[v��-�B�R]�9tam��,�!0����<cs��z�ۍ�l�����-���jJmk�����!����n������o�=�^���^������o~y8X`O�_G����E�x:���F:��`cC�?���kI��]����4f0U�s�շ�!,��d��|H��Y���( ��z�zZ#T�vw���$_�0���g�O�}����7�}xX�i�>B?J��L�Z�Z�A�`'%?��O���&%C�b��_��NC�� FFwI�L�ĝ�|����8r��ܽsK��Rӭ(��:gN|FrAF�<�B&� m1:�PJV��<&Ċ2�h<.���Ĕ�������k
���x#�p��x�7p��qܽ��ϜC�rs��k)@�
�8,׆]��7ܓl����NZ+��:1�J�AÎ������{�x��6���18Ѓ��Y��.#`�Ǉ��2:;XT��]��=����[xM���j]�4�=�ޡQ+��%y�Ǣm�
�r������%��w:�9zG����>��S]ד�cر�rI�E~^�6�!v���dmY �Zs~n�d]�IIR����K��Ҝ�Ǘ�H�P�^�*���e+֞�0���$��`T8�	�6��5]O����P�g��Q9�=�"N�8��[��\���޼VVB-�ٸYh��ܴ�d������A���Y&ߚn,�Ȏ�n��e�}������������+�N9;��!@'��7;;'��uğ���-�}|���3��SHڳ�,E���NW,��K������!%jn�U�:r\���۷03����H�/���>E�^F��Ŏ�~���+��lG�k�vv(���1��]���tVk�]+vj?���C�H��އb>��G�<|T"e,Tx-la͵�N����
i��>�Gؽ���Z�}x�}wd������Z�g8{��/�]������C���W^f����-��a��A{�9h;�,�����}���u�_|�H,<|4�_�1�>���J��,)G.��;e��w��G��%���@��G���B�Sn}�w�u`fi�~vO'�Q�zKvax�.�؅���Jr�c�<��+��M �.V��4����R6���@��K3��k<�}�Ԇ
�\���1U���I �5���Ab��uj���â>Ӆ�C�dй���%�O��<�WΟA)���v��at���T���Z�@�R^��X\�*g!uO�&��J�8(��d <�=�r)c��h�hfpzv����;���AL�.���׮���4V�U(o��>�-���-�e�	�{B^���{�Q�����bvs���d��g<�X?�y���ҕ�J�Í�7���}�V��J�����[k<M����' �ڡ.�X?�ayf
g?��z�}]�M&��S+�% ص�;��w�P̧��2���孶��l嫇�1��ś��,W��FT���p���ɮ^4AL.,�ҭ���$�_[�bjzS�K��ãc8������t>�	�բT����U}zh�X�#��>>DL.�� �7�}��D��rY�s8�R�
�M�=����{(����� �l�D"цDk;Z�,�!��ׅm�����!�ah��@�L��"q Ђq�3������f��+Q���i5���h�	�w���KM3xo�T�[�z���0��[�/�����G;��y@�0��F���$��nVl���3��@�<�r�џ��P]�z�'�P�r0�2ZX�q�6b�#��W2����.����e�G XHo`��՟�q�����a��~����������O ~�k��r���LJ��;Z+R�͗��_�Rz�w��� }�Ϝ9#&�s0Q46YJ2�۶���Ò��P���{4C�`����$�&�QH�F
�T
!���E[R٫B�h�W�h�= ���������ڪ�]��������c�܎+׮�̗_˂��7I��u����%� HSԽ| k��Ƈ�dD� :gƃ��V�U�9����ￋ�������ۆ�l�)ܻ�=�5SPTowz�;���W��w�&�O������@��p�,��EK4�GN`p�(2�*�W�d|
�x�����~>3���>���믾��X	�ȶ�P�L���*igix�6���p��=��C۰s�����Ԧl�躳�����,�,*؈��L:��n
<�3��b�	D)�1L��F(H>�������X0�̤rYdS�����Qb�̈�.3����a�๞�ޮ��JV��q�1�K�9�Z�3"a3|����^�� ��H���a8~���ӿ}�0���au���Xx���M?�V׹��ʔb��F��|������z�"����<���th��a��5 �j���}�UD[�p��	����07�����{ݾ}W/^P�<�=c#��ｇ��N��W�$!�K�������˳XYO)msl�.���M���y��So,���x��q���w08�]�\3
tri�p�`f#�!�,q&R���
�Xw�	$�V-Yc�]��.�ci(��-P�4����;��g�� ���43��8'����̲�=Ӯ#��|�m.З�O��9A����^�L��q�>���x����CJ9��I�o��_� �{�ڷ^WCs#d�����$�YS��i���~��׸�t�lE!l��n$:��p�Q�+G�E�"YlW�%��癘� �*��P� �E�n��5���?���/a~�	�������r?����}o�B{�0b=��aW� ���%�1 �c�"�$K"A7RkK�}�<�4��. �V����Y�BfC�6����.���fޏ��$%����r�Ӻ����Q���D�>��֔� %F�h;66sX^K�ҍ��r�$4K�
"�x���q���({^Hh4�ߤ��������l�,f�+��� ��.̄~u��_.���)V:��s%|a���EW� u�#�aE ω�!����S �����5�05��O
_���=�jm�v�U͡=��];0��O����l����(u��Cn��ٜq�������AA��:pl+�|[k�b��n�-����	T~���ϭ�ɓ�J�ʖ��>�G�x-�H�j:������u��y̍�ǧ���k��]�n�rJ��\q���Eѵ}7�}��A�t�B�M���=���CT��b�;����:$�;�G�hmmq��l���0{Z��mV�Vc�Z��4��՜���9�C��c���\4k�m�������A��L��[3��-��̚4k�fi���,����,��X����e]h(���ɟ��Fi�~���̈�i�������y�XϚ�'���՟���ꍻx�x�,%D�fG����o0�67b������n}L�d@N0 N�n./bg/�y�ui�9���Y�'�����W�\���6<���ٝ�I�e���0|���ym�I��_��ؚO��\�3��.�N��*?~�(��d�k��UCJ��ym�V�H䦗ʤ�`{����i<{2�<BG�(y��n�ٮa�PKd����6��KG �ozֳ���d �����5�>�.^�,f�Zw4��N���u�tw�,X;��Q��Y�쒨K@��s�i��mh~�V���؍���Ȭ.cj�)��	l@v3��Ǐ$� �\(���C���xT����ۘ�y�`��HK@�#+��=(��µ`dlv������03����.�����{��}|y�+���>�8�
:"��O>�D *���������.��J;'��c;vˎ�ýL���M=��Ι�5��T*�佲 �CW�p���s?][Y��J$��T�����SAςS�#�k`� �Z�I7����(I�mzyǗ�n	�vC��L��2�9�Qv�B���d�	��ټ :;�<����{��)C��������l�_3��mm	�)g`meYñ�ĳpp`��Rk����������O��� _������Wq��VAĎ]�X�S��knwvl�����whvd����t�
���bdlT�K���#�)�b�ہ?��?ƶ�2�RNo�0�������_bym�`X�]�Uη<}��d��ZݝI|�{�ᕓ�%�!�a!ǵm�',���?�<�^6ù���RP8��w#�2�
��������:�4%Y۟i�3��%���1�g���=����߫���~ل����{Zg����eq�e��ͬVP���]0A���_�ų���@�T�R���
676����;oc��]���
�sS*��m�!�D"I�6��V��Wp��#�ϓMw�22�@$֡�� �u,!�_�ҧ��+B�9)��|&Wu��J�(�O#Omd3�YL?�����avr�T��w�[�����#�֍x��X��un�2n:�z���53��`�?S�9'�RA��^]Ľ[�᫗�wg?��߅d�/�w?ʨ��hT

'$c	�e�l�M�x�CA��v-KvG�6'ś{M:�E]�RA�c���Y��#�����{�џ^X���t���R��x�0^����S�4�143�<���!ց� �t���K�-�k?�������G���?={�/�ſʖj]<T��G�s�n$;��v�o�FB���;	��*���fxx�0-~�@���8�~��6������@7��Z��s ]�Jl]Y���������@8l6�5Z���M؀x��s3�����Oىˍ�܉H,�|���E<�^��E:W���"�<����-�{����o!�օt�N/*U%�|�<f���}����/�,J����	 ����}��3�W�LN�^2��u,L=�ܳ���6�,��ա
�<7j5��;�g�N��E[ԯ����t�VJJ^�����n� �	�\F�n�� �nBV7ʍֲ���`R���ym܎���"Z��s��7Kq��l��	����5k���׽e#�I���w���аi�"l�sc�p�Ν;�t&��Ϗ�]{�G?�Ju�����\�6����B�����S���3^T(/r�y�(e�4��AH��u�����_š]��>_[]�[Q�o�.�y]�r7oܐ����v�G��1|:9�a�ɩg8v�8������Μ�
�}���b�8G��bC���;8v오l��^�jP�Q�E��V,Ӷ�.
~�p��,���$�ݺ��糨��]�R:�@,Ǟ�{�``�V�i��^��s)���s����q��U�?��0��t`p��r���kεe;���hx(���.���h+1��4I�5;����/����k�>�鑅'u�lV����
����A��M�Hڋ�6�L����Eb�T�Z�;004�/�gӳX�H!֖9����������H��b,�|�[
ta����~/��m_����78�`$,����'Ot�Á�|݃~�{�jE�����z�어�eS˯��A-2�^)?� s0�e��m���s,YiV��)����Qvdz�{��O��Lz�"�ժJa�{=b߃>�^�4�����A��#;Md��I7�:��97��{>�'ڼ��V�Z�ټ	vcpR����Z���Jf��'��l���]5��e�H���];��Pњh����C-h>��"�ky��v��5[�p�܋I�q��[0��,,��}D�#F���Ս�'N��t�2=W�i�=    IDATqC =�l\��R�Z�������M���?-��D�>�g/]Ņ�7��������Cg'�қ�z��=����=���w����K�ǵ�5��U�����z]����A�T�58Dآ�Öl�Ż��c�k�n��|~mg�?�v��P����ּ7�󣙁7��3H����5α ݞ_�wu��Į���k�䏯���f-Pc:N^dry\ ,@ӿ�t���,���@�F,�á�:!��E�%����"*�L2#J}�9���9���b���3�r��4�oD,�?Ҋx[�l��´]�HvE��@�/����� >G�~� �2�">��QMob��Cܿ}Cy"�a�*g9���CqIp������h��hkU�!�Ë�=qI�W
��`e	���G�U��}8�o;:0�ӊZ>����(gS�#h��3.�, ��Y���^'�����sZ�g�WJU�'Z�K�
���X^N���+�dJH
���<}>��l]��x��`��W��+!]�(����]h��ihFh�\��q�#���up�Y�9f	���������\ʔ�:_it2 �/#`;q��^%ry4����4x=<�� ��I���*!�b!6��p��dG�c�c��ر�O ����m��Nh�u}���ق��]6�5-r2��5!�g�����k��g�
�h	q#I�g5W�cbn3K���X\I���<&��bz~EI�c��ko�M"K�����j|�낿Q���$��	�g��|%�r>�@>[N�A��n]HJ��cK�Q��U�kv��,M=�N���P_�<��Z��!���n��K�ޕ�#�kH�����9f��ob�Nd;h6Zb����bK([�(�Ej�٘��ÍJ�S�F���6��;:�\�R�����L�˛�˛�f-��غ�����-bg#�?߲�:L~��(#	�u��� �����ŋ��g����T��}��5�Ɲ�w���E��mT�GI�Z*R�� x��]m��	Kk惖N���x��a�5fR�8)�$V�W���΍ow ��	�b��&D`��5�������zK>���b��zRd4�����O�o�����g�cE9-􊕪�ӋKK��4!�/����Z��SX��%��t�� ���ɖ��Ájbs[�#%Y
�`w��4Ո@]�V�P*V�C-���	��8v��Hz�=x�;�t<���$�%�q��{ĭ�� x2�;y� ��޷�:?��g>���|��݇C��Z��h��S�c�3Z���I�(�0�R� D;Ѳ�_�d�]�s�����)y}�ɴ��B��T���?��ko�.����3Ih�l�9fA���R��ӼF�JK���<�Г�����I��^�ߗEH8� ����dJ	yh�B��|�jUOj�O�tVRZ���0�4��;���o���ץ@�BnC�r�l����-�w�*���%�=�,(��d8���jd�f��.\�|V�^I�����e��9E�����%�Q�j}�.�v�#���~����d�#��'��/�=v�Ȟ���������,�������5�9�}S�q��{���� 1�9y-)a"��i6�)�j揝8���v�ڍ�JԵ{���"r���80X����C��	�
�(�+� i�bb���)V��w�ù��Ff��7^�WO����z�Fw�^�@,��D�[p�7̬݃� ,�3=fﱺwI*9��N_�$d[ݻ����{�-�W�u��0��x39�r7�����i�G ��I�a�O�ƽ�A�:�u��U���XY
�5	��)�z��w~a_}�nܾ�ŅeKy�fS*ƿ�G�����hMą-Ԩip�x1'`�^���2~������+��t�Z�	�����sn_�`T�J�� �?�C�O�j� 2��u��!����,�^. D�`Ћ�߅Z!����F��.�n�R�p4�7 �?$L�T�޾�Ca9�pQ!W3<�@�QQ!�s��:���k���4����o�k�����s�/͢Fc���k��x�m<�gk�k1�q�+��7|f�[Zdd��}��V.�⥛�����p��y<���F�����x���cd�a�J�o x��7�vG��T��k�u�V��Ǿ���ylo�s�/����p��ҥ���ܝ�
**��bE[{7��0������W5�À/���8��waz�	{:���O >&�?F�{ћ��/��%d3i�M���Ir�����ux;σ� ���&Y�(:<xEÜ&N"W�aja����8�=_�Գ�:=_X�?ŁS�`ϑ�@(�l�+�E&qP�l���y�r��,MOȷU��2�\rQ�pZ��bI�\^��u�g99� �:3��Ix�E9��0�����p�=ؽk'���(���W^��Q)+)�}�Ń[�L3�L�����u�����m���HY�ݶ�	>�Z*�0-�O^���!ǃ����,>(vU,CӇ�-kѼ���m1oY[)�6�Vs�8�M�Hq�"l�3�2�����7���?}�K<|���F����տA�Rǵ�$�!�7Č�}w�xAz.�w��P�G����<�WW�f&�˅��A�v�� <����K�����*,�gZ׍���C���~���O��o�Sp��;�蚟�xAx��|X�R���q��I9d��L�~��.�GF� �mn��ʑő�PX�)x�Oz�ӎ����G�${����2�]Jޣ70�\j]�lmZ ��j��Ӳ΋@($��J�\^�X�-ͩ��K �dE���V[�JeXDؐ1�0��tK+���5�:r��u@|u�3<�{[`���L:d�*qWWV����f#�S��7��sj*
9���\��<������QY�!S�PkO�X�.,��B������s��FZ"7�/<�#��]<x�u�M�t἖������3b����s��KfH���ָ)�*�Y	�:��!����t�����f���������E� :ip��-Y%Cv<���P9(��X��|���$N�5<�Y�����稣�6��|]<|	�	�t��ұb��@ �{@i��_G"�lrݚ�ˊXl~k13@K���X`����0�������v�,��>}=_#A>�H���2Q��/�Dqj��=�  ��e`�ɺ�ݱ}'n߽�;��#����&�z)�W��DNg��C}�S��R�r�JKY,���K��P,fX�23��]�o�o���x���ti�וד�Ǹ�HQuS��*��t0a�g�;�V*��b̂w�V'4��)V�I��:��t�/ ��H[�2��l���I�w�sTz�� �~ޞ��L���4K���G�gI(+3�;
�:��� 9�}wjj_�>����ˮ4�ɪ�I�b������Ȩ���Ev9A�|f$�t��3rY�?�;��y�◿�ח�F]���Dh���/W,o�E2�P8*�-PM��-�q��!���H���D��T��+�1�g�6&���zƹ^�?��@��05��x�U���s�=�V���3 O	����Tr\��+��gp`l;Nڃ�d�Xݕ�u��SI�%���#ߢ���.m�~����V��gf�:�!�8�<4�����"���̊�&�h���p��gQl�0v� |�����!I�aF���bm�kYͣ\H?w��G_g�<4���g�/��W���_k�<|$���$Z;�=.�^0��0��"yIBC���j:w.�@B��q����q�"ڢA�PF�ߍ������z�h�zѨ�y���&Ye[�R�}'��dK��0�b���$�ܹ\5IJ�UN�G�w Wi���2R�:JU&��|vE ~ny��8���ۃR#�\�L#�����1��4�(a��BN>�KX[ZB�d����QcO����`5j(R�T� An�sS�\x����]��xG�A�}� �݃��hm�#�o(¸Z�jH��w����d�U���XG.�����8i�K�~��4��%��فp���ת���p��Mm2���Ì��-o�hT�yt|ڷ��t�[�͛��:��XV���Þ�~S���b<_/<%(܄���+�O�MA��+�p��e%Mnۅ���"S����{��db��ԉ[V�Ai[��aS�@#y��r���Mx���{�0�{�m��V��ի�U��ٷ��v���K����(Isߞ����d&�Ǖ�M��w^�t�7'8���u�/��޾>�zJL�!L J�O J�����<kr�9N�>��g�:��޽!Y�I�R�nf��H ��LjP�����M\P����JE����z���խ��a�	[���2�f3���Z;,�<詣l��W�(�ݰ���E���Q�����܏�~�M�\u�'���)"�	H.G�R�h%�s4�Cjh5ݣ��M��u{�U�p?�|%
�P�JM%	J?�Y(�A������Qh��$>��sl�nj`�O ��y@LV�P���(�0�P�jgBZZL!�g��$��S�\ow�����j�cfڴ)�(w�dr
墜�/��H������;�Wu�bDaf��R=@���a���ȯ\���,�	����BB��^#� �7�I���b�l�էs]��g0�OY�)�M�.��s�y��F�d!��Qi+��Û�U�X9����`��=?����%�$x�� ��NgIYN���4I^WX����&B���{�������֝۸���!�e�R(2��=��h��@7޺UM��O)���ȕ����z6�s���zo���;������7_�k��D<������݃�.xH��)�W��+�o:��:kP�\��V*a�r�\�6}�sf
�f�g�Ѿo��@{3)���M2��A�?	�������z{&�"���m�@�L�1�6�	+/$��Z3F�s���¥�r'{���)�	����dr����ql���b�M@��B�OF���t����
wO ���w����i85!���o��D.�<!�od��+�M������
�Ms�˿3��ϓ����Qad���Q*�R0�_}C8g�5�P�B�<I�������W.�ك;�?2���w�?E5������pv���daJ{^w���k��C�_>��tp�ۢ[�L��"��ü�d{/�P�X��Ք1���K�t��--��҆�����o��Hk7�R|����~� ���cIt3>�ȼ�*�̴�Q�_;�b�ױ�G��<]h>���_�g�S�����v[�������?��y����6��+�~Iƪ3J�JhJ���[�>v��ҹ3������cd�=��:HƂ�H	R/ߐ�mk"��NK�k���M���97R�z�Ш�9$9l��T�Kg�3�"�x[7
��rX�T��JJ�}vaUL��Z;��Ƿ��.:�IӔ�J��A5��hɰ�p� `��R.+����q0��N�O<S]�6M��n�B�J��\X�AneI�����݈w&l	��-��{F�ʉ��KH����^-�\�
��s���"[�lrB1���ϱ��T�m!��I��M�9H�Š��O��}}:px�؍��h���S^w2L�O̓��gy�I8��$����n���hג���&���M�}n�֊��nS�,(���kc	��5iΤ@�_[���᥵�g_���[�0�m~���l	Wn����y�6�h����-f�q��ɀ�%I<ҿ����z3�lz~յ*��؆��.:;q���8�J�"��8�#Ǐ��$YN�Rkm�7^k^'����?GzsSɜ�����\�`��xϨ�>��Y=#t�!�O������)!����w�ٳ����3��TH�ʃ��
�h�{���x�X�I�L:��NIz�R��n�a�?�uH�M�1{�����X��0s���d���qصiNj�%��w\��"V^oD���g��}{�o����.�k�4Jh��(�(3k�Z�j-s���R灅�fzC�R�,���O>�|v����t&�z�dRu-n��[��`)%04�����[�h��GH�E��B��J!�!�ll�$��x�&�S1ˁk�	�
]�$� h_X���@/��������(�aw�t��b���Ͻ��=�a
-�I ހw^g�2�\faJ"��;�Hܯe�ɂJaF��F��"�1U���{L$�'9��<|y�X�YPm72nv�Q�G!�$GJ���5��3���L'�t�x�o�"u��d9��?���������=н�]&�<U�!AA	�b)����Yf��g���W�_���OD
�|��K�g7QL�y��ن�v�U	�d�J�ZCnk4NXN簙+�̦���
���)��Wx�vʓ^y�$�|�U�D&�t,z�gc��t֕e��X�>��ۤ�ZfZ�������Z�m����g�מ ��㾉���,S*���h������w���9����.�5{�e�����ŷ龎��:SN�*��l�3�q���h�Mz+�3�ן~����s�.,+�����C��ء��B�.O��u=s�[�s�$U'���\�����q��=y�y�y�h��Ck�o^_��фb�%������ۣ𹹵V3y�&=���'�;��@)'G�5�ymd��1%�ρ�������j�C,�<,��5�r?���:�������Kص��F���ւ��"J�U��5���F
�Y�`#�Ҟa�@^{1�q�WIp���2������������=<��l��sȕꘘ���Ϝ���3�,���ÑW������	a5SD��B���<�5���]1 ���Q/垹]ſ��j����]K�,�����?�.��T��]*�P,T�bxx����~j�����ߥ!4��dl�Ĉ��&�Vr�����=/F �B��\�1�M=ï�,?���vb�'�D�o��֨m�t����=I]T��َa8>�1s����En<X����ĐǠ�]$�=h��G����2�L<Ǔ�L�/���2��/iB�ȩW�ʛo)�z)]�jh�Ikk*5&��)�2J��$@�AP�W��䁨�X�bN�1��i��|��&��#������$�{�h���m}]8~d?��A+'��^�P�et��7�Q������������_��'O��\*!3lz3�n���;�e�h�~��	��q�߬���P��� ��xx��zy��"C,V��W`�n�v���IuP�0�����y��Z���7��u�9�ʂ���sp���w^3�F���~�;|u�"ZZ;�������._����yd3���*xe����c�v�6]mд\_YVK�m������;1�S�:�)g��uf;�\��m�����T����د�m�vhc*��X[����{��w�烇�`x�v9�p��϶��[w��鄞Y���Q�R&kY5l�U����wÅ*ɇ��F8F]gP֨�UK�N1%k��
&.�qt|��\�C�����'�CQ��L����;� �6f�o�iV��� �R*5%�2��2�:��U]�=�vK��B��e�Au��-�DW���� �C���vpM��'���J�*�������}�P�Hq
2J`��K$�O(�Ϥ�زY<�{w��C:��- �iC����dg��z�w���#�6�
�ղX�[];u7�P>'��R)�u߹}H��-༎�,��^�iyX%CM�+3����>4t�[<�=��f��1�S��s�ZQ��Ȓ�XoZ�d��~�{��a0X�!7�w�cj�M8{�-R���=���3�s\��s��,
����ٽ�e�U,���;�5i�-k,rk�)����;�\��`()�x���*"P8�Ji���K��uX,�i,���%��~i���lC��4M�T�T�,듩L�,�J�~���v��r�eҔаCA��?��N�±�57Ä[�?��;W3$�U�3a���3�����Ʉ� �G[@�߅'^��mx�� ;�i�ۢ��^�؎��E�����C��b�~o{�(�<K�얙��FV�i�[���WPH��    IDATګ�*{�ٵ�L.�."�;ShH%�o��
�+�p��}|�ᇸ��I>��$��}�ٲ�di��O�]1ה>�To�����9����/p��}eҔ^�cm��B�K�&o�E&�P�@�섃�Ȩ�Ϗ�Lk٢֎'��Xχ�wS(�Zl95��9C�־��(SǙM�E�^�c]��y�`��@�X�.���13��ϟC��<���ba�J���A��$3�h��|�Lǔ��$��bF١�q�AdU9��x'vTǵX����^tv�a}#���y�-���ͻ�q�>Oϡ�w����}�ѽ���`1�G�	HRI�=�:zAw��s�MK�B�xp"�n������sgtYk�im�d࿼}�[�����b��\r�P�#iU�O�q:'��a�;nYh�`�Ƥ��%�Y�6��g0�|2��sc�篧&����:���<�wC��wm���m�n�JF�ߗD{""�t���b_Z������q	z�JF�-P��2����h�Ff��w(�@kg?��6y��O�b��,f�11����9M�Ǔ�8��[�{���6�uY6o�4X���B�N�,- ������(V�.L%��W
 1l���B�T
k��Q�l �=G�#��n��a���8x`7z;d�Ie.�b�^���0���MO?ǽ{�p��I��lR#{P�k�`'Y�	�y�v�ދ�'O�em8�ƴ���7H}��J&AV��ϟK0O ��L&�)u�/�J�v,谋� �!^�<~�&*&����k�t�.c�����W�����y��џ�;ld�����Cj�Cl������c���J�h}�J�K:�h3`<�Ajs(�������@m8;+��4L+��/_;�S��PDmX�1mىdkfg�~��X��HP*Nw �@�~��?O��t)
���C���L'+�1	��AÍ���a�h) u����%ނ@�/��}��i�Ɉ=�	x�G������k!�gD̞� )~��xZ�e���[g!zU�ڸm-��+dǬ\��?`���[ ��Q^�!a���B�>��O(�� ��L+��R�L�oO�Ԓ��t�{#�*t�iM$���1鄠��l�\�N���;m��a^�	2�|�ݽ=���e�Գ)tt���S�)�'R���� 4��/�Y^��s4
��C{ü:���d�y}(�1Ϥ��p���u�ͬ; ^]�����Z	�2��Jʪ �W���b˟���/:r�u��c��xϹ����c���5b�}�
v�h����^N��TZ �2y`י����kH�c<�-x�w�y_f]���7�t<G��:�d��%;�L�����G�՞y��eLML�y��W�������DI��w�E�E594X���tj��)�\P��%S����r�t�b�t��1�8q\i��ϥ��^M�ퟎ����<k�������|���0�/����$5s{mm�ۂ<{��	�f�����v-�/mUMZwˊ3t��4�:[���]��?_�̙�j.����k��p�s�_^O~������%�ǿ�D2U��|�����=G�油.Xo�����4i��O>ĝ�d�]���A�%�D'�"�J�BQD"m������Ge5��-��S����2SM�֕�y�|o���YY�3���սu�T�o��Z?R@2���K��"<�::�T�Yܿz����#%�iC2@k���(6��֕�C��.b�|�	�4�'�S<�Y�q��\1��5��>�,J%["	��Ax�a����eqy��?���n���qL�-!����������T���F��5o��OE��@�*zZ��/�� ~"����1�p�7�����9���˟���\�?��]��Rm�v1�x�����w�c�Ŭ�� ��n���nǴJ��l0.�K�T�Mh����1��.n^:���x�����)�BG�>��`��$x8p��"�/"��KL�O����XIa7<<���S*[ �q�Mt Wl`jn	���[\��򚪩��ExB-�w�8���Z;���+!��n�o���Ei�r��.u*Ȓ�r-VKb�����X �gb+*y��AysS ��q&�D�hmAkg+ڋ�N�ľ=#�Fئ�E�v��nnb3eZ�j�zMT��{�q��e��=����	�:�U��v~Y���&/�E�l"������צ�����������`�����͢�ب�-�bj��mm��!6���3�����V��^���(��b�7��(���aO�k5m����{ ~y3��������n�>�*�Š������!Կ /�9��ph��olj�]-�)���@��{��ކ��v�e+�@t�а�-6L�1��ɨ���/(�XZXD�d��~�̑�����V��π�b�:���[�v??�nܺgl}�c�ң� ]�6YhGf +�f��w���ZI�M�+K6G�'\a=�%/��M�	����60١�7�BΚ�!��^$op������?�%��d���'�7�{E��Լ��%�f�5�Nh��M�
%�j�N����E��Q�a�>�#@��s���Af�AO���tJ�ގ�����dǬ�9�%��f��9l�X�r1�$dx�Oڭ���i�}��1��W���B(b:7�k���PC��:�r�d��/ic��k�dz��:;��ĵa��k�H(��F�h�y=xxPkf(���b?�v���T����¡�2;ZY�=�{͡;�u�8R+	�
n�՚4�%��vhs�hz�5n�[ ����}��B�����kXt^G�-ɠ���1����4?�~xv��'!� |���"�����{��J ��,�-�p�3���2qV̠#���A�w~�ߗ넞���V6�)�:���op�a/��5c?��ۅW_=��ǎ��=.KL�?�sm1ün6��������,#I�������ޙ6�HԱwf���%�`�	`�{e�msQ�N������{�-��^�	���[](ǉ�q�7�d��ڲr�v��=kl�`���H�u}cQ��mڵ������f^�;�]p?��q��U�C-�а���rk�º�TU���V� �iM�����2�C�w�v���{�-�P.`�VZb���p_$y����c�`,9��;�I$ty͹�G(��H��*<������5,l�n���@"��;�MWE6�b�9@����5�����?��`��a׶~��@o+�.b�U�]E�U����k>����j\�ᖨ�~u�S� �UC�#�cq�^Y�`������{Y�e�a�y�/��4UY�{�U]�fzf A! "�I���?Q
�BR�!ħBR�$ r �ǵ﮶�m��&��|�+�:wg����@A�r�'��^>s�9�����k�GLgW�\�|����?��k\�z&&u]�����W�����J�g�9|a�|a�΢� ��ݩ0�t%��Byy	~��ܽ���?w�5�������
�z�|�/?�g���?[�W;	�Ke:[�0<�M�x�V���r#)u��'s�x2��Y,��UK��j^�dҸv�,.���{oᥣ�ў
�9B4���i���Y<}��B	�X� �W� (��sY15���ı,Qu~�<ܒM-�ԃ��ýG��;�����<�=|���6n�����M�v���d��x��uLl#���"��<�s�(\�F ��}�*\P�b^�AV� @ _�"�8����{k"��d��)�������q��AlX? ��ev&9��
&7��U��5�[7�H3�� �6�(t �0�ڷ9'.r�m2�tD�p����m/�>4�	y�L�Ο��$�p���t0A [OI5ܴ34/�� o�j�Ϭ,��Q���Wɔ�. �B ă�Y
Kz�P|}�<�=z������� �9�|N�,V�;Yt�$�f ��'|���%,-�!�	����v�ţ�o�t�4��v�Io��t��� �ΓM>^c�5� �F��])���y�\�&�k%WTz�l�u�:CPJ�x&Q��ys�^9C�Z� �6K�����|<�q=�����~,.�#���	�lp�z5�F�ݗ$1)�ճ�y�&=tk��$q�a�ٮ�d����tٞ70-��a����ڦ׶��� ��ϕx2)��U��_>vva_�9�G�����'��R�G�ְ�� A�� J�Ay�ww:/V���:�^3̃�SKU�f�jT׍{H���"NKM^*�}�!������q�l���;����'���<��|�<ʫe�65y��u503Q\G5�'�F�x�Rq��Q�����rbv��=p���b�G�F1�.a$���xJ���W
��t >	�!O-�M#vVP�� c�1I���2۫N"+,���5�/w�W}������>�� 10jD�����y���"�&Ui�ʙ�����g�~��|��z�(�"c΁\�p�����ٚ���AM��G�X���}�(r�29��~d
%�ut���S�x��d9l�X��O�����ɳ������q�{Y�=*2�p.*�W�%�`����Y\p�g�mo��������x�zYS��K�,���{���G�pO��r�٬����3��/wv��UF����.����������6����1�^Ӧ}~�6�V��ƹ'&'��Ώ,�)���}�{:/�;n������3���t�����1�ſ�nܼ�b% �{$ɡ�mH�t ���q0Lb�ͭ���B��j�)! �.���WH�=�iq � ^g5+^�l2>����v�=ed��)��&)2 �*Xdꋠ�'�
8O5����^»?�kdf����{�c�ֵغa]�$���e�Q+�8fՏ6�a���̥�'ݵX�Q��熎��u�Z���1<z<*~x�f�1L�-���;8��i�2���%D��p�ŗq��ˈ��c1]�r�"�AJ��s?��4G0Й@Os�j�	3wc�ڿ��o�ѯe����+��?��_<]*���i���փ6�w�忠���1�����t�Q�P���^(V���Tiĳ�Zv���4Eh�F0=�_�!��w����ؾ�?�D���e�'<ƓG��,�t�#%���8͝��y�W�7��)�(�i�B�� X� ��������F'�11=�`$���^��� �ܡAK�r_%����U��1N�g��<�s��u��S �B����k/en�����"��S�}� ��$�hK%��ݎ�������ػgz��!>I�-�������i�?�%�>���c�۶m�b�s���A1�vh�S~.���З��jxf��7��0(�!g	��ȊX�@O���{��J���ћo�)+�F�L1�ҡ��F&Õk����|��6_�X.H� � I`�e�&�pD����ڈ��[���w��.�&�kB��d5��iI��$4ԇ3�$�O4%�_��4X� �c}/~�;o`��AL��J�H���F&2��I�>��&�d��&�ώ�v���/�W?�K1�,����>��5CeJ�ă�!,e3�%��{��{Z�'�=|�2�eje�xI˫ �l���U�&3����"��ʐ�3K�e�e+(�6� ��<mLY���3i��س{7^>�"�֠R(*��,;˺X��M�I��\��=�@�KnC̘�fVp��n1D�n-8�������ohH�k���a��u�,V,4��d�qV�X� 8���W�e�x�{�k2�q��}q� ��	��{%�r1�	?+~^v���<+Ig�Qʚ��crvF뷩���n��Z~K(fsyׅ��?3�� Gy��^�� ��]d��%�F�0��:���������Ei��g=�M �Ob�����@	��5c�K�M� P�x^O��S��u7��@�G�4&%����ZA`��j��X���_~�UY�=�=�_����s5����}���i���T�P�	����:{���!a��5�#����x��E�@e��K/bǦ8~h��+d1if%�>�3�i|u�&�D���صg/ZR͸}�&n]A>�,�׺�����8|p?���q��]�K2�l�X��39�0�M��]�7#��cv����v�Q7)��w�n{� ������4j���ܘp��<o�X�K����K���Xb�����#�b�׏cR���s�������2@��p�ui넯k�;�]����3�P{����fg�U�דk�_xŕE ����ܸ� �2�M�^3���u(�M�B�<�F�H�֎��Ӣ3�X(� |�VWC&<�;�;�ؤ�_��y�Q�F�5���_N�h���C��Ȫ���5�k��
��N�X	���m���C�5�ܴvo��`��ӷ5��X��]ZD(�ӐOg��f��-�ͨ�LL�ē��a��4����]}��J�y�n�{���F�pl�����ip�V����ذc7�f�-��0�Qx��CР�6�=�av%ё�#\-��~�B�^4X�}-m?ڸ�iF��7- ?�~=��G�d"[���|�����^� �ƍ���X⯻����'hт��I��8= O�^f��j�.�
���*:�q�K<�sN���V|����n�Ʉ-�*�<�Ǧ139#�(�jF[k;Z�;Դ��n�d����/n�J]gi9���<���f�11;���YLL� �Ha��]8���X�i'�ln\��r0�t1=���@��xUJem�R�yS&@&��-���W��.�&�zq�Z��)�O<F�ZFK"���V�b��=8r� �m݈榐���|�ܲ�Z��F�\���P��f.VBΟ?���/	<(s�䑅�	:���1[�����a�M{���S�n��9?7���ٵ�F�bQ�a�C��?��{ڰ#�F�={���4 ֘�j?��7�Q�c�m̜�牫aC��5F�b�lh������Ѧv�s%�ܺ�9e���Y�n'c��	��)�I�� �9:q|����������hK&��'��ɓb�=6����;� ��.�À|>lݶ/�|7n\�����b�%󴘶���Ţ�7������4�lp�����'I� ��B�$j!�ù.)�q�꒾�z��;��C�닕�Lf�e�����e &�F@J�?�YW6��Ba�ŷ��T]z@�d��r��|����|��T�a/�k�F�:���8[���nAѨ��;:���o�op�}�!�\�� �(d65#��fR������d�b��h�9+񐦋�b5���B�F9���xog�Ǌ���tL��> ��U]�,1�8�ǘJ ���!9����'��`����G/�/H{nC�[�g!�� ������QO�s�l���D�w�|K�C�Z7��,$�p�(�zY�A��O2�ը /�'�Y���92���?���~��4�&J�ύ{T�a���g�X>���<��&����~�� ����\z5���W ��L�NBCIW���кaQ~q����4N���`*�Z�Q|����_+�����/�d3J�����8������%��F.����rR��`��:�r�E�ܵSS㘜Wr��x������8�Է�oϹ�Ì��� ��d��31�s21	���3b�@�=�y>�q����-����jmQ%��M&$t�!��g�5���X�����޷}�$m��I�Vp��V@�y]���y�����vz6ǅ����y�ڵK<������x���u}<������sܻ�TnD�l޾�����̂L
dk�|��(�l���*K(�"{3j!TH���x}.�|4 �$�7 �ՄW�Ļϖ�sv��Z�E�8 O�q��hIj�7��p���}x�� ��܄�����P�k*�^��I�	P(d��t&�siL�;�dgW�mX�81T�"\�͗���O�IR;�����.\x/�C�7�a�p�8�Oz���#�/!Ͻ���ٍ >���-���&�F�Ԋ���y	������n��5 ��/o5�����t2[�/
Վ|�&�� ���8�"���)�<o�[�	�)�a �aS��]�j�K���VY�y\9�52S�n���f�    IDATc���m���.�NOab|KK���~ޔ��K��zj���������	,���ASss���x_�8?��y��n޾/��:v��(���4��(q�<�ܼͧ������&���v�H���BEn ��%��,����g��Us��Ma~jL �5�ͦMC8|t?��p����/�5�.ϣ�����|d�%�� sc�f06�T.#�?�37��v����@��s����l� 3@̿�M�=3c�t:�
P��?��3pk��ܜ��%�]cq�ٔcM�Vr5 �k�!�<{6�Y=pd�� Z��j�� o�Z/q�p�D�s���	�?fҸu�!�^����]qI��j�F�J����w�ͭVd���f5��W-b��M���~�Z���g�r����+��c��FB�Y���mHy�����,�Lc���_#� #˗�l���]�~_|�5f%����?�G��G˲sg/!ϵ���5D_� �{��3�!Q�N�@M��.de�`�P�#��$��;]!X��8�U����dF��k��VW�1�{�;K�Nĕ�����v&���u��%~�'U3��:��@0�6z��c�uu�ī���Z|���q箫X�}J"�lR�b����՚k֠�5s�N�u	+�K�q�R��_:c���o�%��>���,`�% �*�{���Ss
]=�J2<}��@
�B!Ii�gfw(��~v����i�T��ja$F�I��3�y���H�&~y�S�+F��f�<��s��u��yM�;$��oSzFO���U	� ȳr<v��Y��o��58��U	�/����=��y	��Ɵ�:Po�m��֭g]ِA��Ze&5�u�V�W�����nx��I���P`angN}���q�w���ţ����/��?��*V��D�Xʕ���?V�BQě��o�~������F._B>�(`�{�6���Q����r�P���=e�d\wkz�T��c�9��IW'f[Lh�,��;5�W��v�x����w�H&o\����d�>�̳�I�A��e�a�>߻�U�s�bL�>��D&�sC��� [[|����h��>�V�Y��}���h1;�H(�G˛30;=#������|�Ue+��͒�eMN~v��m��o~!��r9�X�;���=�垘�C&�x�@4�BK{�
��SK��@0,,TF�x_Ƚi��b�5�ն������V��L�j�U������Dԫ"{Id��5�7������lIav�	�_>�����ym����Ϭ��E��&b!D#A��Y���6��>�3���A{w7�mߩs�ɩ¨T);+�����{�!��N`~1�OFq��=m�Z��;vbǾCh�@�
,f
(R��&�zs�R���O�� ���h��@��J>�0��ˮ������������S2���g���
��j�ƦM[��^fy��a7M��ˈ]#�� �] �XF��c�5�rU� ��]0Q�����wK�%<�;��n��%���6��%&����99���2=�5	-�t7����9aO��9 �D�u���UV���%�����˩t~��19v��혚�az~Q:`"(�')�m��<*˹�p�w'!a��Ƙ���w.43L|����۫�Obyn� ��E_W'�m]��_;�C����Yl@( Y~���8�7S�J�\����.������9��hs�hj��vbA����������[U5vW�%N�{$-;�&[;�k�`��HƀA��;6�شo���{0њ��mp�SZv�'6�y���?8ms�o�5|��1�� O���p� �x<6����N����r��9�9X�g0��c(���&���'�O�/"�MS߆@��}۶�;o��J>��~���iY���ĪJ��,�߽w��R��!���똚�P#��#�1�߇��q<}�Dׂ;;���ށl.��.��?���l&������?FWW~����xኒ�e��2�u�lZ��4��2����)� ��3�{���#p�F�T�Ʌ���x�p*2=��S��D�F������iIVX�	�I�=bf(y���o�"ɪөZ���G�"��@�^ͱN��f^�M��::�$S ����Yܼs:]q�vK�Gٴ��0�f>Vo8�խy���*d�$��;����櫫Q�����8�?a1�~�(�!W��r���Ғ�,�@x9����XR����1I�(Q�]J��r=�{�a�����D�שi����ؾ3�d%������U�>5���y�^%������:77�	œ%/���$u�.ZjOV8�6���&V�%�����s#{k���e��� �7�����������{�F�n�gUB�l0�����ޜ���\h���۱c����ꕤ{�H�\�x�y,/-"�a�M8q�(�1��SJ��2x8:�sW���Ԝܶ�[ڰs�n��yc�/]���:S�8�w/��p�=���`�m�A���~];8�
-�fժ�w��{ZM
#��(�zb ����r[e�������g
�|]�n�1b�G��g�}&�g�<�'���x�=p�������a����k������U���<�g^�_��`	���z���޽{�v��*���N��W{�n�٤b׳"'�J#ׯ�o�ySSK(��Ռm�b����Y����� |����V�uu���C��b:�*��$3ɾ��&��5o�9 �8a ���;"��
���vw\��xR���ր9:ۨ#
�x�p ��n���%�s��Ha��}=���@s($���ނTS�������M&�?|��Ö�;T�$��5:��$��çcx�dc�S��O���f旑hm��m;���a�#S�ih�e�u�#a�VW�JNJ�(������(�Xz�U������-��??�������T��ǋ�Z{��r��ގ>x�H���kdw�X�\]\���N��kx�e�9�T�K^�@�K6c�h�g⤸3�Z�������5LO<B���lr��A�c��j��)�`�D&@�8�O%>x%o��*�rd
E��..i9��6oۮ�k`����ei�����UH�j��@�Mj��)"s�!���W�|Q:I0s䀘Z�5��}����dn��id�5�*�����|'^<���6��9����a�3��i�>�b
|��0k<�hy]��?kʳ�a,�1�V��Ɏ��V�T=�vȓݠn��A���52���CJo��t�8��C��dB,�[�Y�F�a%u;(��f���V^�j�<��˩n|^5�D���;��� �s�������d�ҧ�a�m0RL�(s�;�c�O�V�1��|�Z	{�n������R?��O�jJ���}���)ɢ{���z]��k���Q��>�呫�[\�ƭ[��o�K�ҭ��;p�.>�����7�^���u����ӓx��OT.�4�X�	�O�)�:{���Å����@�ft��Α�A���2�� �J{.�|о��l	�l�m��E��hi�#��	F��wM$�hl;v;�	��b���KŢ�g�ONЕ�q���ևQ��ku���U2��u ���M��2vKy�o޾C�C6./�����w��H
E �C����:�||~V*�G������/�����	��9�D2W�Cg�h,��X2!P�dxa�����R�hkǶm[0�fP��W�r�	4Ȍ��P�zS̹�3���Y�����b�TX�Ľ�ٷ{w�#I`�a�xq�55ZR2��γ���V�L<��8vҹ�0!�.��{�
+6����g��x���<�id+���Y�=K���Ɂ���7��ZĬ�g��b��ozO����X,�}�; o�F O	<�c��{����*[c�J0�=~��%9Ȩ�_ȣ5���Par	˅gtjV��#��s��CI�h�_���gϠR̢%�������hin�����k���kϒ?~�EÚW��oI�9Θ��x��%���F��90=�*�����n��%��4�=b�=�6eE�[Bi��-��99��P�U���<p�Wo�!�7�9Y�ro�b:�x������>��C�,��:��Նu�ML��]&-�3�뎉���+�ܮ:����o���?��52�}1� ��Hg�q��|��I�-fP�e��q��9pTx����B�H��y��h)fQb�\,�"e�5Zo������s�'FI)	.���ȴ3�����];����>`?�J#�Nfuj�x�%�:W��>��K�0?���ؼa=m��HD����=�ǂ�W�Ϝ�V0�\���$��شe;�&��B�S��_���"��g1;����,e������f�0:z����H�N�$��*�WUmp �W���a_kڣX�ۄ�p�za���� ���߉���/��~p��=�����b�� >�)aMW� <3t�ʵ*Yϐ���~z>���2UMfd���Bc �:R�CQ�����af��^)! ��d�}z#W���[�ʊ��@od�Wu���ZV�luA��;K�Λ���L��m����iW	���W��M�����M�#�s<C��"ҾW	H<��� l ��M����d#��X�@��!N�2�߳��
T���O�"�4�d<��d��=��k'��+ǰaxPA�\tVt��^�_�l���{�\)����w��{$(��0�r7&�=��h�$:��V(��K	A��b��g:I۬�p�N�ʏ|��Xy��#���N�"'�:�wU�����v;,욬�X��G ��0�U��T}�_�`bv��?Ҁz�gsEW��Ʈ�����D�ͫ�>��~��lb%������;F��V�K���z���~��Ɣ�����u��i�z��b#�+�i/Ba��t�Ξ�0��W^{M��=��E[k3�޾��g�
|����t`H������O񾆕�O"�j���?AGW���#i�h�I}E*�>�%o��il� Q_�e�zlݼI{��,��X�R��Ӓp�d���*�1;3%�7>��I��x���]ye8�kD�M#�ݚ��@j�����ǛWQ�����O	�ׄ/��#�C�N7�D���0�W�N�I��7~tt�k}7%��Τoe�����\	�8u��D�J�d�W��%C{sJ͂�����C��sjn8R�+*�U�0�m\�)���~���AgG�����|��q	��Jx���Y}�=���RW.]Vr��ͽK�����e���e��۳[��&d���FL�J�|A�9s ބGO���O>�s��������s錠�=m$u_V|$D��_���+L����?���Y�|P�8�5��30�X��ے
�~%�׫�J osT��۰g�^�[���đ@ran^M�����t�bB	L� 4Ҿ�|�\�颩f5!f�� ��hǍ�Wp�¹ ��A9t@	��¬����	�M���C�Tx�k.5�K��M�n	�&ka���W/_�a�N;WK ���aw�τ�ĉ��j�����̤��mcU��˪L�5�
jV���+9w�HD��W_}�M���@7`� �����_�N��w� �}[��*��)aE�&��:��v���@����c�c�I���3��k�!"��M[vbǞ��_�`bfQ�D~z�G��#��#����٠YFEj�B�<��Y���$���ZB�'1�HC�1^o��Y��<(���8�F����Cu_��Q��Ӈ�=r�Oі�a�n�v����E�G{U|~wF��/.�ރ��u��}>W��ܢ�AK��F2Y��Nb|r�X�lہ{���o ��U$2��z'�VH�t~،�F ����POmQ��%j��������o-�ï������>����R��\���U0�3(2�\Պ�А���4]V|���0�-]��	���k��@z�����;3�R!�Ǐ����+{�ř9�0��침L2��'��W�#D�k�*k�(ɎcCh��Bw_/׭8d�.?�|���~�`B8��4~���~�	�����8�������5��L|Nͫ _��;��|f���� Z[�زq����ҋ�п�S�<��	�	�\�m��+��*��d;E�>53-�F�������.X�0���&�Z�$��l�(6�����Ir,P76���5�n��&��c�g�=*��;�(=������c�e��M}� �ǭ�Z]�����3����ƴDI%mK�Ʀ1r�&��}�D�l/V
��TEg���;����D�>��x6�P�W�0�i� ~�;oh]����#�Y�?���AWG.^<��Ir�q�?�"6n؊x2���,�޸��?;��w��!1���طgZ�}�lz��Wi0�q�>>��K}�\�"�?����5�g/\֡^b^����5���RM��r�h�9b���b�� ����kii�7={/���=mm��l�eR6;3-F���{���� 7�S:w y����h��q�ge%q#@�Đ ~䳼��DDo�5�[�N	`�^���fż��>���d��YZ�q_H�#�J��&k$	�A<x2��?��>h��	�D�����-�c�6tuvH���s_NLOI�F��;eOU���f��}�'��rU�׈@�C�J���翙�6���sJ٨�f@6�{y~iQR��{{���H�]k4������"I�lܲ;w�����+�Q1ر�b�Y�� |�a�x6���5qUSWm��j�����n ����}�g�7�< sU�F�����Ǻi�����wrc�n�MB���-�˺uêz��/�/����ؼi�&1��"�4���)5>s�-,-b~9�\��h��d
�s�x:1�j�/c���F8���EUٚM8r� ��#K=5�W+����i����?[�l����F�d����5�u��cY�eܺz������A�2l���0�Cϵo��˷��-��#��|.7��%k�v��sh�9�=u�\�v^�w�<�8�n0L�����ݸ&�r�{��h͟`�ό3��y=Z�Q|}:{1�[��U�ĳKCJ����9��t��G >��ݻwpedW._���RcΤ}����"&��������_�k*��MYIh*���G>��A�w���\���%���p'�Ļ�eRc�9���l�����D��wn�\�8�u$"A�����xr��_����)$�u��:��^8���>�!"	�z%�F8��\Zj?�B�¦oZ�:�6��M��JFD2�=G�Ûp��Q]���:��)`>����Y���v���g�?M �$��=a_=-t���#�� |��}����sM���;���|2[���2V �P�Z�_�Q���笔���Mܒ��׀�����BC{1����S�;h4Y��5�s��N�D�[KǮ�1>�O��ē��.."�sV���d(#�d�=�W�8 O|��w��~�C�Z�x�=�Fw����Y��2Hp	R�E����kʤ�A.���_�B= ���B~:n�n�æJl���W�4�,oPɢZ� �<�R~Q ���{wn�o��->�]����Rw��e�0A}�6����ظ�����Ѡ6���`�͂��޼vL�4�e�)zd���|,���|d#z.ӹ�z���ό���Ć��؀��T�Ξ=+������'��{�1��w�|cd��&�>�Z����c�HCעPL��ѩ\�vg/\0��$��r�&�zh�TH�sd'�"��� ���yd4�)\+a�a����.��~������w����<|pO��k�d�ٷf�HB.2���Ç'?�db��]�s��>��Mt(�cqfShJP���܅�M�$��:^�v�S3���?�cu�����ՙ�.	�.�����~��PbNK�J1����-��u���>�l�U%��E {n~F>�C���탏� :}Ns��i|��W�=K�Pr�����\+�ĩ�9��0L�x5��G&�������zѐ7U]3�}�߹{��$��M$���%V|ll3�c��    IDATsӈ(ыj��30�KD8"���ԅ�<�߽���X�K���'c��pۦ�(�s^��1�dcv��=�&�]�d,.��ɘ{ɾ}�ŗ�|�͆5��"r}�h&�tZׂ��K���Ay��7�u�v<}��|vR�#�$s ���3�^!���5ԔWj�%e�'�{�^���KX���駟� K����]*y���K �M��6 O�)뚳��&��vVn����Ǜ�oc�nr?��z�%�4K{c������^�Ͽ��#j^�zqӾ��T�ԃQ���Ify�^i��S.�87�D����x��Q4��J����|N��	�(��Uƨ�[�q��5�9rDS�/�?/�j9��d����];КjaD φk�����D0F7�R���|F4$�J�l ��rf�G���>��*cͭ��qf���5f���7S�q�p�Iʽ���>澠,O��>�x�;_���-3_�rm###+r�i�g��O�w��Aeg犆�&v�-���^+��#�3��k�%��f�Rꨄ�\���w��b_oznVՆ޾~M�)��ܼ�m�@���č��ǲ�.kҹoߵ6o�B:���Ed��}� J��{�z�sH	��)�W�	�J�S�i��� �0��'a�a�g����<��kCi��#<�G��w ���H�9)�1Ƃ��J������X��DoK[�����x�DTM�ױ8.]��K�G06>' ��1��u*��(�
S�j����X;��5�{���\�"�+�/V�X���3�G��I
k$������|�;����죈����z� ��:s���N�7����/�}�J9�|���k�i��H�K�p� �~��"�2&ʦ82]cp�aʚ�H�:�&���:N>�nO^�.fI��@6��6ώcvҁC�i�FfKu�6GƎ�+׬�&?9#�#7K��lnAGW/z���߯M�2z�,Ἄ�}��On���z^c�c�X!�w�4�%Gm{EL�5�� X-��)[�T@9O�<|�� |��|ay�b�dk�:p��~���+عm#�Z�ޘn�S��xP�ρڈ�7mr�wn�[��*(2��n������Ϳ����20�ݻw�>��ۚHɦ���@�۷ok#2�1��r���n�F
k:"��k��9I0�򋏧n��_�L	9�x���c����|�u��� :p�Q��L��P0��j�P8�B�����x�:�\��G��U�0�*�z]���&SB�ZaI�%�!�#Ȧ܉�7Nc�44�������,~�w0��	v�؆uk���Sj�����է@I�ǻ���K���Ğ}�09>���nah��6�54eazV͒�kF&�F�Gsk'�)}��DM8LL~�;��f��?�g.\�;D��!�@9�q�n �ҨW�h��U�${B|��X��<�9�����=�H�Q�SF�?����&�}fEB��=��#��,0�x-P�L6\Nَ]�+
j��+LX2�RO�1�ܵ�Vp���w��i��8��;w�Q�Zv���L�c�x���`	=&7!k�E�b����>i����܈���2�պ@*'���W���!ǡ���+v19޺m3Ȱr�0y��I XxƷ��V����έ����'�Zq���giic�9�8ù��<N{�����*�o؀�1��pA�-q�.��0����Q{]���״� m����=D8U���/��}����%��a�arNv`KV�����r��z���k� ���� ������K�Mzg?�:��F�n&�ʸ�{a�ɊF�s'q`�W1�vv�P�����k���(�d\�2�[[�g���rRA�i�gfq�����+x������5��^	 g��.��V�����=w�\����¹Ӹ9rUM�&�}"(�sS�9v�\Z�#���COz&|-�Hn<�nI��"���J�Y���ŋ��%ش3�D�8��1���1�9����}BV�q�=<3��Ǐ�,QM�ј���{&��l�$���s��!c+ ��fn0��qo�ԁx2��2�_;o�K��F��A�b����϶o,��9��섊�ә��r�&��0���'�c�n�S�܅��}�J���J����Ϙ��U�!�hn��]��a�LN�czn��/�������ud7>5�9N^��V�%%)W}b�9G��l{5|��Ot'�]���
�{'a(��v�L)(����Sm8�S<p�;������+� _-ixy�,f��2J�%�N'����:Cr7o�ǝ���䕔0�&)D�DR{g�::ѿf ��v$Sm�����!I_�L�~-��"��H��1ɏ*�N�Y	h�@d���l� �h��p�����������ԩ�+}�����_��⿝����tŗ*����X/�,u��	�y�� �-RYQ�Ig�2�(e�`x]re��#u4�W.�$�y$�Ɛ�s�
ӥ��Fviٴc������|��'Y�d�,U���@�DJ2N��5���ֆxS+x��sP��Z�aP.�8��]]�rY�V0��> �i�ƃ�>���f�t��y}z �����_)�Z� �8�Z%���&lX?�Ǐ��G�ix�XX�� �r1Ξ� <?���y��N�RfHm ������ŀH�l?'�3��+��q�����f @߱4.���2�/>�%|��R��`ˀ�C�X~�g&<����L
k<��q�kgh@̀��bXI¬4��]�h��L��#�R�����p��b9�]��<�uѥ�c��G��d��i��/��5T/a��:1�����w�B�~�;,��\qSX[��H��i�s�0Vk�}���9,��LN�mhM/����%�@vyI�T�D��� $�;#�y�<�@�H}so��4���Sgd3Iй��KF�=B@M�V�ů�_��0������ޡ.��ɺ�.Pο�Q(�h^K��yB�	���lj� $K���H3�#�����fqaNS�ټ� ت���-�d�I{��#��Hj�t�b����� u�wv;���Ж-�y��Z��#���|��`U�edN0�W�j���ƕ}(�����-��7_G2ŧ}�+/���ǋ'N�رc�k`s��>�k�${�Ύv47%q��5�;s)%�1�L��EU5��sq
. �i�J'�X�nX`�׆׌{���������Ƀ�Ly؉�f����R���_0*I�o~G���>R�-~�7Y]���,a72�� xQ2b�aT57~3j�f�%�kt<b,3 ������Y �Ȱ��o �:�ͅ��<_|2Ռ��]�[7E<�����$w�~�-���먑)���əE��q�@�R�<�f���g_�ԙ�(�b�ɸ�=s
wn\G��h=�o�d1����4e�{OR���:���ٲe�*��^�ە�Ӭ3���^k�I���H O� ?���g�u�u�|���
A�|�3��sK����+��y.^�ܙ�����`��D�i��<�5�������l��Y jTԁsk��9d��@�x[+~�!ds��`��<L��k"Q��3�����@��ű�'�o�A�^��I\�-��P8�����Y�S�2�T��޲u;�n؈��%L��W�&��V���س�	��9�G��U�y��kȡ���k�5�6xw?��L�I��F ���SnȔF�ƫC��;��;g�v�
gL���E����p�����f�07���I'׫���Icvf��<��*�?)�Y���%����ͭ�H5�s��1��d�g��,�:�N��Y5b_{%�3��rNj�����7�) x��j!�0������� ��'?��r��5 O~��F������;�Xe�ƌ��˸V�c�= O�9%4d�%�Q�g�������f�|B--��(�3hM��<�1�� �l4]^B.��\.#P,�y�\�xNt�*<Ss���-�%�Q5g�!yȁ=����@��6)��˦W���d��W��Z(�F/��W �^@�T@5G��irҾ���d��T�ZA�G;vl«/����{�����_� x)2X�l��ZT��8���4�l:�=��!��d"H	��xp�̈́A���� ��wߕ4���������_x�=|~�7��7=���OV����RSP#CC�q��Is��˱{�>���'񪭤�=we~�����nr�<I����7�B:�d
�x�X&�Ғ�|y悚Y�T��x�1�$V6�8����FR-+ ~� 4�A2���M�[o�����p��)Y*nߺq:��8��%��S�\�Z��c33�s~��J��v���|�6�����1<8�M�d"G(��|�� �O��@���^;{���Ӂ���q��]5�.p����ć�,B�\/!�]�cWG3Z��hmK	�..ͩyU�l7��~�
�l���U�Ģ\G,'��=!�iƭmZSn�fIU���97T�s0�~5��5U�f�#�h���5�9��� �ޑ\e�]��7��![p^�A>.���r�pX�]}H��ꗝe$��aH=5�zP���yL�,k���u�nUpd�N�x䀴�_��W/]T�A�Z���_�����g_�q�M���o����r���@٣�06��7lTC,����d��2N���٦kL�' �qH�W�qɀ�	��N����s��1d��	�n޽�{IR�k��x���%��ǟ
���"���&�r�4x��52�_e�]eW @q�?��'�0��q�H�62ѵx����<��Қ���8^�F �*�y��2p7�� ���}M��xژ�;pй�ܸ��#�_�]��+q���|��r��d,�k��)�A9��@0"����>���7��p��Q5��=�5�ݽ���nϞ]"d��y-���ؤd��&����t��ր��`(��|^�L�izs��4ʙ���3���?WR���{��c����g�ݤL�_�ǕJjJ%�D�HO������c	�'��uX9�S�+2�1U�ZZ�b�^���u�3�=��\3�i�*���sr�X?��B%�����b̳22���>��Ԣ��1�f,���o$�$Y�ڷ����{115�OO~���wԷŸ?�0/ϵ��f}���$6nڂ���X\�brf�<��"�����ɣ�-d�f#��1i�iC* O�'M�I�eU��d������)s�q ����*�����5�j��զa"�H�
IX���Z�R�0IV�9SH�HFB�9�"���IUt3�Y�PB�V$����X������c�)�����Y�8�� �8�I�?�!�~���0@x XsS�9��|wkC�	t&�W�������Ywǟ��AN?��b�;�.������V��b��X�C��f� �#NF��l���4W��}5;�ۚ6z�/��k�j�r���˞�9$S�;K4�i��X�?�MM�����^ �L}}�i�}5im��%g	���8ufS��[�MF��&]����V�!�ˆ��J0���7uR�����j��^�%��j�a�*�b�Qtj�4j���O֨��e�B�/����_uC��&᫕0�߅}{v�W^��=;���"�5z�3�]�痭���2\�&Ԑ3 ���g6)���$�ix]�E0�0��O�V<r��_��9^�
���@%˕Jb�XD�[��1����s�dL�$����~��m�z�?�P˜r��|��3���蹽�4z6���'sp�� �Wi���Qs?/��d%8Nzv1�K�n���~�!���֊$_ ^v�*��~	~g�)�J	�����x��}U�t��c�0=�O��ö���H��H6E%!{Mi���ʜg�_�����Okz*�*��_<{����X?4�)��� �'?Z�;K�����G8w�*�so����?@����\��2�������Z�1����JC��8rh/�t"�!�]����q�)�Lu.��%�P� �&'%���F���"P�h���TWmYŦZ�
���E��1??��x6mٚ�������o��{��瑌9�J�<�"{R$��=�x�\�%�m""x(ifٯd-�-hnN�u�VU�MM�A�|!�E\��w>E:_A�޳�*vm��]�ўjQ����[Z�d���_38 9ˇ}�����`��8�� ��0��:2���9 33ؽk��\�'�ם ����Lzo\��^��̒XD�����{�{�T+��clؾm'�]�8+|$;Ƨ�1:>)�w��9k���w��щq|�����:��Ӵ�.���3�W-
h��7	��1>α��Dn��*���[|ֱ��	�6����h�%n�i�[�����l�ŲF2���o�и�Y�W�#���h�/���P���JJe�ٻ�Ihn޾��߼y�X�kW��)���Wi�L{RV�'��!\tr���y:6���9�Ͻ�v�X����S��ܲhm���d��U �My��ѫV�>�Qu�35x-y�8ٚ��{j ��&E26�I	�S�L�\��褄�k�1�7�(+:�*�$�#�����{�S��L��O~�=y�
9�9�I'�n{?LZ)�$�ojqS���l���k����`��O~�%�����1c$�7j^�\��qEkΫLHV�9�q2� �K�\c2��������3V([[�q��شy���g_��Ց����o��j��fg�Y��M[�ax�&�C��Y�;���������V�7d��P�X+}u��Vx7��4��л���Am~WQ��QE��RDxq���PH���~��\��U>~M5�S)���ı�O�i��G1!�5�:�d�&�	6���y�H��8���ä���s0�/	�� ���7�Lj+sB-�aP� �/&+�V8[̰�������Н T�|A ޏҟ��w�z ��������3��L��2�@��
�*��nF��!�`�a��6)��6d@��p씖�8���eO+�)���D&.��y�:�q�M�A�9�ϳt�.���N��&ٙ,C��Ph�0mϨ?r����a-��%h�6I��̎l�m����)Β$3G�,\(�0�ʖJ�n&�ޟ�'C�k�U���,�/�Z�>�r6�J�/��Z-8f���rJ��YX*�����ǫ/�������M�e:ܐ%&\�L<���{�#&XA�:A��/�D,�P@ٺ}���1	<����i!�)؁b`j�y�3p�ع]��(�9�>􋋲��c8P���J����-� ��]O���/�s�R��o���o|m��|�<D��±3ƨ�Iʓ�����w+{{�3(g���7j�^���c�D-��bWn������ƭ{X���S��t��L
KetZb':��Ң4Oht�*>Z�+�]�C%���h�q�KE��vmق��>��wt������~��^X���嫸��\N�:�k��s��vl݂�O����rv��E]'6B6�av!�w?���ߖV;�j�Mkg'>��Sܸu[�xЛ�FqW�3���諂C=8z��v�@��ٹ)ܻ�ݜئ�k�ҌI���9�\*���sx����)�[ܷd�M{ʽL;J�n2�l��5?d���Ϩu�>��3�[(���g(}`��Ǆ�1�b�#a���رMIQ�9��v>�k-W���?{�`g���'���2��L7�<�ū�16��x_�����!P����Q��-�mXX^���u%ݴemoi������Υ�Q��˸s�ƞ>��6mV�a!������~&x�+&J�C~Ǧ�G�\�k?x�H1r��M�ǭ�J	�>�䤪�T�Ȏ�\IIN6_��@,�āCG��o��Ǵ���SU�L��\��<��3`%����F�XW	�U�h��F�|U�� �0�M�����﫪r��c��=�l��b�:�9ׄ�7��Y��,52�&�_�j���T�=Dv�N����%����v���T��u뎼�	�Y���,8� N����%IU.�P0�x"�����eK:9)��j��!���vlGwg�����H�{�}�+����Y������:���� �����dٮ3I!c�yn�)gb�=G��K�V�    IDATϚ�ͬ����ڳa�g��<���n������_k���,1�c͆T�KƝI�9��s��f^���=���9����g?S�D�.5�H[Ն���<&��:���u(��y؈�h�\Ӫ����ܼy[�����a�64��0=��Ͼ<��.aaqY��8�riyN�����\6���>vM�<�13��|��aIhb�f4�ڥb�ϼ�٣I�CQ�Bq��uF����|�x'Nw{Cd%���$���<cx�u�!�+ 7@ȿFp�R�S(��ЪU�5]��,ĵ���rی2gʜ�ZG"�!���@/�C��A�����=�W�F"�S#��ݗى��� I�V��3fG����ܣJ`�#���z�T4��H �{ZЕ ��d9��~�Z�����_?��/N�t��3��l��ۙ�?Q,�Y�C[�����L����5�ި,�x?ȼ;mR�e[N���$�(�3�"�+�r�/�z#����f�I�(�i��w ��E��I������l��C���4F��c8���^#���sx��ˣ<�z6g|�B�GE�.������|.(j�>�;�d�i��Ü����T)�G�V1��N���p��������&^<v�M�������]R�,y���5cՙ�}\�M�u���5A*���b� %xsta��,8���M�T&eP����O�:%�!�]_z�%}7`-M����գmP�D2��ݧ�:x�r-3h���&��YF�B����i��d2�Y�Cց3�_�=ٰ~�>���<ݪ�x�\e�Ʉ�6|��Ep���\�qK,�Ʌ�K�����p�,HY�#p���Ҫ���l�E5��\Ȣ���&E�\��[���ioV��q�W�S�V��'�Ͻ8������b��%w��Fzi�����cضe�^/���k2'S���,~���x21�c'R����0Fn�����̌C((�`P"������et����E_o+���g�4P��E[��'��*����5bt	��������6{�uyM����5:�qZ�����l��
�5��y����9�fϊ[�0@Slb�����#��^3�'@ Ebcty!hg3�l��#uNC�)����,Ƨ1:���E:��\�b��Aٿ�}3D!����KJ)��~���FB� MN��U�M��~�{q��\8w�o��밶@Ϸ�8��z"D�J긷�{�0�~-bNv�i ���;�� 44<$�s��Y%��_8������H�c<֤Ë��L�͵���'{���mtl'?��5�Z�\gt��P�*�ʆ�C�8����W�Ь쳕!z�PxU�
��a����c�-�9�QdN���cL�g$������ 칟�b\= �(�i|��sp ^�S �&�g#ݑ�<�7�y�[XRU��o������`U;��	L�L�J +T6D6���ψk#X���3�4c>%2�lP��1�"_'�am?��E$��LYM�kW����DZ�^I�'d���F��\��l��g*;=�d�YbI�fl�4a�oVt	�M�n�Mڝ2��k����r�����g��1V�g<�U�ccz%�L�l}�����Hg!c 	-�u��RG'VϾR�ͳ���3+�l&�⾣u�%���d���x���>nܸ���>l޺�H��������O>������]������ڛ	�ɽX(�����H5cbnISE����!�#iB��Ux:�T(YM4����
�sV����yͪ�*�M�����od��sTd��a�ѽ���M���J"<��e'�"�����T:p��IZ
z^�@�!�%�%�!�t{��Nf§N��8�'��$��r���ZS��}�9�2��.���}&&��$��a�*aZU��Zř]T+�hJ��)���8��� �\X�����������6������4�+�v��x�@���ڭ��PuT�����?��+
h=��,9u�b)����"F.����ST���>S�5/"4���:��<I�c0��ү�\�s�C�`��^Q'�q��v�I�UZRJ����y�U����,��b�1�^���w��������_��K>A�\\��T �� |�D�H	v	�Q�JO /���|N �V\�Y��(�ӚZI ���}[M�m�1y�S:���#5�\̀���S��I��@����t��M��獶��F���y�Nw3�i��C�����P���%�f���� J O���Q�F�����Y�k��㆘V��2@���oz&��A�`H]!�{hv +���f=H�"g���҆�U��X�,�үq��{�p��󒕐����hV���I�%�"��(<�i���l��Us"*)D.��C��l%�1��kO��g2�P3�O��R,)NP����[�:�T�����f�����u�
peʹJE]Oz?3���㽏?�/��(Wsw�ҥBQ�<t���jIje���6B��'0rS�UC����`��,�C"�@OW7��4�H	S��J7F�ajbrE��{�5%��U߬��	��6l}06H���4�<h�g�v���u�D� ���g�>����(QW�u!��J|n�P&RMX\J�-gl��M��P����rEN���b�P��&����x���lmSo	e��������>��3�K0	&�>73�s��`r�)z{:q������+����'�߹u��/����I���d�#���o��Y}�_&c�ڳG�Q�2r��2���>>�z]B1�����\L�)c��{�>���7169�/N~���w`�1S$h�v�3y#��k�m߂:�MB�M.4�+����y �ML�1��->��p ����M�5��+��\o"i��/��M ]��%��Ȼ��Y��zyO��EBp�I����n�=p@ �����؛?�}]g~������}%	� ��d�"EK[�XVY��+�Te�W$N%��T*��qe~JU��#�Y�I\@p���h4�{����<���KJ��U�nt����~����<�9ϡ���s��(�,���m�� /�} ��c�;HZ�<c�L�obtL���߶��ۺ�� �.���	�m�O�v�kdm��z;z��7����Rc�1D�Yг� U��_�-�y��v[ٰo�r{nN@�Xp�T�]�tV��������d�y�YD�Oh5x�\_�I�(� �D
:y�X� ٤�*0�w��Q�
ᖞ�o\��������NB�(1��D�d$Xl�7#}��P��Hx��$`�t,��k�y���ֱ7T�ܱk��ku���v����~�mm* �E�]���ƪ�q�X�FK�����[� �H�-����!O��6��c RW��� �&����e�+�I02?_ iɅ��}	aOoZJ�z�>4���^RK�/F�c�.�$u1���.#I�N�ޖ<�ġ0 Q�ER���d�+��J9*�n���V]�����&@�3P�ޱޡa��.�֟��h.k�#�6�5�w�OJ֨�_�Y���}ӽˊ�+���ɳ�?=����Pn�q�I࣑�mݲ���T�A6���+�~ER�#�o�&R� ��5Gût�{��6w�,��y� �Qè�΅��$�a�J��-[dL0?�NL�2�xBR�`N:�T����&n}���_N[>`�����c��OY�.�Ա���M�b�|n��a
�[�RU��[s�UU6 �].h@�t���jŅ�^�h�h�FA�Xa��z�v�����?�#{��axu�V�d�.�r+�w%!��&o���Tڨ0�9wVA>��æE��`��l�0
�w�P��5U�t�1�H]���86�;AT��+�$���BR���0�Hop��!8D����z>%Qu��s����K��5��M�!��nyr��Lm�l��� �K�����+7�������CY�}FM)a4a@x&k=����O^�����Z:���]��6,M�_)���q��#O<f���v��q�ִ�/�]�˗�ڵ[���RoI�PoP�2+o�ۮ�{��cjxF_�_�f,�h���R#b�~pJ�jC<����L&N��j@B^���W�D�ݰ$,<e�&��e�1�Mp�.� ސq�K��t��&�SG�����a�TI+	a �< έ@O��vh����߸��_���a����c)��B �2�d�v^{px�֋�τ�u@+��G��4�l"��X$����R��8�z�ҌZ��6��#�ٯ���/~�s��qӎ<�}�+_S�=��/� ���VSs��n�BA�pjrT��Ǐ�a���k� <^�8-�[P23�� ���U�\�٭3\���y'�cFG�e?|P�6h�Wr���=w�瑤:J��(�pQ:t�Q{�g7����6; x��4�d�0Q%���XqY�X?�lr�I� >�[� �� ��{��)����E ��DD�'��Q�a�;�߅��f�w5Gp��������<_~?�ݦ��1𬱡�Q;�����[���M�L�h�A4�hWj���d7nݲ�{��OML����b��WmiiE�<�"x�޽6:8`�/_�3�|dw��zRq��aJ��Ԅ�V���s���;距�gmrlԲ�z� �� ^����x���&�G���x������Mo�4��}��=�����6T#��*D��ׇ��}0���������s� �5 �'��%����~��(� ����"��H��9ڃ��z~��+Ʊ�<��3�W�ɐ�>�ᒈ�i��s!w:�m��.�X�io�������֐H_��keG��a��f�&�&��#OY2��[w�7|�AN	f��,��wN�|��ikh�SJ�U�/Jh�w�o'm	��9���*��DR�$� ��2u����HZo����u�
�X[6�m��fSU��>��k N���Kau�A� P�B> }>�%���<f����H	7�1T� P���xr2��|���T�:K�lǾ�C�X�萒�T<j㹜���gM��N�����N��68������$��۷>���;��;��K�X O�dfj��'�<5����(���Ҥ>,z$�τӐ3�QYT�iwn\����lWϝ��,ܪ��(qy8;}"@0A�k(�p�n=�Ư�R����'5@"a���{��u�H$����
n.N߄���9K��S6>��<���LO[�V�Z=S�j�M>C[ �e� �+t�#�)o�G�3C/s����2�f�
��iTlp�G ���m5��� �gFS�*����fY��e��賶���=�pH|�U��夃|��A��d�z!�5�aB#��f�z0'L��f� ��x?�%t��|��y�A�dC�p%`���@��P�o�|x���]!�sU	7�U���h�i�.|y�F�a{���	�j-���u{�ݏ��g�l��?,K�7!��sa��)��AƉ�����f��+:O�l��G-3YX�֖-�V�a�҆e�I/�zH�Í����h\�V�ƍ[�hLo�.�ڕk7���V�Y�Z�{v�׎>e� �U��5TrU�/r�L�j��]�}O���K�Vm�xQE�
S�����#�i�� 5�D����c�-S�bG
���1�$�	��я��P�F"��`�L,��,�ܓ������?ȱX|�1:�H7������Z<�Y�A>����EݺpL�*iY�X�zxl��TNX{����aH����$lT��G14��;Kv{aՊ5&�� <����U���'O؍�Wm|t�;|�f�l�Z}�d�g7��m3�c�p�����V,�����Ļo�@�W ���}6w��ݼ~M���uN>��;��I�sz�HF;������-� ���1��$��g4��{�Cg�ډ���\iXSL`V�>��ٓG��׾�u�9w�^�կ�ҕ�:/���X���_���K��,��x$c�/��U�Pא��ɍ].`��nw�n@^��:�� �C,���w��0t��W����Q�=�kUxnx�M��?�%44^KB�^��#b[n�H�v��)	��y[^Z��y��V��+�.���uˬ�M�Kz�م�v�Ɯ��5��]�w؞]���'g�~j�}�n޸"������W�v���	ai�Z������1�W����W�"s/"}���	^8?Hh��^���O�� ����*u��c�M�ĕ��|��@&^/�3o7�Z��f��x�	f��C�	>��رc＿��\.T5H����\ժ@"�0��S��yz~��]�7Hn�1�7�{��p?B�Q�&��$����܋�+�G��B ��S�^\Z�����lm}C�B&�6\íH�1MM��O>m��}~|�x�X2�^%�hG�%.4�����1�	�3�-�Īc�� �I�w����b�3Y���|ځ1 #5l(��X�`�|d���-�ݲh���Q�iԫ6����V4�|6$���k���\,��P�����Iה���cMe��Ro��%��}�7\���*�����-9|,mKَ�ڣG��̎"�Hj��{m��\ݒF��_=mW��l��O�mX�'��s���/�x���/T�Y��R�J�R�^�t:�ANlP����.���;7����y/(�"h߽~�>z��;F,Y4M7�[V�M��d1n"AЕ������C.X/� b�3A�Q'r��|��~���9�	���>��F'�N������>o{8h�V�
0q��j�,2���Z�ķUs �lM��+���� ^���P�a�NE ������B���k����\@�� |7��i��$�V�,6]M$���g-Rٌ���T���c�q�x��j	�G��{�N0MG8w� ��0P#t��- ��!7��q���:0�vp��s���2��U�Ps$n ���I=겜"P��� ��T������'>V@\�(�1�] ����)5�2�l��~�K62ԧ�����V^[�\:aӣ��w��?�mJ$��n�<���h{�������z�F�'�
r��{v�M�ٰ���W�zҶNO���5�����Yg�x��,��;�l�����FI >��;�,SXջ�!�"�p]�4v��MEm�Ԙ=��n۶m�2����޳[s�tm{zrJ`�ܞ��zA� Oia~^ֆ����,@��\ޭ� �~�)f��Gk'��a~&)d��wޯ��g��!T����&yo[�&�\N@����A�Fb�|ҳ�#���a���)i[\ڰ��]�s�oʊ Oe'ӛ�\.nؽ;��
#45:���+�耘�YK0ѷU�\&�_3SSv��)���푇���kW��416�aT$��`|���CH����CO<�u�	B�S	>�<�g/�B�ZU �-�2��Q�r���lv�\���ѣ�g�o޴W_}M���%,k7��g�>!t��H\"�аޝ��P�}��ݞ�-�����������م�]ؐ����*�E�������	Cw|�[m����4�q���9�/�=?<>�����I������;w��g����	�f�ޙ�#;W{�3� d�bY��u�{�N���mx�����U�a���I��b% �����ٹ�F���A�>3Y�� x�OK���v�P��s�-Y�9T�4Lp�^��w����}�W�����}�NÂ��}<�ܡUǘ���*ͦLV�G�fn��=D"�d��8�� �����7�Jdq?���%�閉
�!�)
B�"���`d��A��u$�H�Hq�W�� xh�(��+W�v��%{�w���=s�I\^^�����\� �a����[^Ӿ�M"����L���H�5`FS9�bc��Q=Ȉ�˅F��yl�8��ι?�F�j�k_��D0��������-^]�˧?�7_Ֆ�nZ��M����D��0#��GI�����l�ս�}ѭ9=6ܓ"��=:�C\�$(��*��R�S�'���P`%H*o�	��j����Y��t�i#�y�53i�و�"��+�gV��S[F�cpP�����oO��������r��H�T�Xoϐm�K��    IDAT٥�/ x4� x��YT�	��՜��%�6e��E:y�/ݺj��S��pF��X���5�x�M�w͑�&�Ӭ�]<\s��3��lN�y��w����	U��	�Q5�:�}q�~����"��
�;����,���Sv��l����MZ�޲:,\�	M���Z�3�hB)�0�iA�:���
���/ޖ�$S.=��}���g�>h�iIh6�ҹ��[x��2��W�#�SP�!�����\�j�?:?7���:l@�F�����<n�_`!B	*lx
�h#}@�	7S���0%<	�&�a1؇�\��;��ktKh��  �5~�\�� � +>�s��[;���BU ���>�������v�h�)��p4�aܸiʧ�n+ ��.�6H�*�5#8�d�ebԦ��4����P�]�~��
k���� �ebƖVV%�ٻ����f�Ţ}���r&)������{��j�l���U�b��� X>8uN�땺xz9��IƭM�MI*O�L޲�^��u�d�֬7����f쑃{lb�Ϛ���,߱��;���lmeEZoŠѝ��U���.͇'߷뗯h=����C���:�9�P���M�LhD,냍o�i�EHFx�F�z ���Ghp��
E���Oo�I"��`z��F-��tkk�L�ϊ���;�>�����/ZF��X'34�4	֛֤��a��ˠ ��h�L%4�����>tPZ��W��'O��C���-/-��˗���mIe��ާυ4�܅�2n�"Ǣ�
;�jS��8�=��pC�������[oIj���7%�Ų-..9,�n[>�/�s䉧mn������=��i����4�5Ը�n�ݼ�n-m�4��fw����d�] ����8����9��tq�U%B��Z�b�������_���t�n0/R��:ҿO��%+���aु� ~bzFN-�Cڛ/\���dM�l���)���bM'�'mrj����kJ�6�%�7�dl��Y۷g�-�G�x�n]��D����6x��=� �%ɪ���h�&FGl߮�664�!:H��7�>s�c�_4��Kh�?�bgp)���?�l�j��O,�)��ܹ{�����?�#T�8������g������_V��s�V�I����o��0r6��8�Q�����1��8�����S�����'��"��s'�z2)����@4��3*�Av�イ�����w�>$!���Z���	��;K���'��coڍ�s�!7�S��ʪXx� ���G,���mIh�r��Cܤ�=���(���@����uls�i1� x5�ʵ�5�~��/��������o�ԓ�p�; o�Lw�ܺ��.������^����-��U�l�=����C��#�ͯ-����N��G���g:���$�.�I	}��J�* N�}�H�N�?e��Ǎ[<�g�����M
��y�!�w�k(��m�֛2KǨ<��QZ:��_M͎��khh�����-?y���ִ�W��d�ж��Q�:�Ǣ�&�r�~��<�b,$r..4�6�e�F�l�s���_��K�^,�Y��������+��.�&ADٛ��F� ,'G%��Q/�2?��^�-7���{�4�9G��Ք�ʗn�t�Q?�� ��&i%�{ƶڡ�_�y�bټ[Q�$	�s��
�~�G� ��v�,��fV924�]�
�G[Uk7�jd����4���6:�c����ɿ���xx^ /�t߼�9��{�p�s�e.<>�+(:�^���������A� ;t�����o�Ī���[%��{%\����TR@� ���c�8�tOn�� �'0�����`���hC�3׶ۧ�בDY��qNV�/n4*@��Iє�`��p隭�j��S�֛7�k-KA�)�u��dZ�>���U�U
V-䣞M�,�NZJ�.m]W���>vHvm��>e��60ԯ�e蕕5M����ޞA[+�-l�����m��-����}��+��`}��M&�`��5����vc��ERYI�����4%�UY��T�����))"��*R�fC�Y�>;�ݑjvg�������3Iip���h\��Gt���c�[�޴K��wzs���/�V��wQ��'o\�P�a-�)�X�G��p�$���3>� �k�矗��	��h��&��#~H�_�ܻk#�c�\�H�;GK�C�ܲ��e���f�r�ڑ����O��d ]G@�Z,�]���Q�41ii��e���0�/?���߷�nܼf�|�%Ԅ�J�dwn�u 5�|�R�b.]tzwH5�g���WzZΉ�!��u�6����}j��O���Y�ljK.�|�4����G�ȑ�(�w��"r�}&Ow&w6�21��
(�3&&&aR?�������7 � �~���=���{�~��l�ۘ�kP��E^P�w�7 <�!.�,��y��% ��S/Vu��ȥ�H�-�z����G����)�=?o���"
������ 9{T[��ຎ�Mؾ}{T�B�q��M'���)����o��{��q�v�u5�wZ��FFlv�N���U���������ǕDس[ �������J��>�"�����pn>��@��\:A��9V%~�va�M�����C��ޤ�$���~�+��X��I{J <k�c���w�+�N��a|>~�q�����̙3Z�Hn~��nr����縐�0��) ��,b���a��fxYhX��1g�� 3���ҕ��kG�>j7n޶KW����?�O>=�	�ʉ�TQ�W�S���|LLNڡG��x*msK��Z��
N?iC�&V����\� |1e4�)�a������|@�/�v�컦��m&����"�XU�U��\Ҳ��]��}��˿��9�#�'�6j�U�U6d!	a{���
��u����%���{֑`�Z��%�Q�#�䃥�$ؗ���@R���VQ�@��-74c}Sv��#�s�~ۨ:��|ƶ���PODX �)Z���I�S�����^��_;�7Z��ﬔ��u���-��)��JJ�O��ю-���zrݨ��u�T�ŸjT�[�}�>}�]9{ʪŢ�Rq�b��n^��\���H��{ OB�N��]ۃ� �f ����q�9��z(�֠y���=�7���4��	'�y4��z4e��m��מ��X$��r'n�H����72�J��3x���a��D��Ed�0�73J���^2k�,�,���rۚ����S���폿�m{��G��
3S�M&�vW0�B�\�L�c�����!��k�9 �P����بc��� o	�<x�sh�y�/?��\d �a�Ag����h� w�	���j����)l�����+�p�F��i�<���������ᾇ�{N$� W9𕀨�� ��ʴI�����5x4� xI�|�y`
�v�3)��8�t$�$�<�Q�Y�F���+Ƒ�^{��n[Z�c�>�T ����n9cܚ�����;�F����[M��5���H�z��E;������x����*�%ɵD8�L���]�y�~��+vweC �i�v����!��LO�E�@8j�kg4��z�zR����*�.�䎀B��&�*��s����Y_O�:�YS$�L
��ir���o�t�(i�����l`���;ד���ೞ���r����������~���63;�=6�0���b�d��wmqyI	zo��˂_��N/ ��5��&?���I3|K؃�dl���z.�qCD��|v�!��x���M��0^�=��\h�>r�n�ݰ��?����Pf�J�J�(�Vꛍr{�첇���; >խ�c;9>fO>��6��K��l�R�7����lqi�U�T��$=�{_��{B`��7��`
 u씋I,"���0��b�)$40����'�[wgmn���!9'��-��P��m������&P�t�	�w�Y�q	�;�@XIP�l@b%��:�Q����0����ߝ	 8�{�n���pq�v|b�{�I�[ss600b���q����xI�ap`U?}SL�i��.���j̼y�ake�Mݲ��{��c�rwގ���ͣ�o��Fd�g��:kS�v��Դ���ȸ �����L��H�yl�e��擄jE�����{���ꫯ����ezF2�R/�-��[04`}2��=����C��|�����;� g�PՅm�Y'~"2���u�� ��{��"�	2T ��w��=��'�|��H���)�E�Z���O�9�0�s�Z��^���/����Gj�����;{悽s�=[��$������	?sU�D�5�u�=�����f?���!�\�Pd3=6�D��|RP"�gM^�5<ɨ�‴)���P�jlc�����8�a���I1 ���c�֫�i����)L�];�^}��v��)h8��7k�=7IF%�����{�cp�§����;2#wO:b/������T�$�V�4J�|��O� ^;M�P�[4����)ߺ�z�	���*C��Q�G���H>&�u�V.��8i����zy��HA��7h�����f�����Xn<�Q����U���'��*?�� �w7l	�;AXN`#	V�I����oIg�| ���0���I�d^Z@f�Pr@/j��=��z`���Ywwp(y�� �����#�_G����Զ%��D������.{�߷���X]_'*o�vJx��*NrR�׬��+ͬXJ"���d�����o֔EZ�,��fe�6Vn���~��>��o[vl�O*  ��ũT����Qu��K�U�����$����<'h�ǧ&��5�D]`>y<A�`�f��9��S*5j�k4�h��@�� ��g����JY��98F^��')����ۛA����q�a"9� �x<�;�Y�{9P��6�.4.ˈ�<7���p7������xG���`?�����Z��S�姟�M�[o�! ��g�.�Y�ElxdP5����VϞ9o�JEz����ّ�����߳m3Sv��!i�*���fQ$�����ؽ��[KViE,����)��t��QT2���͋x3��K�a����܏u�g�I�0�O� bݤc&��dW��L��R"�}
x縘Ɗ��J��?8 �.�Nw����X�#�W�4�C���΂���l������ցg��Je�xý̽�3 �&�T�����~��Z���b��U�[ڒ�>�D�V�;�H"n�d\���T���\�8�ʰ6�Q�1�
MZ0R}���<`O>���{�c7o\S<౜3~����r��'�m�X=1e�}bo\�)9�bC�l��C�裏��ب��$��y�ɫw����6�H��z��KT����ۆ���K��Y�|{�o�a�[����(4 �
C �B��}�gם)��z�|b\H��|�B�/Lsf��=�_g���g������})'�L�CL���V��#C�վ�e�"���#�� ���؃_��px���/Ĝs��}�AK�bXs�[��F���߮ߜS��а�$?=sV�f&�^1���DI�zz�ҥv���6��u���#�>bKwn���^��k��kE�z�3�cSS�c���ݪ�D�"z�f�L˶�ĔAo�S$�������u�n><�¹��Z�|Y�����f� �r��?�� }x1˩���/�\0J��[,�}�I��� 餯oZ�ޭ�:*�>��cp�>��ψ��?�я� �~��[���ޟu��&n��
!��{H C|
	! �s�1��W_�_����O>��]�2g�._������+�����6��}�gf�����Қ�[Y�J����p��(PI���O�BOY�MZ4	�w����x�2�,�ghw/Y���:I0���}�F �������|��ݺ�����W��3k�,a��]~�����>%���G$�1�31���~����J��Z+Q7a��y���Xkզ�c���wq2d^ϭC �[�s�H� �X�w�fv��zچ''����v�F�lf�߆rf9����
�&"����:���_�����o��R����B�e�����a٘R����Q�� .1l���^ B �U���]��ݾqݪl$D3y=4~���A8��yjГ���߂m�&C�?]Yʗ2���)u�v�5H���8Ѝ����J���%����դTB�]��fv=hO~�Y�+M�2S�Z4��&$`�&|�;g <��f��N��9 o�jZe����V�ZZ1
0��n��}�;���;j�� ^�65|��y�<(�O�TcAS��ڊk��3�ф��s4sa������%ZAt}�]B��f[B �c��qp"����СC6�ef3K�=	���Hhi��T@��Pf�A���ESC���!$
<�����܄ ���q%%�C¦�j7�x��UO ����y1�g�_�wN��+Wo
��a��vJ��52T�4Ԍ恓��N��F�5HPڷ{�=��/���[�گ~�Ɨ'�
�33S�ӓ�d6i��s���t��W��ۺ��������gN��S���C66���iH�A8i��~[+�헯�ks����<�������+�5��W�	Y���F�~I ɉw,����-c6;=b�\�j���,ߕv�l:%��T*�� (�l�@�t����Z(Xo.o9�gyB!�� ���6�W|�Bú����Ԉ�۫��J����v���M͢o������y�G4b##C69=��s�e��Ȉ�H�/H�Zc�XmDlu�l7nݳ�+Voc3���bٚ��N�-�=�֗�+Ɂ�$�PՐ&iʼ xkʅ&�I���ۡ/��-S���h�w�h�8�Ǔ��f���` t꺚��d�Hp��ݻ�{�v�O��`����85�GU�	%K펦+��@���gg�۱�^WR��H������Qͫ����hCD:��橘^S��F�K��4��q�1�{eddرl^W�߈$��7�Wp��ɭ��N[�'�D��ƭ�s�>$9�)$Ģ��k=��z��q�B`�Y? �Ь������ъvrbx� <��yD.@W�߰��i����7oI2�c��\���]d�$0�c�6�>����X�RV,�r��쵍�;y�-��zQ}:F�+�4��{�ٖ��J8�$��Q윝���[g�Ψ��^ۼ�a�] ��1���^��gO}�����%�%3���oK�źZY[�t:�1:�\o�%d�J*��RQc������L#s�i�=���8=����Op�aO����O�_AH�j#���dq� ����=���2ϐt�6	M�D��܈kvь�Ήw���������.�H�[�#7V׭�x�t:��	���L���ldd\��Ŋ-���`���/e�(N*1�0�ɔ |<�+�����@��,�xrB�; <犆X��]��I
{ ����@�zUU��\Ғֲ�W.��7^�[�i�:��!����ͺ@������]qR�fbJvDʨ2�~��p~Ta���t�z�Yœ����]\�Օ���N��guD��N�HQO������m���~�\T?����m����s#�2�S���2������ś��z�j�6#���zÆ�'m��5� ��;�}՝�X�P�Pq��J>��.��r�*��m����X-1����d��\a�O�5v�1owd����5s�����E�d��W�"y��/'���ka'��g7l����ȩ�KI��F-�k{��G�l�cVn�g�Z��Alwlr�"�{MzaMc�q,�j��|. <� \`��o�׭�ذ����WUڹmھ�Gh�?��M�)�| ��&� ��f[� l�b����zt�}���1���D��8��EL$�Шs����o����`�������4 �!�h)�5$��x~4jhofѾB�g%�`m1�X��#���!��`
���5, >|. <����dR � �V����.ٻ�jWn�[��:���F4�6 /��bo�F��    IDAT9�	�Ij�5���wn�bO?�$4'�{GRJְ	�H<:�vߴ�U��Z�nkEi�b��'{�Ν=c�x����nO?�m��0>�����h�{��Xn����]�z�ʵ�X��ٟ[������k��ǟ((3���]�׼!�IK%bbF�����3_y¾��n�db��r׮߸��֓�X�\���w4����FG�u�h�\�����Kjfu���'i� �I��?��ݾݜ'�`��6at��Ц�LhF�
,~��7�1!���"P��G�Gz�ԑVy٥ 1@οs)�(����+���VQ�j�f%fh�lͲ����z,�rѪ���R**f�`�b�G�4Ep׶�63�Y{�R�Rq��qi@�����  "Vk8��KW.ڭsn#��
��c�=|�a�����{ԐxG�Ho6�zU��Èu`;f��5����r�������Ն�h*fջ��^h��v��+vXE?��i��7�n>_�Ӷl�T���2�63 �p�]�#����������A̖m����� ;�� ���T�V���� �	�sS��LnV)��������P������$�z$�.~{kOO� O�b��M�:,��鳟i�Ӷ]��Rmڭ�ۖ��b�$_ׯ�T"JUt˖i%J���_/��. 9vm�f��V^[�ӧ>���.���=+׬\*��
���-�u�.XKk�o�m�̌��N�У��fwmޙ�����Ī���&�>&���� �!f�ڿw�<ѩ�J���Kpn��ȁ��z1ρ���s a\Ӑtq�O�wǆ���k����$/��F&����g�:��?�� <�g��\q,�W+T�C��{��xY�-{Z��Z���K����XĞ:}Zs)�Y��1Ig�;e�[�j�S���䒁=�M{����Ϸ�^�F�
^�b��5 �X*m�|�b�kD�(��r7 xU����5�ɕf\3f<��B����%D�&�����$�~ɾ,��m�7����gw�oY6��P*Y����|����0�xd��I������Vs����7��I���f�ٱb�b+˫���n�W���:Q!	�3�r��MbE��T[�姿Q,O���ΩΙ��DZ%�����;���L���" ��[o��{��*�D|e�f����C�Y2��2MZhec��&L��AvB���1������DXj��� +O3Ý �� �i�`�nyN).1��C*�ʔ�|8Ymr�M=,�K�,�(�0r�79p�!MpC 4�D��0��a�VT2����{�[��ת�AGՉ��C������@0�� �j�����-��,P |��%4�5+��3�K ����}����fg�u��*��&V�MF�7��ĝ��'a�?��1��N
��8� ��p����e�����0*���)�4��a���yO��/�� ��	+J́y`��Y�" �?0Vì�4�n�4�A7�1�<�X�)��@p�4a���q��*<�L��32z�/���bUÎN���]��`���� �4�5%��5c@�MѾ���}!ӈ��-x�ɖ�.�G�ԺG���m�(�'�'��3��Duhu� _�D2#��c��sgN��Ǐ���[��_��|�K%�aZ4I�ְ��qz�W��g�������_�w�N�?�E��Ï�J��;�aQeFG�����Sb^A��s)��Ӈ�}�-��ؽ�[���Ĕ=��~���mׯ\�ّ�a����kG��{v��7�
�噘�Ɍ���;	��lF�Q�GX\w�C�]��c��rd�������k�~�5���X:���m��% hA�֋��,�3�!%J���f.߲�?�`�U�x�ʍ��ќ3�Y<�\��/��|A��t���U+�
��!�s�a���W6&b�|�N��P��;��aI���}w�F�Ye�{a͕�)Y��"֒��ɌH�r��?,�`6�)�X�{H��bq}_ZX��j#���. �j��"���nM4s/�3��r��/5��J�R$ߎ����r�r� �P>�fM ��� 8��o8�.��͝�������Xd��y>�I�.�_^Y���_>gX_������^���Ī��Y4Y��������)xFR�H?1�{��k��HR���IP!�Á��k�D�i*@7���%��w������4"/��k��23# �ۓ���1���n���.Z�Ƚ���H�r6�m���n����Ш�ݵ�{{$sU��OZ�9 xU�<pؔ�h��k�BB��+�H�B����OiaoqT�C���{�L���>4��$��gӨ��Ժ!I 6R��y]/~��yO��@���{�>k8f����ZČ��5`-786�}�gL�~���fu�O	�B 0#��L���{�Uj4N�{��r*�����A���#�P3g�!Ҳ�aJw�HIY%��D<�)�R ��Gc��#�A�Rk<�^/	M�۳B/��ڣ}%έf�uA$*IK*q������1ˤH��V-oؽ�wt�47H��ڸQ� _zQgN�NL��.Յ�n)]_~�����x&VSTL�qauK�$�R�l*q���s��'��H�TN��װS�MT{qj�!c؟��B36hc}1K�~�,Z��|2���OCS=���u�����ݏ���w��R��|����,U�p�8d}�����8�pq� I�����Rpt���,  ����=�@e�l2��AMm����QE�)Ð���c�^�+>�^S2�0��~7�Nv��i�ΤA?���`K	�&��E6[א'5�zmT��B� �?��0��hX��qDc����*E�������%7��3�֩j�]��]�J�" iW,֤�u�J+w������s_���7�a;�Mk:c����O2��1jnBj��]��x��U6D����r�8g�^��f� 7:A+���p�*Ҽ�0���;_ 7�Cpg�;��':/��ߠ3#��^׆�uT(3R��d\#�BZw�8����=���MfS��m� ^���'h��?����H�!c3�@���R+���?m���>8- O�����m ���N�SHfY\��D�*��G�<f�oݰ�o�f�L�v��i�dB�uL�d��jBkv��y�qkN6U�8`頒�w�z����f_�+�Ѓ�Z�LޱL����(��క����w����������{Yž�˗��OO+����V�5�T�+!'(�x�.�����m��`_Z�X�K�QX���1�������PK�d&'�-�DXdј\hX�覹f�8 �/2�}�+�7ج�,0��1<.����>!y.�'��~��*����
0���H.X_0��4kb�a�I1��2����-����҆���^Ml�4�΂�ZSe�ɴ|e�x�g���(Y�k֬V���&���y$�eT��c�����_����H���c��!QR�p�35���烙bh["�q��-�����AR�ܽ')L�����Qw��i��U�9Y1��I���lv*���q��7�+I�$��!�fCt�K�|\�q@t�\g�'&�ä��'\5<Ɓ3�{��7�����*�bSH �Ru����` � (��xEu��"�`��^ ��+<�o�^ֵ���c�v�v�[]/��؈��MYC�b)ۨ�lmuݖW�T��3�@rˎ��7�h�ؽ�����r�֖���,ӅF�(�3%*H#c�6�m���O���Ӳ�	۵s�:�>Y���������d�
9g(��Ȅs��j���Ğs����I��IA��s}�w�{|�u�����k�`��:���k;`����q�to��Ǝ~�|F�)�X���Cś}IS����4W�}E7�p�L�ì��n��	\��H����g�V��d��/~n��~G@�9=�j�Z��$G���=��b��7GcJ ��?��&����Ws��Ea��eѤ%syK�z��,��b%)j��d�Q0h.3~ֆ&�z��Pu �r�XU�KF5��^+i��e,�T;�y�K����]��KV�����8^#����3�O����H�v�ͦ�NbK�c0�,2cj�gOt���_��,"`��ƚ�D�Q7꒚jkK��F�i�>6d�=QKQ��o��^6��wM叏����I O�o��ϫ5�F4�_^,k���i�[dAG�& �����t,�I��&����Rv����� �L���&M��A�����c��� 7٧tKn�-�H������M�h����2u4%M�� �
d��7���_�1�\5��	v��RR�jG��%"'ɨ�*V-��֢�EXxM$��RS��А� ��*(�3q��W�l���m���N%�;��
_,�кKz���c����?Әh��m3�&E��+��������-A�=A/$��d~�� ��x�6s�h�es%��xxd6�Iw����i��6�X�9Hh��?A���P���}�}N�ln���y�v%@���kX�V��v��e;��Ih`�Y���w/%�Ě�̧�ϸ&j�������v�}RCx^��K����sv ˷�������*A�AY���l�~���>{N�=��
��?wV��L�|��A;�o����t�/���M���b�>o��0��o�B� ���s� w�b�.)��⑦E[5kU�,kZ2N��\.eE<ݳiۋ��ؘ �훷luy�;�D:��ׯ]3��9��kG����I��g`AY��m��Khv�v�  X��1�S[f��L/\Y]�l/�`I��KLi-����Q�Cr$�)+�:b����5#k�Ӗ��[B6�15�� �mQ�n9���78���JY�'.~6���.�CJ'��p���_�G��컋d�` ڕj�*�ȝ$�xL��E�,ƙ�����3�ĥ(�r�*��*e��˔ �H;�6��P�$;����3���Ҏ�
x�t���v��aǠq���N�;2�P�!V�9މ�1}/��8Or�Z^�1*�F� ��mTs�T{�`���Q���=�U�~��}J���U0'�>�<���X8~��""|E���a����w�^{��G��<~���ܓs��l���ܨ�i\��Lx �B+����Mhu���YacŪ�U��׭U))AO '��{�h�6�Ke�6=5#�1�A|���q۽}����X>��T��
�z����T�:M���vxǊ&��Zӹ㜈�k"(��_d�$E<i($b�Y��1��б�����U�����'�	��w�Į�D��rN��c⺆j����~b�"��5r�����Iɞأ�G�XR�K�j������q츝:}�6�U5��c��R�&����$�=�؁;�/Ǽ��h�-f�v�F;� �%,�����Yɨ����b�,[���[uR_���j1�9���x��tD0I� 8��9CI�!fk�Z���'��p�.\S��ȋ����:�UX�l2j�'��;�JH���wa��~�[WpU�,X-�x-�$��u�� u�$�8�� ���"���b�z�;i�A�o�SӬL\�,3�fl��g͒m�:���{�d��1���?�a��Ɖ�^*�s�����JՖ���oضm�mã�������9�7�/���c���h#�P��^뚠l�F m��L40Fc���54�1��	&�!�r�N��)�
7��K��\<�"B�>�d5 �N�f�R�Hp��j��cT�(c���J���J�Tt�{�_l��pk�U`�ؠ��3���g �ntT�ɭ;�~���J֪���[�N�$�W�:b����Ï��bb"%l�9hP|���4���Q�]�X[ۍ�.H]�-��Y�C��GH� W	S,Y��0 ��Jp	\��+���G��;����0�ؐ��O�o.��͆G@$��a�Ɉ�Q9`Ä��s�x��k,I������n���S"��5Bi0*��W��G��ڵ�Vk8�(G��@�Clt{I{��q� jF�s�vlϮY;��v��u{�WT�~���������1�;��q�W���Q��>���ܽg�L���Li�q��]�r��l��ɉ���φX�j�f�w�ڵ[���j��X�F���?���^x�E;u�^��s��R�2i�pi")�y&֩�P�z{Ӗ�&�T�P����[mtt�&��%y����Gv��Ӓ�(q�R(ƻs} P�t�y����q��H5�d�m�a�g�l،�654�FM�N� �yŔXܦ����{Kwe��5&R��!9A��!�HHV�5�P�J��$��IX����_7k4l�rr�s��C4ܿ��kD�h�r*fJ|YD� �Ɲ��H}�=AF#��'��S=��P���낻��ҮJٸ.C3}n�L���8��iW*V�X�f�l�T�;1W�j�|�;<9@�
�`�����`�3ez*��7�0��1uΊ�*�cT�b�I։iH��!�\{b���#��'z8��C����l��� ��Q,$7HFF�6{k��*�!i��1M�1S"�������x���Ao '��� �r�G9��M��Tk����������{@?���voiQ��ț���-X�#z� }����ud���8��:զ�UkT7�UusZ��1�	�#�)��ձ��1UL��-�J�����ٹK ~�����#\T�Uq�t�7��܄a;��g��������sY�z�� �I�� ��s� ���ڹi����B*�5$��:��7������Yg�>G�,U��A?�!F.!v���d�����gM������������������O�.d,�g�5�����-,j.@�D"��D^�zp@VҠ�A��4�U�;ÁF���?�	�k�NBe
���ed" �� So�Yk�3֎e�!n%�I��G�ΜF�Pq	6��y�K-��e�Hr^3��l��}����;��^�U��O`�$=��qO���D�Eec�s��UB03��'	Qbs��e[���xż�W�����o`@��Vo[�ִ*���j@���XB��o�D
離 ܱ�#�pl�4l<���[�l$�d��N���^&n�/b���c���������z��R-iw�]���A����^�4e�DdX~ ��'/�Cp��h�:��-Y�a��N�w~0�d+D��F+��H����Rш�r%Ȁ�1�e���֓���}��u�=w���X�i��z=��u[.�g1KY�N�)Y�����Kw�!��Ee�!��c���l��Y����9 \[L7,94�M�dhXu���aT%hll�-�,X��b��-�aJ-zٲm�:c?�����G�ȳ��>�H$���,�_���KZ䚘��Sĵz��;�`�iP����d���mҥ�x��`�hcC`�YQ���f�dA�7�g2B�K`F�C `M���z�`������*Cw��`�{>p����\�<���\Z+�j���'�ƍ;V-#p���%ط.a�'�te<�L{q%ݎ5pö����s�}��ݝ�_����e;����[/n��"�KⲺQ���5;��Y9���ھ�mjj�Ξ;e��e{��~�e�8�ˏ�y���r��e�d���ٳ���jUM��ys����?T z��ם�E:o=Cb^a$E�<ME���҉�|h�m�6��'3n޺j�#65>f+��b�=}꣏���O�a�lP�/���ߏO1
;Xr�d�qu�sm�P�u��԰�^nx�ۀ;�>?��]k�\���0zӭ����!�R���I2���~������Q��T	�
Oxb����۷흓[� �Y�E�%�^"\ � ItژJ�b�������*��N�fu��ۮ<--�F��"���������LC#�;�/T3���z���N2�7��
�@��k�2�V�d��uk�K�Q�Ir�g���)�ǣ�Ͻ�����NCD����*^� V+M��0>�i�,2Ҷ��a�}���H��1��A*Blp2+-���k@2��nX�s|\@pEuE����    IDAT��š	��U(�;Ʌw,����^7_dr|R�y~��7��$�Ȥe��8��d��	����+U+� �4�m�n۳g� �]�wT!.WM�S�!Ö�d�	�0��R�d4�Zp@C�m4�Z)���-FkH"I�
8q�^�Zc3�NyM8 y�޽b�I&U��8'i���w������\�9��"�Rʹ�܆N�Ĭ��ȿx�5�8�����`w�0X0h�5�����# s�	2��@`��ύ�=��,\�@2u�Z��V����:��G�Kˠ����H���T��������;�P*[��䝨n�Y�_�v�Vq1*Vu�#��$�R����5N���f������\�|Q2�r�n<(���ub)�'�fєEp�a S"i�L�R�^K���BIь���k%�}�΄A{��:��IdX�����~��	��㎩�]�����_�J
��vf p<�Kk��4�'��h�fy�o����Sեiw�,���{@:	:��k�+�V�ZuRM�iGLO�s�Ƭ��ĭ�l[�F�H^���2�+Ub(����|��D���e����p�F�	��o��N�Rx�'���S������������Xh|����6m�b�2�^{�/���Ve�	iԱ�t�O^�^���N6&��V�j��t�#��&�tS�g3��1���٢L߶�t҆���Q"��4�
��H�����a�V�(�ŋW�W��B�.�e�T�zmxbĦ&gmd`��&�(lu�l�F�/>m;�����Y�b�Z���	�\���:�Hʕ��9����d��$3��:���2���"b��.Y�ʲm,�Y�M�*,~��F��[���t�;vn��G9�Zv���*i����Yv��32qj�sO7�wZ0�y*9� ���� 9���طY�ם��^����#���,5[b'�C�8n�P��BBA����*��7�v���*���AR��1��`E�vIH`R�����LVe2��vkួ��v������<k@P��Y&��D`^�I�h��#K���6��e;vm�g���� �c����%ٱ��:k��b*�!���5���ho�uҖ�,��t���S��D�#�X>�ж>��t��q#�#b.^?�����
�l����?�t*o/���v��y�L�� ���Pj�s�{�i��`�}�g���Z.��k�/����lfz����v��i[_]��޼���Ra��X��\׫����"Tz��+�cn��K�\��z
�"�蚾�q�*2� ���z�m�r�t+&>s�ddX	!�~��H%����Y�T�j&G����F�`�>����O~j�w��֐��C��L�f��!/��axHO9�7W)II�&m�5i��&�z|4�Z�����J�~$�����T��7�G-q�NF�,C��lamH$]L	b�� Ϥ^� `Q�ذra�h�'2���u�q�G���q�A��|�
�w� Ļ��#ֿ�o�5Kr��$�?��䐘02H�*�p-|\3�b����(齸�l�L�$����܅�\Y�^'`N��2#Ê;�+K�@Mn �TMs��?=~|dT���zW�pǲ}n�\�azW���� ��LĒ�V�5������.�I@���|E$���*��cP'�sm�Ќ �2B�	� _/���w*�Z��"�gyCL.9�bI�{dfjZ?s�14i�����k����-��2��C<����昸 lhŀ�U��=�らAث�k���y�Z�8��c\3����:�.�K0O`���0z�*0���(=�n�ְ�p��%�E��R���(�c���(�<L�}�=�Y�9%I��rȫ�:�����#�r/����9�~��v�޲��$C��$lm��*�?D"$��E���ծ];llb\�/]�l�b���;�����?d4��I�#Ղa!�N�F2��v"-�\��Iw±�H܏�בS$V���U6�P�	�Xj�G��d­���5@��>��AV)���#�diV-�2�MңY�t�m�t�2��-�[�O?9�޻��U�\#b	U]��T�d�1[פ[��,��#�c�6�s����KFT�7�بy�XI$I`*��^>K<���	a�h�a�D��GR69�k�})�5��T��J�|��;gf���G���O��㱷�˽B��5��%�X�[.�o|��'�(�w�/�{�L�������Ѡ!�7D<��Î=]>��k�asW�Z*b�crĶ� l��G7@&jk������$�r�W9{M,>�s̞��Ԗ6>=k��kF��H�y�}
���)���$���˳�߅��� cl�hG�� ��Me�x7����ѿ���fc��E)��	�a�[�%+,߶X�I7 �'����<j�'b<x@ * x�W�S����� ๩��n/ �C�h�Ԅf(���^����X�<?�$ ���X%Q�zB �<�#��5���9�0u�ƪ�l��
v[</���ػ��{��q�v�;H �#PE�V�6���.JBs���Vܬ���]Mv�d�� ��Ś�� 8�] #���c�w�����Ӷ�z�>x�]�4���;�����w��������v��u���̮\��.�}<h;wn��?���g�왯�l.ekk+�$�*��"����^�_��K[��*���o��_�9^�3g�[����=}Vi�m�\�|��L^�0@Y�V�|:a�}�v윕.������4H
�ȅ�9���4	r|l���B6�`��/_��*�ڂt>5!�>�gs
	��U�U��Ib�b�`�y%�q7�D�^��M�#�g�=�g�g�c�N���."N�`Z_/����ry%xH�33```1ً}|����_��F�R�>�$3Vm�U)��%s��z�z5s�\-�͖
 ��a�����L�����,�63� \���dJ�C]| �:�MW�й�~ꛃ�\@���&g	����%��b�=p�:��s$Sŵ��6)!kHn�zM��S��:UI��������j30����`�����D����j�����+n
���p�Y[[���M�:@'נ^uN��t�!8�}��'�tE��r���	3��zz���6�ׯ��,�"�`�'�'�E,�*�����49���S8�����C����{�U�������������B���d�bT�6A�+�����ד��y$���[�|�몮6��OOw�w  �ͮ��]��
>�Az�R���%�ܐ��K�+� f?m�}�������m�9��Nq�AE�TM�k~����/�
R�����v��i\�� OYx2���`��o��8�m�5�{Y�1ϓ���.p]²�K���v�)��>S���]1��C7L���RP^#���Ai�}�Ĕ�����������^|~^�������ܚ�J3����e���ʻ=�y>_�Υd����'ϟq`�JP:342�y0j�9�͏l6�H0.�ٍ�N�ƻ|�مeɧ8�X�ѓ���:^^4sf���s*�0�Xbf~V�D._���;5ߵ�����޽Ax?�u?Z\���:���|�r/��t4]&2�[x��R��fØn�"�ţ:ü)�s ��-%-�ȹ�_ׇ%*�R��������u&�lE�W/�Q�"ꫣ;FwG��(z��X\��G~�K.�\��$��z�%��T���sT6P´���B��Xg7�ƶ`��}ض� ��8����ٱ��CEU(�dnZ0s��_��B5�T��1D ���(�Y,6�������c��'=�v|юe���~����??M �|��G�H��n�޳=}�b�#K����x��c��R��JqMHJ<�ڐ�r`�Ϩ�:b!t�b�P�e���Mܼ�%�;�x��}ؿ{�*�j%�Xԏh$�J��gO����)�9�Ȕ�����*�D[�HG'�l݉�=��70�r��]�@7>������e�h�F���S�j;��ݥ����{��ӍC�w��~-��8��*i�Ī�<|�� �S����	�*�qb�V���?��C�KJVNz{jI�#�fn�ksZ/ø � ���@����0��T�^��na�EeoN~v�=����B�a�q�=.�Nc�Q'����kn�N��BTT%[�f�gP���|�w��l�k`��:�P��61�2���p��ܼsb-��w�*(���xz����&�!�4͐%�[����^B�����ױ}|3^8��]I�Yb�~�z�CH%:���s�����q��CD�q�޷_!-gϝ��p~���bd� ��M0�Ǐ(�|&���c'O��'��@��y���N���3D�	����q��-D)D�)��M��E���Y�43J��>����`P@��-b��[���\c�0�F��JE�OƓ��gO�J"%�I+mr�VJ�=ض�K`A��n�f�]�޺��+ �D�ՆU�E�Q4��;��.�<�h,�R�xA�e<{�O=F(E��A���GҼD�ݽҥ����+��OT�Џ��@�&��_��o@k<�@2EKS�$qd��L�f��2�A�o�2�ǁ��gJr��w�)������:�nl��ݣ��Q"�j�際�$#<����G7'ĂUl<�5�"
��c���k�4��K�ʮ`�?5�,Х���yMƅGn\��lѢb j.YF(���حM�8�y��Ŋ�fMu�4�1�Ȇ�o@�Y����+;���ܫ��Į?Tp1�2l:��\�Xܑx`wVǴnlN�f�i/�ʏN<�~���DÈ�M�4����Y�j{�7$��$��ic��z��j�b��Τ|�m�ʒ�'<�$	�(�	0�.`��/�>x';�~����1,�Y9�8>"��	�X�:g7η8��͛��9{C�.�<Kkr5������e�%'7�L�\J0ύs�4ƙ+8@M	��ǝ>�dĹ�y؁�0�c'xf� �+<܇\QgB����g\���@�k��p�Ɣ`������xN����|>>��䔑���Č:˃�*.�)`�o���jW���'t I�����}��|�����n�5���H.E~Y O�Y��Q�Ɵ��o��]��C�֎{�%\^���#�Ɲ����f�����XRָq"��<�fJv�Hн�7F�b$/�R���&h;�%���s ސkD��Uv�$�3�E3;a��Z-t�¨2s����0ԗBOGLn~� ��K��Ïq��9��t$;ѝ�^�<i]PW��N��X*�k\�V����֑+W��ۏ}��`�g.W��K
����ϕ�oB�$�0iԞ��+ ~�?" ��; ߨ�r�:����ѱS����_��o��_�����[���C _*7��ُ]����g�|�=J0�� p9��C�Mބk ��/oLx��s�{���`��o?� ~�BfQ�4��Eܺ�%�&�}t�y��ߵE ��W��y-<؋\8ww>��J	�F��aǋ�*�*�%��M�wh��ضcb�.,�WtH���Ŋ�:�pC�­��{�o�a^�1i��KZ���.�[��Tn�^25Ҫ��X�D��� |93���'��k�6��i��z����غy\���t�Ql?��RZj���)v@�1ns�鳠�-���g��3H�������֣�jg?��@�+�$�9����k���wu����N���%��c��eq��'�z�X�B�h����G9_��9x�1��Wo���(׍����ޓ��͝`	�������b���^#`�s�V���KJ�}����؎�Gk��ʗ��b[�v����$B�j�Ο����eēػw?���p��������+�����-��R��>��k��_��̴\*��v�����O�-��q��u,�i�&�f���^]̀`�ɮ��:��-�Iv���#D�A�T!�C `�:Ye��.Yy�J�a{�)�h��ϧ��e�������� �HX�A����i|[&��gO'�##7�i,�/ ����t��04�9�P<*f�]�d���ކ�B��7.?-�r��5Ǯ Yx&gr��d����59P�&>&�ȹn�,x�8����+����pE��.�|��Z��5�#�/h�3E:�7�y�I�&D�#�;M-�3�6�ȴQJX�k��DP�D�f��P��T�FI ��Bvq�z�p �� �'X��;�k;�W�����h���nCd��1��k�� ���jQ]lf�d�I��trk�#�f�@!l�|f���]�r�g0D�I�vf�<���)Ɇ�k�W�&�&|B��`;�I�>����=��^_P9�q[�gͬ��g�ʞL�E �pT�1?���������kJ�&�o�Ь�&����)��$v8��d��1kUUq��_�K,V�@�h�݇[��1w�W�"�!�v�$/�;N�Lƛ���Q�Ð��s>|�������"�/>�{4�oʐ��u��gV%+��p�!�"���+T�<�y��w{��}�vI���ݡ�ǂ�+D��n�&y��vq�w����HX������1~��w13����a�mD�!����'=�;m^E���gjZ ~��q�g�5�������f^\�J�'��Q��̘^�v���"h�W�5�JHr*+f��ʅ�C��d�ז}w,�HS�w�;l"�^���N�n�
��HfJpo�Zn�?�avF��'�XЋT, _�,��G~�3gΩ�Eg�M��JM��I��Au�
%�ryץR�+��%�u������"1l۹�_{]����6i��B��q��\�~+�!O	M<��І� |k!����O=�e$|�]h������0�\x�P��Z����ޞAl߱���ƭ�x'h� ^�Pm ���4������.0.D"L�_��ۓU���@_�&��^<����h�a�e�@��:��^؍][G	�C]��ޥ�{&]��W15��R���-��E�j��Qi4��/c9�G�TU�M8щ]�`�}���rb�E��U%<C�d�E6^�)���3>�=�t ����+��Ҫ�Fr�׵q o�)P�{e˧Y��Q �W�P������S#�A�M�xG�����ؿw7=z�K."�K#�I{�7)�����dZ'-�M�����k'qq������Z\��a$k�S���l���8<��ZU�Vzß;���Q]��}qogR�>h��m,�A{;�w��{����ͺM`L����I<x�Cc[1����K_�����֕�n�G����ɽ�+�������S�Rk��1��?�kc~�96��`b�8N�:!��S�,��u�E%_��=�+	t$��ؽ��-x��>Ν?�cǎॗ�I��!-��L����[�d���t'��	ad�~�w� ��.\�*ǑXg�6����k{��6<��Tc���5$(iy[rE���l,�)C~�t\��Z��z���e��Biu����;��%�lg�]a)�1�������d�T�p�6 ��|���iW+V��ԗ�}�6�^<*���W.c%��"�a�h �JR���1��M�s�](Y�#h,l[Ih�\ShaK�,��8�Qn�^YV����$��6�w�:���8�ͬ���l�An|��Zڢ���q<���RŁqr�#���)��zEP� ���k&��a.A4� =��~T���5cQ(��Lŕ��5� 9|Z�6J���ޮ��3]�2���,<�\5xK�
z�V�:`3B|f����K�+uqM'0��׀N��N%2, ��&������e �gyZ���e�y���9���r�g@3�A���
(�i�k&�f;��iU���z.{$��>ȴ��"���lgܹ5$������F���l#�:?v��U���|CG*,X,Z ������ب����v����P0 �e�&F���Ҿ^���]��;�'v	��X. ��2�|�	��7�Lme�_�����s��|�i���w8c���X ^��R�sl�{�F&b^��%����cr��ߗ4P�oL�������
�֦��d�}��2]%��!��r�"n߻����K�"���
�W8��P���@��\&����C�c����p��}xj�i���������    IDAT?��FW|�A$�!�T�C`�5��c&כ�/pY���N�O���!��l6�"�eȿ6��l���`7O�o^�>�G�P�z��D�7�BJ9x+Y��t`疍��!�o)k��񥋗q��E,/���ۇ�cll\Ǚ3.�>]���H^q]."_*c)��R&'s���L�P;�����/`t�f�r@ 
(�r�J��\�(R���5�H�K�!��$�|�� |��?��fp�r�h�ԯ�?8y����ŷ�� *%/��� �������7Js������25�Կ
���p��L��L��������q�� -@ҿ��.͂��d]�86�a��l�<��cm�M��U-$+x�hs�4[~UI�3��4�=W����<2�*r�
�ҥ*����އ=�!�ݫ�V�Z*58���(1�r���� %j�\
���5�J;';�U�<�����؁hp��O-���s�3��6hV
ZhZy�։������|�8�=�~���x��� �*#������*�F�]��@0��n��mdnGߧ��:�&���3���j��"�p�c�ݢ��{'��kr~��5��1W8��u��;�*oi�b8��:V�z�J�%Hgr���5�㯽��B�ΜýGO�M\$8tL�e5uOXФ�Vm�F��ŉ�g-�/6�t����cx��������dW�\�FP(�<:��&b��|g	��^�����ҹ4<�����t��K�%�y��|���dQ�	��3{{��s���y\��%.\�&�_8�T��aW��/�Nط����>`�F� yv0ܹ�( �x�3 -H�ײJei��?����f,h# ��[���D]��Cl;�X���ge4[b�,�$���.)W�p�{x0<�	��(g���e|��gvP� �V��>4|>�R����2j��s�22�4ḑ�p�d�S��rn`bt�1�B��a���AO.��N�����H�%a�S>�Ѡ�}dq�Y�ɶ�\/Aj9^{�<��а���0�.�@��!�n�H%h���e��E�����,u�L��pi��T7��$�^V �:t�R��O]ŝ�*N�KG|ݽFzϒ|]ਰ�V�tHs� �w�X$n�$��s]'��ԉ�8�ҕoa��������`I�$U�� +���c�Y8:B�9U�!��	�R;]�z<��s���1i�aKd��������q���rOr�VS��<qX�3<f>�q��cb$�w�+�Hq�����
������"A��k:>�I��<���MZ���;��+l�qjg�U(���ϟQv�Y(2��J���3	<{8'+��~��8t��9^#�5�q	��}j�0�:uJ6������K�����5�tC�n\?�ʿ�=�| &����G����mg��\�$�4�:S�v�I��г��j��ٙy\�u��8���S�I1`�D�PN�Q]*��HیqC&)���>~�R��ݻ��}m~!- &���	p@5�&���b�]�%:��M��l��vo�B#�7�=���f�qr�,z[Muk�3%�
��)<x�q}s�Vv�l�*���Pg<�sxv�:��E"�û'p`����HDL���gS�x�
�޹�B�]��{�"��Y�sMw1��s�����r�R�\^��c�#�%#3�%0�y�^~]����S ��/�R�(7j�U ��� ��@�}	��� �N	M<���_����=�\|���\�.�������̉ ��� x�n� ��c�i�H�X��0��VU�h Ѡ>T1��)Ο���9tƣ�}��Lj�uCo�c�ؾm]��2�R�:���Z��>�Bz%�0�?���1��h���Z�!_�ˁ�\ka1_Ƴ��;�p���x���`[#E��lqa���+�&)��mx�$^�d�u����@�i���e�xJhxg)�,��|jF��7�H�?Y�E��6��{��7��}W��/�Ǚ3_��c1�Ά�P���v@\����ͦ�Ξ[ܹ��s3s�s�4H�i���"���n<�Ww�+<��T�ܻE��_�Ծc�S�X7�x8��{��=���1`����2̆[����_m�����r'N�ƍ{���?�}+|v� <�P�B��x"9�`�h�u�kӶ�	"댗�L	�����ĦQ|��7���U)r
uʭ���'���k,��v���L�6�ZCZ̮��z����w��\R��tw�J��FW��4H$F��ͼ�}w��ǥ�7�"d�^�Z�r�Cv>huag@��f@%4FkM͈�\Z�w}���b$쇧Yӽ/�@�%XZ�]RɄ2X 	���
��] ���ڢw#�3�?�}ͭ�F� -�`��cU�J��r�]������c�n9	<����3g���æ2���E_H�U�]6 �jP�6ڥ��Nc��3��	I�(o!@�=O���'0Ը��lj˩�%��X+&y�l�>�RI��&�j��+ G�BY���q	�E��{A� ���`�κ�9���n�5^�l螱V���$9�ag��,�(�a�c��Q��ƄDKPj�[YF1����}�D/G�
��'���::Q�O&�獰@�|/<�6훌r�l2EV�Ӫ�y�%��>B�?^��ڶÔ�sד�]�ƪ���Y�ѐ�7E��M�ht:e��7�Bn��Z������	q㼗/�&��A*��*!��kB��3@�)z�':RM�FS�}>"eG�cVk:Fz}$$�r��px����\D@н���i6$�q �B].4Fo <�W��m�-[���B��3�ļ��E;��U���뫝�q$O;�͟s�����|�p��v$��?�d�۝���&8s�?�:2�d��=�"��p��<N|��no�~����e����q�����t��.�k�� 8IrX+�����Y;2��KZU��{�/����˗���S�%��	e�ho4�I�ϧ9�Ź�U}7�S�M�G0�0��J��}�^i�W�jw�x&���]Ht� ��&*T��	VPG��(��]�D�f�P{�w�j�p��}�;�b�x7�b ��h��մ��S����!�o"=��.�A~a�!�{�Ʊ#8tp"����a���۸s�LFG7a��]f`X8v���������{$��t����,�"����O��˹��K������^F�sr5�u �ͱPr�V@E|2���׊�s���������<y���
���U��C�t�Qŵ�E�\Y8��5 ^����z1��qJ8�A_W�XsS�p��YL={��3�:��仒1���3��n^���T�S�iaa��j�v$Sr�)�J��?����
�ق��t�����m�]=�}�E�x�e��>�p�>�#�P+�2�8�L���7�U �!�BQ�az��+Ȋl0Q��L���$�'[�F-?���s�J�2��R^�5�\���;���6��ߏkW���?�W[Ά�ǂy7�J ���[�+�@��쀻��9���d��־ su�8���{.���JܱX��6��na_�ƴ�v&޵��z�sT��t�N�@��l�����?8����Kuk���S�K5|z�,>z�2��U�%����f.�Vg�������9[�� �q�����ܲ�=��s(�\�^\`�ù�0
t6�մqD9�S5��{nv� �ļg��x�,M��H�$��1Iґ_zĄ')��6X�"?���y��m��Ig��!O@����̺�e��๡Y���R��Fv� ���p�F#�ȥWPd�C�dK��fԬ�ն�2ʫ׌�4�
�B	��w'�g��1CND�BNZom���S�*;�NU�r&���%�JE0�A����`�D��gc��e(f3X��B��+_�Xq�@�|���{Q���L��ᵁdΊǓ*��y�q�wZ�2U���pHr�Z�$.0S,8��*���c�P&�˴�b��-Y���W�e������;�1��Wh�P+ڃ�=�J����x��Qdg�B�ܪ�u�����a"D�6����[���!f&��x��1"0e���L���:��,$n0=�� $_?��;��`�864P/���|(��\ۼolŢB�a�ӝD���}[��`A�"�����80)h�&�!�q��g
<�K�&T�M�~�:����T�ɂ��g<g<v*��
S��c���j��% ���ȫ�ȄD��*�0�,��?bU�=�06�n��`,�E}�=b�)]ٶm�!m(]���9'Vr�N��-�:o�˯���k�8�D��,<��d�]�7״�_~o���?�v^�'���s�g�ݵ�v}��q���p��+8�xʸ�ziM����X��ۋ��D���u�m�+�u)���7�^��ɓgx��)N�:�;�h�)���zΎ��.�yT���:*f�-����0�yϧ&q��}=���&i��W��J�.��#�$0�h�����A���`LZ殺��*[^+�a�˥��5�o�ZJ�eIG
��#�E]+��'�%^�=�0C�T9����kH�ɴ�T,�Zn	��|���Z�����11:���vk^)-KY�Ů ��CPA��,h��32�Q�=e��MNMKƵ�)�����7��0�Y�\!/c�l�	�>D;z��ŗ�����G�����J��
�b)�J)�i!�c�7����T�U
�ը���sɐ��6����!V9���3�.��.qáU�=��Є"	��<п
��Dp�6�"���nj�טr�� ��=�(���K�x���<����#潃��XP���ח��WC,� ��YTYkH�/�T�}�蛛��ȑ����ggГ-U��X�0��G��BO����6�7�Ɓ��YZ�IaE���h�n�6�ө�76��T�5]&�^Qx�
[Z�2u��ZM���+H2�����_|�Jaaz�S�4���6����^ŷ��m,3N���p��U=7�7j��;`��H?�)����ƷK\ܢ�$���z}!���?��v�w틸�:����^|��p��58�׆l���i�r`D�(�훜�1\�t~J`�����:���<z�t�� �e-:@�Ц�`�!ft��������p�xҀ�&-5=H�S"öq���
Sn4����\�J�h a�U&v�>�*d~�,-���'*
��s��f���ҕ��}n��!S_�S�Π'3�F֩�={�%Z��ȕ�,r88��J�wU:da�@����8y�@u�~�L��u���粯S��yBGf��@�չ�$����sׯ�_��Ɲ�]~v���>��G=�"�)5 ��L4UzI��Tc�!�L�Cot�w�Q�e17��ar�|�= �v��m�\�V1�W3�'giX��}���7�)JDc�� ��q��_7�%zd��Nh`1�9n�k�}� ;)���ǜ�=��s�3
��w�WA�����FC��lF�{v`����, Ⱥ�kơ�PPhe�aY��Z��&=���d*����h�n�)/��G5Ѝ0fĻ���_��������:T�J>C)�a��y�L���!�o>X I �Z�.��"+h5�4�C��;��X3��n�Ѯk�X5�զ$lɎ�Xx�^y�t��ÂW�3���,�ׄ81:�s���S����� ���u�B��J�J9ͦE(K�0��H2�6�z���X4� &u�G����;���թ�Xw���\��0׃x��=���� ��j��$�F� &]h�TC���.��n�p{���wg�_���}����qT|�.v{7�u�n� ��ﵚ �#ȴvٽX)�
��)�^�0����cܿ�˙4Ξ;�;w��ц.'�W��:۔ ����"ƙ�/����`c�G5��lrw���3�e�JS ��1���|�($  �DNvʂ�ˢ!�y]&�r��z���z��^�,IF�N�5������:�,�U,��!�2ǣV��Sݫ�b�H Q��n_��W����b�7�2v����F<�)G�\:���=:?�$~�o߆-۶���G��+鬮��i�4Ttbhh�B��ޑ�M�(O�J�!g��[w��ob��v^�~���7��5}�ya�X�"H"ʺ�B�b�U)����ۖ��_�z �ԙ��͔��U���;148���`8.D��>#�tŶ%�|ly���$8/7xn�M���c��#<�us���a;cxQ�G1�}�FG6`��q$b,-��?�+oLz3K�0�]79΋� ��v8���<������ϴD2�Ky�,-���a�Gp��K�u��gE:�)J���f �E����K���:�C�Lb-̘Ī�n^*h,��c4���zt���?����v��s�)�������O~�ޞ.��;{33S�r^�_a�,xv��h���YuǢ�j�ۘ����֖���[��zR���.N��|���]���(��,"�pmJ~OzCˮ��AZ�`@�d��"sC?�O>�W��@gO� |���ǟ��oT8�8+g���>n��jͦ �V����0���0B�ل<-龩ΧW��A�L�"$�e�W��!(k�nyE��8�44< ��!���St$���11�bl�N�ͮj���$#[/[6�Ԧ�T�X"!��97Z�QCIF�����\5L�2a��l��M�$��Ⱶ�k�2�3��Z�cϓi�WL�U@������3��fj5��k{7�m�k@�Fy[������,T�k�Ji���u	�LIeJ���M�D�J��N�j=C>����&e��P7 J��ƳZb�����%�b�C�N#�y�s$ڪ�
����8z��~�9�v,4g�3 �球���I�Ĕ�y=�z�t�$��}˰씶�88|�:^�Ϩ�h���_i:=���Zmavq�o�³�i=%6�s��̍�G+��@v���Ӳ��)��M�4�<-��"��{v����`�-�h���*��yk������ �l���d��.�j,��<�^QV&]���s�w\�4�zm9 o�\[/��&4�äR.�&s���ړj���W�{,"�(�[:��ZC�ڴ)%@c�Y�e๗��M�	vn��ȷ|V�9q�UN!|-�����o�EǴZ��
��<Pf�%4̝6��=���~�N�g�ǝ;���,<�_��X�*i1@[B���uv��io�;�ǁe]��v��R�Ϳ�z�⓿�f��c����ҁmmv�um���s�����߭?��sl�vк}�2��a���QW�ݰ2=��L�_�4ƹ/�/���˘������A��<ztl��Ѧ���)��-Yd>NGg
�[6����3I&Y0l�؉|�n+��Q���w4���G�D'L�P��aN,
M'������#'��4����,��«8������,��:�H! ��Gz��2�! "���4��?���G���s� vnF1���M'�Ai,�y�7Zr>�g���M&����}&ŷX��ɳgRv��t��u��c	>W�\�Rz3��r=��v�PB4Շ�G^®�/)���I/�{Y�}��U1�a`xC���;Q-�Q*T��� �桍_|�<%4�p����g*�Ӆ�I�#7cdxܰS��	�ض�6tǓ��ɛ 
��.4Tu�E�����Fa$�������3�|����$z��	z0�ߍ}��bt�TJy,.L��)~���UM]�M�h"�=o�Zg���	Y]����Ro`zf������Y,e�H*(V��_Ɋ�O����o`Ӷ��U(J��>�.5k������$�'�tT�֪�'�'�$[I� y|l�UL<�� <]h���#Fs�Ԃ��b���C��:|����IX�e�n�0 w-e�U��<��l{����v��΂������@���Z�ŢY�J�������b����1#��z�on|� D�Pn������r%{t��%���E5���'�L?>qJ�Itb���5c�g)��4�Qmj�Llgb1����ϲ�u%����Q�J�GP/�O{P�W�zw0@)��/�\3�m�r� �	����:7.���b*����%�kn ����    IDAT�q���-ْI��2,�6/��b��}�󓦦�e,����xX��b�&75��������j��!Uw�����������mYń}m&Uג�J42(��\6�"I�i���H��#2�'HvӀ6j�㝞�F�����%A}�U���HI�ł��;��]�I���I0����*6y���"���AV+�]�q޻,(+�����Ǹu�H7���W���FGU�R�Nʪsj�9䪼���C�8w�".\�R��n�J�Ǝ%7~jz�w	�<�2�<j�<j�R�woߊ�#��jf�cE^H,P{��	;E��u�Y��G�KG��'��&�RWok�D<�T2��r�YЮU�����|I�T��7���7W���� 1�܂Skn ����Zā�z�0��,�g�� �'����|9�Ui�ȎMȤ?Ҁ�ݭ|� �eY�x?[kc�?��< �S�I�xe��,�	�+���,��b~2��}0r&j�ۉ��=��
YN�ߴb�zʽ�+NJ���vƭ�NS��o#i��Ѷ�������y�|�s�b��\��^k���{����^�JMۤXN"���*�}�t�U��}�zn��ٕ1�F�b��t���)�����sܿ�X?g/-0>~$�'�wX0erY=��eW�r����E�R]���~rfR?#��s�n�
U�,�;��Ax�1���ʂ.�D4�4	o(���՞,�S���hp!�d'H.ÔU�W�\�_@UBݜk'��y�D���1�;A|�[�^�,����}r�R�6t���]�9>���Ǹ}㊎c��D0Q6�)���~;`��f���5QE��'-��wcb���?;q��:?Ėy�˨zBb���F6�@�B�����y�����q"�Z	�b�ڪ��C��:�� �?}qi�O?=�gӥW8�vb��Cذ�,`�r��N��_��ɸ�s`|v���<�<w��\�&���GmaFy��t"a�p^<��8c���y�A&l	U+5��,�@���쨚���@_��<���Wp��m%N�-������3�ijM�?r��B�I�WԬ2�Ť3���w���e��X��*�p%��k�m�r�JY��L�@j�l���V� x_=gl$�&�jA�5�.%c�&��J���;oIF���=��L>W�ְ���,f�s�z������}��c���ŬP��ۿ���B�L�z�����7���u��}�����_;y
��.vtu����^�s0�˫�UMoߊ���B�|~������z�q�lɰ��FO1��k���@@�}����YG�c�LZ!�x'�Nݟb�{L��V>T�%���]4��
�keij;�	��s�Z���Q;Ƒ�P(۴�hd�ٌS]����f�QL%&����H��0u�N��a�(����l߻�0�%�;�1�~�[ə�tLk�p���e,�m�"ȶ�A�o/Fݵa����m���@R���(�^�#��ŖZ��Nt�ƁFv|ƊGJv*0��#���]\Bva�_DE�RA<���۰{�tww�=�&�b����z�ڵ�^�b`���*�[6�)@`���զ������cr���"�s��ja�����&����/j;����ǟ�G�L���\�DO��I�倗������K�����~�}�~��i�s��F�H�
��I����`i��#�^B!��PЃ��ǿ�t� ݊�YTJ���*�������/���çί��x�L�zq�m��7��@�� �O��0<�/}�C���vl���
�����k707���^G���� x��Mz���o��#p���æݝ��NI#����"��-L��aa%#��z�/�lYJA�88��]���
����:r���l6	_�<�g�p��@c$jH�	|r��舎i���Y��i�8��5�j�/NB������됅Y�cǎa|l��6;x���gl'Wځ��h���Zt$��;�����vɥ�ޮ����'ο�~��3�����v���~ǽ�m�����;��]z��a:b�+E��jY�����=���Ң	��� �B#� ����|0�/.Ȓ�ȱ#�qr�ս�B6'7:�P;OF��>�;������Դk���u,.�h#  O�;m������d��d/Qz�G�f�AU���5��t%�1��X@��7݆xL�u��N1��V7�KK� ���C)���* �&r���n�G�0��}��<xW컯VFW<�}����C�M������Yc�-7���%yn�!�焅�x}���;fiJm8c��=��A[�N ޑ½�����G��dKȳ��y������b��#�X�5��+ȩ���	��	c���Mx$5��f9&����C�����ϯl��Sg�n>[y��D������T�\98�A��A���WE�k��`��+�d4
b��C|������AoG
1�v�^.`��=�Q�w����DZXY�C&�"ƨV%@�F{H&rs ȶ�C��	[���qj:�!HYLg���4f���)`q� ��/an1����6��W�D��(��op،�[�DX����M�M��� !�/�2&�4��	�8|�ת�J#k�Z O|qy
�Ҋ����.��s#'�J ύ����º{�Zy�p����u���2Q��: ������b��W��6K�v��c���,�{�v�c=�w@�mnAji�A�s;ǽ�f8vEL�M���+۬#c�*��p��E�<�����`���w�_�To��ً�u�m��o. h�t�!�dܲ7H_T�N�aj���2І,&��rV��[���9G��T?��>�i�F�N���0��8��;����թEhfjZ���Ҋ�=~�=QVF�k��c��� �m��Iisg;��M�<��J�"�$���p���#)pO��<`S*i'�6,�\�ŗ'>��Α���r-/�n����{�K�5�:��v���`;Z�K�ԛ�� x��d��E���]a5\zy�r#G*o�`��.x���OD�X��Ezaq�#�������%����"��e��Udv�t��2�O>��S���х��سk/��܁H(����cinV�]����䓏p��5x��d2���G��.�^6�,�L�Yr�����;��M��w�ũ�O�`�� �Ԡ�3�Z_�� ���Y����o���1�qWo������X9�M���''�����N0OF��&���d���ہ?������^-�V-�!��, �a�-,���?����Ug� ��	�՝3�~]6��rE�%���[��غyL�o�E���,���	>��S<}2�y.1�ԶS�y�e/I����F�C�F�	�ٵ�z�$�.��x|�=Ѫ2�)��7q��ec)xH� �:�]����I;|���� R�ד�A�^�{CQ�X px�Og�r"���y�u1�%�K����)e���hS�#%�F����{��|��Wq�ȋ�
�Y�7������D���ݞ�}q�H�]�<�n���n�I�6�h����iֈRWk5�\k���������rk�+����^��� ������'��t+Ւ�%��IFZm=��*�"��4V��-�`zC8H4����.��3���z��N�N�<���eǕ�IZ)�=e�gIuj�u=��2����T/��$��(j����;�5�p���bF΂�3S��R]]z��d�HJ��k��n�/o(���#0�iJ3��ӪK�NiWi�}��Yܽ�%��A����	=��D S���ֵ/��,���
ELb2�2f,��r��(��V�~�vT�0����ō�.��u�����)ܺw'O���JF��bUN���n�<p������b��\?���x2��@��!l�ЉD� �V�X���:"��u�w��ȈGa<n(�����t����>?�����˙2Е���=��:���Of�x�y�ؒW��s{���_EoW\/�ε�8���r%��E�CG�n��x�+ �iS?&�!c�I���H9-���Z�VU�:na%�P�8��M�L�L�c9�C�B����XX��ޣ'��Oˠ�,|���_Ŷ=�P�@#�}AT�a� +�X@�ިH>C�\���=��,5�-���ϖ��69R�\�r. ���/�ӳ 5�ӾT���gL5�W�S;}td#�g�p��%i���� ޱN���*��Xx�2t`���݅�u����5��_��/���N�P����/yɺ���p�y}Q�@=7W.x�^8M�(x^S���/�|rڄ�x|�����!W���q��]���9"��Bh���cl㰮�p$��C��r*��Q�ȄGF�S#�bB�i�h@�0�d��q��]�R%�{P�4�-Em6��F��e'�ݙ@<�>~yaQ5-��Ϭ���^ߔ��Y�z{z���-}�#Attv�T�b���a���B>��X��l��(v���[�J��>���4�nHM�&����S�zqرVÝ{4l��B�֯�h^`���=v흤�s�0�v��u��i�9T������e3�@�-�uM[��!	�f��|0*�f"!�F�i_Y�GzaFJa�j���+ w��n,�����x��������'藿��O�����ؽ���`xx�z�n^�c�����?�����i�,u"�ǌ��@k�t�z뭷t=�<}
���
���>],�\���R�	F�LV��E �����C��ʗW�w�W�t��������`�^U�v>��ѱA����o�s�6Ki�I���:���R7W(��.\�,��������B��5���H
�j*F�P�Ã*�>�����*��aRƮ�U����{O��/>���ZJ�M1ݜ[��^�?3@lҶ���$���H��G�;?��	���x�_����/�_��_��i�B�W�n�� ���0��x������S��8����ҢpX ���!\�iq�{h/�j�L�#ڗZ �Rf\�4�l;���.�:
M��ke��K<x� ^��;��a��2E��+`�Z�wCՎ�q�����\�����lWȭ9�N(+5�,fví	���:���JE����;�ȁx������X��k ��[�;ҩ]�OT�����E��ں)D��")����Jj�2,�	q�M����4��UPa��a��Ho�7ng��X��^��,�H2qN�C֔�x�ضu;*�:�(�aal <�xJ�Z,�AD���u�"��dLs)n���{��A��@�����S�
�,�*�^s=��I��H�ohF7!�ݣd���jL��E9;F>��&�("�e���&�!/���֥�(�,` ����L�oT�g,�A������05�+�p�����KW�HĄT���/S$e���NS���ùN:���ab�N\��:>��s�-.�Y��)���0�e�>��[����P��B�\̓��#"ު ��`��<C=�ש�r'a�_u�\ش�S�g��y�Ҏ�}r�o�������غe7"�6�r�޴&NZ��ALկ���kz���	wlA[k$:�49��
�Sj����S�����y�P�1��y���011"�wΉ��m��Q$�'�R���,2Kro��c4�l�c���n(�t&�H4�/�H�Vp��<�^PJ��R�+98�2^|�x���l�ܠ6͋�M�umR�����zQ�hdIҋ������HB�K�ӫ�$����Q��g��@=�0�����V��9���P�XU�tz��Kz��/�ý{w�f�u�W�t̶����1\aXzÔ}�o��L�W��es�At{� �	��]�з/~n�u�^ �?�{y<�$T����'\��x�.&vlǁ}��s��1��RE�u��Ć�q���kd��>{7�ܕ��cԫW�E�#Q�z����A���M��C3�ץ�GUЦ��l��Ec�1޺}'N�T�(��- �Ec����z��A]i����G�4����zf#0��_;'&B ���/���?+�:��%���	y�FS�r�m@�N���f�Mڠ��4��.��,�c�a�y��}�j��
�O>����@�d	ZY,c����|�"z���b�:5���h�z9I��Z>�����H�AUj9�N������;t���
��&82��2���yY��88)�{
�~�u޿O�>P�.�/|�v����%_^�������H<OPL>{���"6��i-{�����Щ$r�}1`�~Dh�Y7:XZF�g�%C�6:��W�^#�5Sj$�u�,�-�``H�E����çϐ-VT��M��~�ǻx�2��z:�8]8;N\���[ �x8��@�
��z�?�O�#�ۉ\~�0�i���CҦ��?���>f�4��a)�A����쇹�8���V-cnn�H ��������@�Hg�H}l�֔�֝Gx���0=�d�|aT����ȤP�9��I��jaanJ&��=t?���љ0V�|/F�Db1,,/������"�x�n�B�>�w�ͼB��B!���B O���@��	�� �����x#�[�G���ϡt����i�'N �k�E	�q���]���2��x: �4�Cˏ���Rο�.�� \֘�ܪ)��$����8�&x��:� :� �W2�F�l4�HpN��]���ޯ^9�8�߫\GבBn_s�y'tF����m�u�#s�L�9�<ރ��.�a�8'#�96�����skPu*���gt�\�	�]��8��΢��=.^��ئ-�������.4��k^
�T��r<Һ�3����0�S��"�0�V�,�b�Z2�v�`t�nlٵ����gi0Va�(����ew��W]!�Qoo_ǝ//�3�PoJ ~���:5��7���=ܾyK�-zYP
O�:�,~xS�M��>��Q���$\_ry etu�`מ��6���8�K��baiK��32G��SRpl�{;�D����
J<��&�~�ݳةb�+���.���7˥Z��=����Hj�o���������s��1�Gl��-��5,D���}&`E�fv@���j��`���:^X����5t�Byk�{�n\�$&��U[;\l@YA��l�����NHV��8��R7��9M��+h�Ts���u�vR!��[���%��H���%�P��q��cܺ�K+<|>�\��ξA|�~�C
~���=�i�@���l��Z�ۏ����G����}�Sa$�_V�ݽ���A E�\�f���k��o��W�[x�����������'S��M������� 7??�/Μ��̌$\t)� +�U�����n_h�t��$� t�%��Xcw o/���8��Θ�-0�R9]@[��űn�����F�=ύ���A���*��zp��M�?K+�(��9�B���;v������E\�vW��@�Z�g��(��+���7�|S��w���N�HT��|�$S�t� �n*��	RB�74�C/�(P��w��+�j�l�v���c�@?� J�D4%�YI/!6��|oz�J~oy�(+j�+�a�]c�}₮02��N8�N5������R�"YD$a�z9{������ZEұD<�B!��jx�G��ъ{5��6�W^{G���k7���I���M�@���
Ċ[��69��^���;����m�ņ�8{J=��)�0r������t/1���ޑ^Á��:�1�9�=	%AX�~. ��ѪWѝ��7^��#����#e7\�vM�o���6���I�6o݂�N,e22�X��e4���j�����?������+O)A<�H��#
	��+{qQ�m,f��xy^󅜂�8�O��۷�)#�/W�ؼy�fm؁���y\�re���"?�����p�<>��3ɽ�X�f �t+y�Tc1�a�r�FI@��qC/�ݟ�1�}�*�ΗQ�N�������޹��}�)�O/��ba���O�,f)n    IDATn0��Z�z�˞2�^���ҋ������a4kE�.\-k���-�����|��E\�|�Z~�{�Y���9���h��V�Z�Qv�s
�����o��c��q����i?�1��ߟ�K)�X�&�B�C�M6��--���0p�2-I�L� g6z�^V�I��v4*�2䮴f����bYj��������
b�~"AP+"�G�qcZ%~cbx�}�A��E`D�'<%�\����gYI;���91�=��U���#����4�~�z�0��ev{�W����u��!ǚ����}��%��Z��de�Nz��7�z5����Q�,2�H�y-�" I@��t�Xa��}�f-\�~����� ���U�M)A�Gs1]��Qg
�p=�<-��!$W[���Gc�3ۂaFL���J��Y���$'mz��E��dZ}���^R]Ȇ��e��1����O���˨eP/g���(ߒm����&���w�a���ؾ���6*���{�_4a�0����׮x�zg?���i�$��J�wb�6���+F%+�p��m��N��˽��d}u�^�e�|6���Q�afnN��k��*ad�e��c��س� z�p��E\0����,�MB�.9�l޾;�DW� ��&rEZ��QƔ��B�<H _�Q/竵R��d�/⃗����Ww��ٿ��7�U=Q�t�`ll;b�Jrq��H6�c�M��[���j46��Ҏ���.9H*�H�<��;�{7�!cCW��4N�P��/���v�#�i`�:��y=��xш0��!V�<)fh�CUmQ��d�+��F�U2�4�H�ɇ~<y:�{��an!��3XH��
��������6�-WPж��d���Ҡ}�9tZ������x|�&�'Q�h�!���A���z����@E��
&Y6kX���H��,N=D��36���f��ѰIZ3LW ۶Ohh��W_�ٳd��czfѠa~Y��-���Rkg��p�0kg��BZ���k>�[�5�7�z��_��_��Kd�A��Z@��YZ�Y��<�-�G��۽}{v����$�8u3�-r�W���ú���r�y�t��<�{w�]�u�۪����+x��W������l>'�N$�@G�K4AE(�G�����	b�12k~Z�5102���w�h~r�$���B�%���;�V)��I��f�§3K��#��g;��L��i
�9 ��7�=��i�����b��@T&���p(BF��L:�J�D��B��}4���C�v��>����A4R���,'��L6�Ǫ��n���n���W_����p��]|r�s�W������/���J�����/�-��&]4�����]�0�doi�뺉�y����\k�) o����7��H  vt~�4މ �^]�8�x�8^z���ܹ}S��|Oԣ �x�+uo܈D�KZt��/�W�ԕJ���U�<���~����G�`׎	I�8G��5r4�躼|�:v�M�e 1��y�<qm�϶������������ó�S�����Y��{�|R��0:�z�{����|y�>��T�UxS��l.]��TױE�C�#+�eW4��ݑğ�����^��UA���2�b�X)+1������Y���Op��C+Mm̔%�������k����6(j��޷��-��e���Cb?O6�F���ū7�񉳘�_T�V[���y����%V.fQ̮��_AO*����;��w�%����2�#�<���?����K�*��.�[�����״3V�4�N���/ �c2�<�d��+����R�T��u��e�����C��Q�j�	�3�,+hP���q�$mv���b�m��o2�N���AÛeڙN��i�f����N;��:9�ܾ��������ﮅ�=�ȷw�׺y��f ����:L��9�	�k ��$4�x�m�Z�qPg!S725�$=�k8/��{�$��CQ:����WT���,4I��g�R�I�*�I<� !;=;�}�$O ����i��k]
�L�B�!u�5��1 >�'�������*�ma��-ܿ~N >쫊�dǍ�\���
���v�s`z�7ab�!�z���ơ�zͨ��a|�U��I*D#����'��/a�+��d�vn�Ɓ^��S��N�������6``à�r"Z@2�|!�_�����Ġ&�w\T�KXI���;����08�Q���K����cLNqF3�EJ�^u���ۺ;h3�Q�^��Z<�p��0�
`�`~J�r��V+�]���2��� ��8qi��O^���l��B=�!ց�MHu��`�[ۦ2���
L�T;�o����� �Z��kgl��@s��q������Go�[Lv<��`
��n�G_włѾSkK�2؞Cg}�ZVu�L����
�m�F�*��:�hi9��G2Ջ@(�瓋�}�!�rx:3�糋�VZx�{�������c�,��	�{���5f�Q_�jO\��Sai�9�u��Q��A+^�1�nDb"���?~��@�UB2�@%3���(W�P��� �h8f <��jU7>���[?@(Ɠ'�p��%��e��YI^�f����]�A���
Ϊ9���BmC��]s�i_���s��Or]i��I�]U��U(x� � �&����f{?fw�	��"4��zV�P�f��vfw{�@� C޻ʛ,�Y���^!�ݣ�|V�{��{����u`49�|`^^c�cs,��ֵ-����&KaBi�N^��aBg�F�1�|�s�*UI��UL���w��7��n�{���>׀(}�5���TP���[o�W_�����ԙ��XLm�P(� �i����0sQ�L�����^�V�������6�>{L[M��'�߷s'�ܽ�k��Sx�t�JŜ����a 閡9��@T�qGG'^{�������1���� <�[������f�^�X��e=n��}�5�۳�cǎiH��.G�px��sbĨ����q|B	�|��'�9�W���@-LQ��X[�պ�3��C�Yg��P�ک���C'ӣ�psM�y���.��
�AIh�����3Lnc��p7Ȯ��3��G����h��$�`��L$}�Y��E���}���������)�q}a1��Y|r�����oق�[G�etX]Ƶ��W�O�Y�x�"�ܺ-tdxPr�&&>H2����[����W�+1s���cO&�}�𺼘K-bq--�j�s��W������8s�T�&�� o� �i�N'#v��ٍul�W��?�O����;��RV���2�D���k����՛�����f�,�Ӫ�j�̖�Xp+��`	۷���o���p�SsJb�Ȉ2y��ǵ;��ǧ�df7��nHv�ݙ�s_(ļ�2kr�I&�b����˙�V)�,��RX�$�+�8v�.^�o�U0��Wì�b�q�C�� �-g�B��.�E�E�S� �+@�n~ʧ����-��5ϔpZ��|�ZNZxVr�X�{�"p��
B�1�i��|#�Z>�$S��0"�;.�m�,-���';��v��v����+x�����濷A������)�k:�� k�io���LV���j>�����U����ù�}�e!;�hL�$;�A|6�AJU�ҭ׉k���<J_J����%�8v�� �<�g����I�i��/`-�A��@0Aww�������E�oD �3&4�:�%ZE\�	���|!�w9)�r"�q`uvn]B&5% � ��e�Tj.4<x�mp�p�ZᏵ`��}�ޢ�%��2-j�~H�����X֞z��0������VB_{-a�v#�{RMC㩅Y<QgH&ەZk�*�a�\����@4�5#B��٩�[XHaqi;v���;E0����w��������gK�Q���Ih��n�|�X6!>���{��G�� _*��c��ҽ��ʨ�!���b��N^}������l�卲AZZ��B3���桔]~W>����
�hj��_�,��H5�U�n_å�g�U����h�`C}�ص} �2[�i4�9��9Ї����}&������Cs�c���؊�������;�|��6���E�����I���GX\����<�旰��	�o|�;���KjA2��� �UZ���(56謡�:�kO���g�(f�����*%�Q�D��?���rPO������"� 毣�]���8
��JƉ�����u�l�k*��2~|���ӆ�v�
�ݺ��"M�JI1�v2�����*��:���l��ڭA7'���g��ٸl���w�������g�8�����s%gZ�v�����N=(�M-�F��eK�����^�:`J=x��m:�U�upzx��������p�]����objjF����*eDCa|���q���8�N��Dkt��ݖ�d����u#b��P*Vp��us�Y=�ޏ~�P$�㟜��̬:'�,�28���	ܺ����	j8RM /M|���/V�Xdsy͈*5����^=|��?��OƐH������lk�����,%Ly����T~ ŋ/����̼ɼ����K�w#�����Udsm�<P������c����x<1��&�a��w����SXYI�s��0��Y�����b�)���3�����3�)1#���7飍f χ�A��|�חR�+���y����z��| N�Q:�qi�"�������CL��i@��c�щp4�����C��G%��`w��������:�mt+���VV���k˾'��.H�I�|�%�|����V�#�ۉ��Nܼ~MI������jq���4s�XBH-�(3�v��+o��߿���u��e�:�	j
k�rp���J��4�,\�����9:2d��_�?��Ҿ�32����7�ˋ�)�7�� �n�G��Ґ'<Y["�g <�e8(w�U4$��~{voW�ç,f	���ewͅϯ����1<��A(�*0���6�B.��ϊ�*
�u1��?�ُ����m%q�	��H�@�����~#�bv ���#�776jȯ�#�Ikb΀K@�$,(:��& �t0�Ih�޼U1�Vq�)��W�w��f>
k�X���� g~l;?Ze�|��eU,�N�<a� <�&�4�b�Q�ty�P4������	�@�*̚�Q�߶��~O_vN5�_v�43�ͯ������Fg�M���d4����1_��8:KkF�o�$G�MY0I԰�m�s��ұ�Xh�<�xJf�o߶fiwl�NW3�}����`:���l�J�x::{��/�i&�'���XHRVJ ����&��D����GPw0}��?F)�̧1��6��B>�7��YRr����/�@��H����>c�E$Ѣ眻/Gy��s���U����) ?�� |�Q�`W+z;�Nj��몢T����G��u$���N�k Z�*^�f~xψ	H؅�QI��7r�#u��w@6�>oH ��)<|��n��<6�Ux���z��ۏ��^�����3Ӆ�&��P�4x��-�J�ZC���}O��?������������	u"i��葇b���l����s�G�B���ey_�������٧:�Fz�ѝl�@O7�z�}[�Vf��?0^��W�`腾�6���"!��nJdZ�8�f���Q�d����Q�{���bH-����$ƧR��5�r&�W���}�ex�Q�KExJ5� W�.O�Fi�������HM>���G�\�; Y�B��'
G�݃�u�qH���-򠻊D��W��0�lzE���˾��n��aL�X���+����7����XJł\i&�ce�)uUT����2X�i6�m�g��9
�S ��v}�fik �����~�����l ��5���l��d�Ȓ��W;�C{g��tH pg�[d��qP���'F0áW���K��B�޽����\�KCx�2�G���#�_� ��OD���kz��M�4��������[x��>�Ǐ�����[ӽ�������L��b}e]��<�X&� �����ax�F�@I!L<�:�M.t��]|~�WWі�¡Ç�xp��Oԕ:���Y����D�"����n\��O?=���iD[x嵣x��7]��������_��ݽW/]¥�.`ue	�d�1�8���n�{���w�����?��y�ɾnݺ�c'O`}=�% �)��-�f��|�?%Z�_��[���睮V�k�Y��J��ԥ�+�wtѩ0�뇇�,w.v��^L!�r�K�H����v|������01�����mow����y��č[�t������N�r�0�<  �:>�m��md�����ӫuE _,��Ǎ:Μ9�b�C�T�z�:�YȲ��^Ûo��ONG���/�K$ZZ�!%t"c����`rv�Kk(�٨ZCgo� <�K�]��ON��KBC0&�(�q3LJ-z�Z1���R1�����^�g~�������b�P�.%�d�o�y���o�d���,���#k�1v�ә�榄���سk���-C�r�M��9$�s�!�äWo���>8�{���GT��pe�PɂS�[�oh��]WaВ�����_�4, �y!/"J�Q>��S���ϿWr#�A9W�F�clY�3��{P��Y�DM1��	�5x�9��1�1��\���5&[zО�b��Ks�q�����ec����� f?�6�cͪ�e��*���y��Qv�FJc���H�<�Yp����tp����O�!���l���Pj>�A��1��dQ3�%ՁHL��I��5nK���4W��+w��29X�E����J�Xc��ӭ"<�`%Qr�βsv{\"������{��B8t� 2��7��5i}��s��?�8��ǡh�������:04�U�NgO	��m��Ʌf�{��1I���P��#�<�'��af�!j��ܗ��D��F0�����,y=����oM�J�3PfMS�^���H�h��Û�p��)�<w�aK'�b$�d��$_L�h2��"Z�q��qO�&�/�-Jy�)��=۹���ܒH��o>H2#ʰW�2�_X��0=� ;X���4�o�E��W����R\<����%�b�î:��2*ōB��=����	���?�y��������W}hI� �@4�* ρT�dIh����KO���ꎺW�m��ܼ�������+����K�:�ׇ��N�b��CC�XY����,���5 �;LY�<U�P�J�h��
�2�'{�
55��?�ryZԕ��q������Ԋ��u<���GS�I-cvqs��x�Cv���E��� �����+����bʭ�p��Iܹ�)��8�94Jy�k,'�2� ��At�oA<�a��>�!���5�F=�ױ�0���
����6W� ��͜ߟn!3�Bv�]���QYK8���+�v�2&�'�eZ�U5�<[�#A�"��tX������xf�|v5���Ŭ4�'�۔_����@ �6�n��S�!2ڭ�z��e���O�d�۲m�$	w��x__OK�F�X��� �����6�{��������h������/�#���#������>Ѐі�ˬ��b}eYZ�m۷���.���������8v��iSE �?�w�{O�Ï?9���I+x�>�2��މ��b���ڭ���I���s3b���ۇp$�+�o����{2�x�UL�!��§gQ+��o�nt��P��M��N7���mh��P�s��5�{��\S�s�蛘����O�(�;�~��m���7��5d�����k����O��΃1��>�$�!l�jP������������}��@1�+	2,	ןP�[���4�Ge	�t������?�!2��u��f����75Թ��t��=�9(�vau~��ED�np<ѰP    IDATר������
��W>+N�}���]�z8u�,Ξ�`B�(8��Ŋ|�%lݾSSX�x�m�Cz<���rb�h{��[G�d.�,�$�ք�ʜ��Y@����=p࠺B"7f��^]AwO�$4�C�����E��p7�E̥��pl�K�0�=����_���=�:��:�=u�,�j;ɖ]���z���y��9��d}9P�md#�������øΉ0y=v9Lw�����f�L��!E0UK�l��O]�Լ7ݪz^�Ã�xa�.t��hn#�i^*_,���C��|���gWnHZ�e�����b�+��]OV���*��� �O�CD�4i�%Y��@k�3]./�޸����K_���7�u�b�<�?��M O�e�s ��h3�\��r�Cb�I�78m�目N�3�Ǯm�(n�����<?-� gm؅T�߲B�d�d<fֈŌXv>/J_�C��I�3oB�̐榗zŰ�ԃ�g����^�pmfۛ����T���_"��w���g�3���\	뾱3'I��&�����,ѵy��a�CiI��+G%[dqř���N�0d�:h$��P4�^q��ml0��Ni�[{IWG�:�$Oy-(��+��$��"�:��?0����lJ�^��n۱K��z:+�m��h�r��I�ֆ3�`��hL���+wgv�i��p��?��Z����=�����,�D�Đ� �VDZ:��Ȓ������������zE���D!�-���g�^8-�h'Fz�P�Gjv+����ِ�]�����6�?��li�3�����wq��m��\�n��}�رc�� ��RX^ͨ�aġ���i�g�XKgQ�9N�#�ޅdW��
�ò��(��Dh��h������t���rq#_-e�Gc�����{��2���쭃����2Ճd�ے����#�V��6)`�� ��:�Y���k�+��N8q�!��¥�'��ś���_>���]�۷"�>���	T
t�S+�4YvE�[-(V���ݛ��@x�yS��Rx�葀>�Aʕ<\^�$	��"n�W�����O�J>3����F�|�m�����K�4rܨ<^��P��Y��ۉ��<��!ߺց��8�a\.؃�9��݇Dg?�����G^�^��-�E���rjJ�Xj&�/�j�l ��<��b��ƃ�#Yx�ۡ���׾&7���%�%�?��jJZ22d<t6A�&S`6$nƺg*�����Z����Z�?��?��6o��ܴ�M��y���	
3q�T��n�XL!E}��ø�衦�S�%y:�"� �e�D�j�yi%i�<�f�)7K�Rvq1�o}E �����3=3�dKB�h�����6�]{���W�Eja	�O��g�`�	{Nz���D`��c��d|Rߗ����xa�6L?�����tu��u�y���j[G�R���HR05���w�⥫���:��;F
�p��5����n��@�
���]�غs��Yɼ� ���nݹ��OƱ���{ᠺZ7���ݷ��߳��������I,��#lߵS�.ښ޸s'?���	#��p��7���_{�.]�G'>F&����P�xJ�t�y0~�F3(y��3��Sâ��,6���s���5	
B'��Q�|�J�0��~/��#��\I\N,/�"��, !�w�h��C/�ݼ��R�DT���٦�����u�^��ttw`���7Ћ�'ch�װsdX ����r��1:�����K--� �������G�^q���a���-%T��;L�fq����t�o��o�HQړ�S�D�ZGj-�k7ocrzV,!5՝�]��_������E&�ҷu�8�h]�����,�9�e�=����+]\������#�I�S4%(1\�
�8����x<1/�����z���4�s�2���-��Pϼ�":�3�6��2��+T��Z"����Ӕ_9|��VSqܓL �����yY0�������{�A4أ6�����
��{}��8n�}��ԪH�\�f�~�`�k��\z��Ѷ�,�:�b����-	M�]�Pn����f���c��o������`/z:�����	�MO������n�V��!�j�<����;Fox��gd�t܈D��{+�OI�7�rTWΉ��
D�U�!�yg�ʉ�z:�`�m�L3l�����M��?�^�� ���H�|-�Ye?[�cuE�W*�yy/�-�"�3��a�~�w�!�l�ǯ�>����xL��:	���X�-��%�'���O�WF���-�V�ؾS�DS3���ҳ�e+}�6Eo}rJ>x�lxUG�_ �tUa�)B�ׅ�n�=Vri��Laj��R3h8Jp��%N��jA�Y��F��َ����q0�jI�B�y�F>wA��X�n\�ᯗ�m�}�-�ߘx|_���hH቙\�r]RP���8�%	�q��nt�=V�mղ'����؃h�EO��KXO籶����y�/,bqy�y�D�;Iv���C[����W2��v��@,����oxKB�����CQ������g�8u�Ї�>��R�q0Sr��u�H�hr�+UO1�|H�Il��d̦fx���Ҋ'[�uF���h�{Pɮ��峸~�B^'�����ڎ��n����Ћ���-afz�º����f3�0ܬ8�Ƕ0/�*Z��f(!���9E����A���V8�,-m��x
��˘�]��'�H�s
�x����C/�#�/���|�0��尔��Da}��:�Gw���]�:,�%������G�=��X�6�R���Բ��BpW���B	Mj����Ͻ\�N� ��C�b���&��	��[�NĔ:����p�����+a�x��s�5C�i����Z��@��3�BKs���Ŋԙ���C�ؿ�U1�oR6�(���������r�G=;���@ ����ݧA@Z<^�v�)c'��y
�
�!��"X/��y=�irP�ƵL��}���*Ic�z�(��Ξ=����[�3+hmM��-)v;����Ʉ�[F�������Z:';���!������̳���C������w�"ܽ�H0���6r������JF�l����F����,N�9���Y�b߁�L��ͫWP�sAg��������;j&)�ݾMô�b�������o��n�=
�]�zM�[�1|����/]�N�"���f�ʍ[����.
��믿�7�~/_É��$Y�Pk{�Jo2��f�{���_ɶm�Ϙ�IR��B�m'�h,� ���HV���g�_�h��ĢpRBG�I��rb-5����n� ���2G���7��K&����Jm�������dSL	��5ġ�����W�f&�����h�'p�e#����J�\\\��'�Q(���֪b��qH�������,,W�(c�u9"uu�+ ���O���"l8��������Ӛˏ�/��؄�l� �wv��տсx��y��V�2�n4tp���D$�=��aϮ��0�RD,���f*���� �(���T���ɥfwj&����8�޼+�2LH��lڼFl;BjN��j��� �r�Gc��7�*uB�ig^?Vs�M[��}L�Z{�����[� sj�|k��������x��FCEJ��
��g����*V7
x8>��wI����^h;	vC2�Jؤ��G�	�Ų�43,J��"����h#�'#ώ�|7�l���r�[Ύ/��얤Wu�j��	�.�=$	_��S��&m��f�HVQ2⥏�W�3�)��r����� $M�9�5��|SG(,+d6��}v�{=��o��_�_�`h.��L�Ʀ�Xʚ���1��f]Xf���6�֓��
�IQ�J �dY��.r��3�����1d��<���^D�o\c�3�87/;Jιp�� ��R���v���s���tappX��-A'��>�?q����3�Ix�y�bFiu�(a�cB9cZ�r@����r�3X��B��v��V�	З&�-��=������V�9�|�f��˕��w��\N�RBs��	��l��@g^ܳw��Az5��U��e
����<\{$9���a�����d�Y�,�,#������{64��x����2V�60�Z�bj])�3��� ��F��]CݎDG���MI����}�6��C��l�R�G���_�����������Z�ND�m�C��D� ���tFg2Ɓ�h���eEM��\h��뉳W��V�G�s�p���H//`t���=��������2������$
�5}�r��5F��������E"�lo꯭H��5��
��\V���11����k���J�15���rZ��ө,��5������;w�T�˜?_�e�W=U�X��^�-�o\��k���� �JpW��,���mHv��iP�����*Mf^I2�Q�,ceq�J����{��n�d(8��4P�n\�8��f��,�<.���c��=��)u�s�&�WW�JC[I1Az��4k �²�X���.i��}���4���m����(�Q,��jo��n���PR���
��Mr��7�D}9��'p�5 �>0���̧q��]�.�H�ƵJkOjŝ[ND�~�D���ך�-����kp�"ۦ�E?飯��s�N�7��%�FgG�4���ܺmm�J�dA43���7�����
~�#���V|����'p��y� ��5�C!���>l������xx��<w#� 1��8����Ӄ-[���D��S�΋K��r�6�Wֱe��}q�$'�����ш�2�K)��g�h42ʖ���������mߍ�;v�ͽp�<��o�.�v�Y�����xE���4�χO&q��Z��{��{����[_��W��Ï��S`xͷX��6�7^�_��eL�3Ť�7-!7DcU�$�Wa��.`f��&o��% �t9w4[�P!�Gwnq>����'�{��n��>�x6��PRŶm"�*�CYL%����6�}� �����w�n1�O��:�bxv�X�Q�273+[9����헴��;3����t���K���_��\7n� ����P�9���=��c��]=����ki�/\<��O��"�Mi�m��>�Z+j��7�׏*ˀ!/tg����'(� >�_~�h���������q��-�.c�
^�1�\f�I��|+�����9!@�͝Yݲ���0��`��e���Y,,�<�)�V�+-��ف�T����&�173���y�UD9��� ��"�r "'#�bm����8u�2�3�=^udX�]�1�Q���7��ܷ�T�d��$��C&�,~��L�#E�<�bk^���`*�K�y���(e�4�4��� ��FŚ���#Ox+A\���e���E@���s��'2�"�*E�})��/!iE����=����$�-�	�2���|�MRΧ��E�~�\����y*���[����1\\���K)����p���M���g&�ST��;�=��MgU�s�'9�df��Չ�W.!Hj���}���DL�n�PB��%� �X��4;HV;�/���O��o��ZZ�\Ke��O�=P�*
����O�1�� ��e>n����`qA=<�R�

����$��DR���\	�k(V�
2����=�l��~��yq����z�hOD�01��'�G1���θY�O�v��ݿ�r)'��>��R�"�2k���Λ!j��q� S��.�t�����Bz='�}y%���E��f���� 'B�HK�h|��\uFw�E,���>�$��k����o�c�$4$sK(��s����۳�_��SB�᧗~��k*6|�R�m��Pe@����0��2�+|s��Vب+�Q6�*�'f��p��?`=����v�$����Ǝ��صs-	R�I�.΢Ī�X� '�h{��g1A] ��=�e�*��Ig�
����C)#�j E����z���7ֱ̥����'�j]2���{?�9���Q�ְ!?��4�J2�,�B��X���߿�U&�e�P+�=� 
�%G��/�X<��6f���h���?��B>����,*UFA���(C�M�F�<e������A�d�r���6I��QR�GzHO�?���4*���T;�}����,��2�-�Q��e�ؼA>�In��� ��aO7���{3�e*ك%��N�����bfɖ�0�)�K,(Ó���``tT`pf!�ɩ)�fr(е���Lo��1�{�b���tLu$�cRv��Ö��ٵ�Y<PV)�R-����[����8v�}|��d�J)X4P`%*--�����������2j#����k���'g4$��(���={1�Ӊ�/*y��뽽t��J���2���n��ٲn�+>95�L����A�T"�ٓ'Q�e��GtpؖRn�����#�g���>�-�����޳�v씴��3����-��hID��א�
yH� bH���=�E:W���Z=�ڛx�ko�������X[�ȁ�HKk�%��,�@��$4���� �S�L��_$�!h�C��p֌��B�lq�Qv�ܮ?|	�����qm�� 3���D�LP��S�*���%,0�d�Ii�-�Ç�-px�H-�Pͯ�ŝ�x��K
l������#�����$�BF��(���?^^\2�8K&�e�3��e���� �F�i~��erzF]�l�����լ`h�FF������~%f�ҥK����Oc�d[�/�bd��UD#>=�2���;b9ĺ4?'��0��dR���\.�{*udry��|������7�A��d0 ز�*�kN�5@�{�[GF����F�A�q9�����_N�q��L�ͫ�Wb�(�*J��2N؃�|�M4J9��=���V�բ��@(�:ش+-��L�&础4�'Μ��3��QD��
�$��"��, �4J^3�D[#gF�c߯ཌ��� a�e���[����4,H�:6.sd��\z���D�������uͭ"MC�d��Mg��g�H���5��_,<;���نg���T3չ^5�~>�Y[,��O�����`��Cγgԗgٛǿ���������d�M�IW.OVא���3J	)E����p���:-��Pe�N��=Y�������NZ�!��"��E��{w|�a�'c�Q���J#�tt������g.e5�3(���7�!љ�Y���u�&[�Q,VTh�L�}���� ����i��R���b�x��#��?��A��k���3'��T@���c-�
���:w9#A4�3t��)\ȧ,�sy��v�"����?�-��Gg�Z#��Ķ-��C��|������+��vcEνޤ��5����cR��U�����*vb-�[�˖��d�KK,������l��g-ҒD G(ю���ݮ�E�����yy�|���9���	�9��ѧW~�T��T����w#��B8�P�!��}�J%�Q�e��0Xd�m �L��CE��*Z}n��.�O�ᓏ~���it&�lmAoG'��a�;�ݕ���<V�Sr���%�:�F�)�w9���]��&еD.T^0��]]hmo��딮�@f���@ �����j�3�]\�z���m;�����6X��9t��Il�p�ϕ����榰�4�R.��An~���A-�J���!�6��L��J%ߖ
�S3&�Gjo�Ԙd�� �ɕ$��lLEL]���kȓ2#����Q�g� 9�Nr1R5&�P�ЦeƏhYTj#V����3������� ���F��iĴ[U�>��)`���s �{��C��ǫ�u���H}C#٢�3J<~���U����]G)7�x�w���$��'��v8�9�X���Z��r��G�ƛG��^��|t���KhKD���ёL`��{�$�Ʊ������ב)��o�7�����N�8a�t�i1�����}scH�&����    IDAT�k��tw���u�<����)U�r�2>1���dg�wI�u���;hO���JJ� ���[N�$�!�#xq9��wưu�vlٲ�s8{�&'ưup ݝI�v%���r��gMh��$��,����)d�&����k�����\�!�?<[���h-�0ţYk���y���� w����W�Ǽ6�p3��tKz�+B��8�
�!0*��o�2�	5��N������B��B�V�V��-pj��^%ͱ�+#�`0�ExX<�ŕe���3ڍo��*z��q��'���%�z+;J+��g�Fx0��:�7Lp���}{�K����!���!�7��{����$}��%+\Swn����<l���T��1<��}�=�|��\Ǉ�>@�� 6@ɿHdC- �j�5�Je��>͎����"�cuq�OĈ��HZj��ѧT�Mmv�k�b���z��]\�tCLy8���b@�%ճ֋�6�uc�)�6����w�nl�;UO�*�E�~��R�"O��l�n������Q�k(���A}��>���~�bz	�/_�ԓǒ~�Z�q(����3�V�,� >O"�!��'��ǧ/��O�`����(v���Y\���҃�b,?{��^d����5��=C$��u�[y*4��4EO<ɢ:\$rxF	�7$�$ya'��\6:��O��Vc �I�e��rR�I��$��q0��í�(�y"�JEuf���%mrѱ�w6m7���{��+�擔�����}�96�>�\W���HN7�E�?H.�{��g�&��� !Yo��8<:��o�<C);<:�؝Q��3r����$9�ᰞYv�
��f��>/:;��1e��פ�+|jyE�:HQ�444*�drrJ2>�m흲�d�i�����c�gZ�a8�2�*��ꒌ��p?�v���7��\�� �<���l�T�b#W�,0*�4�}Rx� ���宣T��ݯ��~G'?�=��?��d�!/�۰k�,�i����mLM�k�Q2p{Rg%�����Z�BE"1�s_���ս���!�ݻ��\�h+�L�<\Y�����W7�����Kv K�Kt�`h�vt����!�+���XxS�P�n�������xG�t,��m��[V�������g����F񥲃��� x�rY��V�ޖ��G�����r8��
T,�ta5��׃�X[�������{������&&i���v���3�j9'�N^�_�yJM�Q��v�1�7Q�H��L�k W(jB�m^���6�"_�&DP����6�l��.�`faI%�^}���M-\����C�p7��u�K�Tr��P:Se�k���H�vn5���='�m1��F����Q��U�ϭ/��U���5��R/�ꖬ9����,�+鍇�,��@�����hGwg"��j�7�x�hIe1�*�8क़j�5;%]2Qp�y|V�U!��{~cl� �V���k���A:)���xdq��.�+�����0<���=h8=x4>���I��x��<8��v1���;&���e+�0El�S˃��r��������4k�����}{���K�����kPOW;^=�"��G*��K��$�6�z���`l��K�#�w�?�� ��ǎcvz�51�/�݃��8f�FzyV�۶�`��m��=���T��X�K����$�=Q H�� FwoA����W��b��[�"v��qäm7���U�ON�Fsiyk��l݁�A�����铘�������]ho�#����pg�'5�����q��edU�%y���ƛ�W���>���ix��>�N�ז)R���gkI˄�)�U�ϲS'¹
;h�=�4��ʂ��b0�@<"W*v��s��Y^Ffi	��kT.K��!C���CK[oi�R�.P�����u�;R*�a�H7���Q�ޱ��YL�=F��H5�Hd��b��=�k�cA�#�LiM$Z�o�^ه2@*57�Ϯ��{�s��l\�R=��,��5}~�^����m�6�}~�">9sZ{�f*�ސav��qXl�����׿��4��$Y��!A�(�Fy�E".,,-czf^����>�z[,y$����u���W� ��c���+���@g'�Ev���.~��2#�m꘴$;�٪9��}�>WW��̂_�~��BvUz�| ��_�LDΕ�>����:���;�m��p���L5�
�u��69W��?s�
>��<�5�(e������&'�H/���x�mԾS���H1�����$Y�h�l3._,��ř7�A6܀ak.�f�ej�֞������1��(�88?��A�r:��*�S��y�Rϡh�2�����@�S�Μ�tg�;��g�m��NC�?�7|qp�y`o��o��u�_�{�9� �^OP!�tΣ�MƝD�M�\��,�X�1}Ը���d�׌����m[�����+��E�2�j]�3��ʚ�RC��>N��7L��_L)��g��viܟ<��߱@�����P+��k��@� ���*O��S^üa��{��ء��:�\����X�r!�ET0������5(��D�)2��#�|'C�ʄ�VK&@k,�Ζ(�~v'��-��:�!t$"��ܳcz;�H��a~vF�4�l�0�&Q8���'O�0?;��K��a���^���M�Lk��C����h4��f��S��ZV]tv������r�i�������{��2�3����tJfM~�5 ���N��%9G��Q ��ێ=��v��O9���;�?<��f��/�=Qt�IB��POց�7`3�6O ��n�x�� �.+� �Z���x� p��Y|��)8�E�wv+��>�[������05�� �Y�����(�17?�u�eI�7�"�zhǖ�SN���8�҂\� PR���O-�c~q���ֱ��V��7��^:��|A컆8�~-T�{lk4^X�d��+tNhP��G��ӆEf��?:di��n���	���8������bcm	K�3(S�s�[�ƪ���(1��̡��"��
�!H$�I)��'�kC|��1��O����,�~�y���Q� ]��B**�5_������<�a���~=��|�fٌ��*D�����a��`�dg7����Ʊ������r��ڮ�d�jb, HKK1s]p�CŞ�@����3�2�����d�|n��J���ߍ]۷����8���X[�Go~����^A4��}�m`�����巸t����׋��܋����{�.�G�ygkK��^�G�^�z{z���^�j
3ck�CHOƧ�+>93�x�{^܇m�G��^�Ջ�m>o��� ���S�! D��v�&n޸��F�x�zD�����}�;��<�;o�[oA,�cǂZ:F�˗���7��������u'�?r�5�|�(n�y ~ee݄�-w0���k}=7�����5�U%��zsX��61o�\D�@�j���!j��U�Mw����� �!�O���YziI?���ԫZ�f���=Z�G�� �U"sg�TS-mIx����*F�;��ї�w�.9ޔ��y7�W[R�TɎ�0 s� L���������NM�z�{���˯Fwo?��
��&�O&� ���I;c��kD���ׯ��͛ڋu�h#Xk� 6��@��EW{���[8t`榞hȍ�����Q��r�d����4OL�h]�Q�e����!k�|��Vs��j� �l���"��������hkE[[�lV�Z���>�W���<�8TȮ��/]�(�U�֕i�ݷ���}������W�Y[��b!��6��,�F�d�v#ޒDGg|���?�v�.\B�Hp��
3G��� ������qX���f ������K�U���б:Av$Y�R���~k����^A&<@K��.��-�!��ila����%�C�ia
� !IE;K�C��2��J�G&SRc=���������Z���X}��|�����H��|��,��<��P�`TRv��E�c��"�TTy8�e��TY�,�4��XxG��8F�Бl�ߵs;�^'�f����.�p����$i�$��7�׳9���w)��.SK˫*0��{Q���Q�ԕK���}�9}�#F��Bhx�>^�N��<�n����"I~��p��M�)1� m�f��x߄q��sg��$���i��:��<^��ua~j���0;� C]�h����bx�ۆ���zTC~ɨY�K����&���Ǐ$W�Ԛ��d�m-�F�	��eu�3�2r�
J������,6�%8�<oE��C�'DϖQ�����i��"��B�s��M|W�(�.�D��p����:�pH���|ne��s��;s���W*� �;G�w Ôq1R�H ��&^��dH��Bֶ�AVY<C�uA�*�^`��m���},�N+�)�c���=�h�j`���1��`�H����Z�t]���O��C
���HXm^><�\	3��f�P�`5��\�UjC�-����W���jnGw�țo�{x+VsEd���|%��E͖���e!+�8�S�%{@�
�)%-"�6���ly�*�,�{x��$���Դ�!}`����+j�K� xJ^�t���.���l�d�Ҹ�i�/y_w��1�Ѱ����5�5��yh4��T�!��LT�>ݰ��FF����bP�҅q��4�6�ן���#`|g�,�w�����X\�:O&g03����U�
���(��h�_A<[m�ct��*�9��a.�$��bv��Usp�G�n��X4��_zQ:�K��������8�ޮv��?��G��3r4q:�+u��gr�O��n�}���~,g�Hv���oG��ΝX/�
���@�e~�.R3��g�65�����ti`;O���#��&�2L���ҋصoR��8{�0��0|�������zEP(��
�^�"���5'�-���_�淰g�Nܺq��o�8?�o����a���h}�Y�D�R�Q]�3��O]�F�w�#O����`ۮ�����W���Hv޶ksY:c��f�������s �hV�fV��r���2;J���t*r/q�<����3���4��G��e�.,�>
a�j�;U,�I��8V���\+��!���W�oԍ��]ȯ�%����!���!�∮HV����ݦ5�"@�>�O�9,ƳR+������O��-���yG��b��}H�&�/�T�([����W)O?fB��&�O�əI,,�Àz1���d�Ⱦ6(�(�����_Ǯ#X��@nc�RIod��<r �g9S�sndjf��v+�9��5����-�t��f'��?�5�_7��
���n�����Gq��'Y��3Б��)]<Ƨg0��B����/i[����}.��w��K�q�§ҿS���o�"�P��=�,#�!ρD��c�Ȗ�t��_���|U	:�=2�Ǎ�U�E��sm{��S�j���_�0�6�WYl��?{�IB؜�MFܰ��ym΢&#����]��g���?�c2��7|,b�"�� �c%����T"�E��d^�}&�����7�Ö`� ޖ}Jv�a]+������2�����I5�?x��4H`W�:o_(
��/G6�̢�P�$%�ϧ�;�]ˢ����
a��B �mdH�	wn\��=������}�<x��&��]�)�Z�۔���m ˂4���m�DD>x�H������P���Ʉ�XG��q'��sLc��h(Z�A<���F#��r��dlN���µV-�@*u�IX<����o�S� �ă�-3�	j�<�n`���r�|�;���8/Z�A�+���L&��EҺԃB%�p4d�^�Wg+_b�	fff���}b�	�YP�ه6+�iLL�avn�]�j��)�v!֒�,K0�?C����[ikv.
��p��l�u��}�7���Q�}4��wGw��v8�{~%���3��~x�>��Wu�{�����J���J�IB#�g3O�z]~��.4 S8:Bn�%=d��q��9ܹv���xL ����m1]pzp��a+�`%���KE�	|�D".ƄAE������7R(��GO���L7�rM�o��<_Ff#���e,,����4�{�p��kضw?\�(r�
�v��8Hs�k� K],�G���bA�iNa���-e:}�A4M�_�p�,��4*�Є��M �Z�p&���F�?Ma�����1��a3�~��fn��c�/�a�F�_f�caQR�b�o��,7ɵ�e��p(�
��S��͒a%L����q7I�M����[�O��OK l�fO쎏Xk���$���_:Cֳ̗�N-af.�H�*?��q�����#��b1�r%h
e����J#s��a[�m C_�ZQ �<�89����4s��%�9}�̊4�����ˇ�װ%[e�թM:���?|�1�>�D���RM���^yUQ�V�&=h���a���W1=�0��;�C�A)7$mS^��5�ZA���Éd[^x�q�#XHM	���"�q���B���S�E�n���=��Ĵ63�Z��$�p��!���;�p�֖���8r� :Z�:�y����K6�<ۭ��8~�2��vz9��Thm��p��E�A�vj3��us�=��=����P��!��ᵴ�$"nx��,`e;�9L�nZG�^�M��Hܤm��tF��3N���ָŒ��� ��Ϗ��!$ 3 ��V�:,.�$͢�\k<���v�^2�̀Em|^�*�w�#�t˵��+�%u�U�[)�[���O'ڹq<_.�M�>�A]���m0-�?��9����6�n�a3:����H9�^Y�:�EԪyl���_;���vx�v��GB�GJ}4LI���d;�YY��ü�3M>�~v3��>?vl�mÄ� �<�$L�F/7 �LJ�CI5�~�	�\�(ˡbey��aljJ �dN��+�j�НYQ��Ͽ�M��u Μ�L�W���"c4�����v������vcviM ����X�p�1�u\�ʟ����OY �F�{���'Kl��mm�m{(rj�g������<E��m��6�k�YR�0���|�Xi�kN�d�E��{�SN85�iW�?��"����u��߹em�C�Vf$q�ͣ�cM ���x���2���g6�ER�.��UwH ^�h��l7/��t�1:�tѼ&�~'��`Й0�I��<�i^��HD�~t�yt��m݂��^,�R
a�q��b�wf��8���K3b�|V<gG�l}!�_X��;bȠ4ڴ�t�;;N��3�)7 �E0��8��B�c'�_#��J�냇�>f
cS�Ơ$͢�9�y�R�w�p�|��|]u(����ZV�+�!pa��}|���X�|��Ǎd4�(C�<D!DCap#.U�
s��z.��
c:wq.�sB$"�kȝ��� �P���	<x8.k�|����Q��w��+�;�lG�Ȱ�d��?%|���=ݹ<��Ϊ �`GT�C|����x���^��w�a�����?}s���/����«ي�#;10�]�~�RM�w�Z�����ʭ��A�Zf�S���mۅ���|����4Z47�g>>���I��>1��]�hKƑ����|dC�r�F��"��Ly:iD�3Ѱ�q�RM C�����#_(kj:���Svu��idrE�od�;�J�Pضs/^}�h�ꕴ�گR�a*�j�fЄ7�Z.��Ky	5�t�s@*�ZM`�Q������>ÍRC�%�8a]/"�k�5@fm�Jh
���@�� ��6<=�M;R���#G�(�d�лɈ��I6��l٢��d+F����)�3Jf6��Z�+�fQKR��&��mݣ�i6��f e	��\r�������紆w�3��o<���u���;�$���~w^��%,�e��ސ훆�4X�4E��)W�<�M�lIf�OYD���<q�&O�S?�_�(>vZ��i���ۃG�`��=�-�a��?��w��6��l!s�����*�\��+w���&��Ql�M ��*=1��ے����Q���}L��W�ﾃ-�C�>���n��&�i���    IDAT��wܲ}]-X^O���+�q�@����dR������M�=Q~�m����(��5�Lfӏ�I���ޭ8�o��y���#���)�kڦ�{<���`��R�	]7(h8��+��G�0AlC]�lf9|a^�d�/;t����QCK�{s��i}m�)�L�N;8�ޯ/����K����ֿ{���8�(�rt�lu�f����f ��Z0=�g�I4�C9A5=��=�6�����
��<�H�n���5���
s1�~��C�����(��𾲓Tw��4Q� �ˍh2�b��]��,/ehf��\(#��U ?�Y�	��u`�*�����Og�� ��r�woŷ�~-1?&�׀^��Bwg�S��$X�Ʊ�.��/�xfv��v%D~~���v�J3 �Ŧ��ּ��D�n�n�i���#+�{�n�P���{w�(��L�����GK����^���[��Z3	�d5h�������\ٙ%v�������{�h�}7ٴ3����I��j��/�ag)i#&&�
I3�cI6����i�r@U(�Pަ�Fqν/+�fsXU����޽�|�;�9(�����7?� �'�q���e�H�+!�I�EO�l���y�U��W�����5ܙ����S��4��AJGܨ!��x�e���}��My��,5ۉ;�K7#!38�-<+x֫�R��ˎb
��8�C/���vtf;��+ �j�i�5�3�d������0(��^�ȧH0�uMS���$�<-=����`�8��C��b妭��^U��:�: ����K܋����Ƴ�rNM*I(�$v�g�ndJcI��V7��j�Ǟ=��+Jݥ���9;r��9��+ϖ�Z|��aYp޻wW|~9k%yi0���.���3���~561�����O�g�X�:{����|�ciE9r .:�y�𔕉y�y����*֝�>�X8��N��(�v2kO.;F����܅ֻ��f7�o��dȍ<�'8M��q������Qƃ�_��矡Q�"���_C��'��	�qU��p��m���`�]�8��?�^��~hdX��� �m9���`vn^��Xj"��E8֩=�Y2�1�e��)$zz�-��/l�uDY#$bZ7��0�b�7&�C��B:�u��k,���7O���� ��o����L�Z����S1q�8
y��x��n�N6{�v*ݬk. -�����?��5�͓&�M�wpץSbK�����W�}���6Ɔ�1><�d"�D� xj��I�SU���?�	4�J¡����\q��^d�U������5d�UT�^i�����n:����������?ı��Q��2�8ݲ�ۄBVN�^�+��RQ*�v^f%�E��+Я���2�͊������.��v6P���n-�
/S�o\h
y��v#u�|m�ws!y8h�E�Nw67ǛWi��zj6	%94>� �x,�:��M�6��{�@�͐�ɮӋ�a_�#��a$��qC��V'0fZ�Π�)N����Vd�e���<е��o@Ce��~i9װ���g+�ء�*�!�� x�.r'5�`�zL)����t�3��'��Z�o��#�C	ME麔�h�������6ө]��7Q̦16؍�}g��#H֡J��q!��;��.����x��J�� ��!���)nመ�B.�|*���5���`;|xR�,þ8�H��ѱ	���.���#�MV��2�l!�tq^���z9�w7q��k*Bx�XS�˴͏~�)<>j��\(��Q7�TT�`gc	�FW���N"�FQ����t���:Pw�������6��� )q?	����3<�Q7�rᜉu�q�t����-@n��^��h�i��D�K���"��g�Y�����a�!�`H�-w��3,:L ��
B��<T�r�+WPɦQIgP/�����AfAZ-Y(^3�̮5FFy�&�L����a׍r9s���Ze�$��δ���àJf@��G�m��st��G����PG\��_�.J�\>��PJ�h���L��l��	�䥸���{?�%�;y?��m�H<�����N?�Sǎ#����,�Pf��ǣC<W(�ރܻ?���@4��3U�Gc
őD�ݔV���ܫ9p��\��:
�n��w��՞��ۇw�G����ϗ�X|���G�x��)r�d����*R;�j���7092�Ź��m)Y������8�1^oz�Y�G@� ���;Xx�������ϩ�B�2{ۨ��:(��S��zn�n�&�vR���̵�n�h�m���&[�Fl��$�Z���:�|�y�ٳEzg�n��R;�g'�;�=v����Cx��?�0�ᇴ��l��w�����5Ͽ���Ն�Ci�q>)��h�C���WW��s�
E��_��8��L�S��Qb	:u��^��y�E��ES�\�tn���e�.��/�H4�ұ�B����y���G/���~J��G9HL ��i�"Q鶯\���d�k����LiM�he�N���W	��02�p���t�٢Ǉ��$*eJB�p�� 'j��~x��3�NS��4���Ho�Tt���A�����P+<k�kl��M���� ��
�Ҿ��V� ."%+��uՔL�t��WX�y�����I�떌� ^����Դ���Z��l��7�"G��8r���T�U��)�*X\x��/�l�j �HBĖ/�! O���C�18>��Ǝ%I��	w�$��\v�y�H0�C��w5Gyk�Y)�}<��\>���3��קw���[����_&�q��5t�ag;�T�(f��Un
v"�M���O�` �:���A\O`ɪ�Q���!@��"^�V�p��ט�w�rQ����n�&���/'g��Ε>��G�|���A_o�JN3@�G�B�*�Ņe9�l��(VLb���N�������TG^�]=s��A��u�7��u�
���bz�F[� x2�|�M�����|$sc��P��m�5��$Vv&����Z�͍(+J�x�rR��A3����; �zo.ZxKʪ�	_�ϴ�I���:�YXx<�wutĨ�Aww'bѨ�7h��.�l6�A�Fe7��3`�s�za��x֢� ���%��Z72�ɲ��AHQʝ]����W my m�����-?jn���F�Pʠ�Ƿ,!��ÍBI��&�����F�ϙM��e>7�������D�Q�_��W	��;p=��r��l��T{842 ���GF�Eh�b���0Z�r�����V����2�Ώ\��x��D��^k�n�j�tcb�a?=����b�0^,?���2�R����ﾇ��4ff����ҿ�e<}�K+K�D8<9&б����w�^�c�-+-�<���ǟ	̿���h4}��0;5�������XT�k���È�b�)C  6i{&�2�G����],<]��2���!�Qk��2b�-7&�&a�C-�p*u`ګ�{������[�����a;�tl�%���f���<7e�Dٽɂ���G�M�`��j.�z� V^.RnZ�Yֱ-̌�����- ��
�'Ya�(�1L�V�X���"Jl�ZL�wy�0���ג��돤��i��C��Q�
vN ����@��J��ÐL�#�P��vt&�Iqs*�p�WPΥ�5q��a���Eud�->Dng�'Fqtr�|V���,�
9T�3�����Ż�d�w����Ut���M9����J���)��#~�u�\�v{;����W����Fx|b�^'#��c�Ηp���ml��R�A�Ŕ����뵋��ų�GhTJ͌F*@\�y�%+��G^�4��}��J?�Je���*��>�V�W(����[^���j��s��h����XA��o\hx��eO��� ^��/��]�&\;��Z��8؜���M=׀Â���[,_����O0M�s՚0P"!�@ÀZl�f
o��ģ!Ԋ���NW��Tꧺ�L��\[Io��R:��O�X�!U�
Z��)����6���Ñm�ko�x�zc]���?��+�����$�x�x���A8c+��/�^�oh�Vx�^#�|]�73 �D@����v'q��1�'O1::,K���]<}���M5�W��3���t��Q�����������f���@�\A.[B�@�i���1OH��n�pT<�����af�[�t۲���gx���Ofn�"Ԍt�t9L@����5S�»�YAn_�c��y�)DYk{\5<Tt4੖��z:�@k�[��V��C�A��1q�b�����)��,>X�sOm4d�y��Q�:�H�X�ٔ�hsu�"}����/C�aP`�q�D��146�P4!�fh�h���G���D ����@!w�J�R)���/���g��e��K���/�ٽ����_��f_����sW��=���<2��mp3��'2��9�������yc��sB� ^����l)W��Ŝ��,/���_��Sb<{�����c�e���}̩������fd��]q��P+�͵Fw?�RLݟ���%�l��_$���J#��a?�א�ᓧq�����y������l�zXw#Y1 ���
�� �L7�W|�n���⫡Q+K�����x؅�d�+X_]B������=�y��k��t6���H�M�F�rn�>��NQ���� �m}�5I�*�
v%��Bw��TJ���g��א�mӤ�Q.�h��Riъ7E�Nn�N+ߴY��M$Y�H,!6��1�}������]�0*�ELF@�|I�*a���,�t���[�G+k����$���M OM� |X�x�w&���Z�, _�����~��891O�� '�	|���ً�~��LՃ�˛�5���.ՆZq|���C:��R�H��b0W_,����	�lm�?y�D��������ه8r�"�HJUlno���b����iq�����?��+��?Sm�ln��Oo0��gω%��kx��v6VQ-�PJo����[�N���'�o��! �⑭E�'vH"�!�=�x�l����O� ��@��9��b<�����������{5Y���Y���ܫ�o���K�'<(QcK�b8(��d\l��pc��$�<�#&�	�����d�(d�ꘑ}��bNl��z>�c��*r���χ��M�i�����4 ��< ��ۼ��a@:?�u��hw͚$�NM.;v��a�;�U����crݩ���V�!'{�Ŭ���p�s �XwJ`	XT�U�&�p��!�~�,|�"V�<B!��ɱ�8rX����}�{�-u�\������Q����S�J>������G�E-�W�w��[@�٫�]�kW.�h����ӧO�б�4<:�C�b�X��Ɲ�X��i.t#q���DO"* ?2�) O[IZ"3����rJ��'0���8$�pa^3Y#c��A�\���:nO�a3U�;E�0b���Sy�t �L����E���^�UΗ�V�`a���O�����׍C�	U�'"��'p�3F��z�`�����ѬɮTe�"g�
 2���,���4�h���L�5��������
���d7J ��{6���j�Dþ.�³ȔS	\	fyf�dX�w�@j ��̑�2�Xw;�Aɖ�4s�r����9/�ִ��~f{n��̊��o���ymI!�Z� 癊��i����8�I���~l0P�IR��Ԑ�f���ܷx���(�@0�vjO���^y��8��j����g�d����$��%F��?�	O0����������Hve� =�Dk��quf)UĴ�e���KD��D6 ^ϛ3�o�4��t��iR�H'������X{��R���rx;c�n�����S�������v66�ݪ�p�j���E0�nf��H��@ͅx�r�nx<�ɰWPizMvcd�zGKv����J��BFC�\��nY O;������0&�먗RL|��ܕ���
���.�� ������o>����t��?փ�g.��o�l��#a'��g�f�]@���TbL-u <� �)c�h2�]WED�l��D_2�Z1�'�q��Wx�xA]g��	I.h#�$E�)H[Ğ�N���H�$�8���Vu!�)���<�^�f��|��T&#F�]$щ��I�<w=�cbr�U�����H��4~X-^�Ed"�f��	���B�e���%� O]<�v}.z*����3�dG�Q�����kl�L�H)�O�Y�Vk�n<�d�h�ĻGpn(Lu���6�]l�`�,��C�3`�.�<�G�Z'���7�xt@�sY��9�b�̺RR�����v�#��a[���K�*=LP�5�ɕ�����g6_PZ�?���Nn@dMx}��.�"�pl��I�v-�'��|BIr��1���������si��7᫔�f��Ix/��N���G!�R���!��G�Srs>��r����V���t�;X\�D��PBƌ�1ދ"�Sb�ba�;�(�R��I����^�s;Ude8l��ťe�����`g/%7&����PX.!�F�Y������[���"�NK��م��,~���N��5�X��M.��f6�4J�-�q�$.�>��xP-_n���T�\ , �����J��
�sy4)�`��I0��]	�"��,��a;'�pv��ֆ���v��h�pO`k�W3ˣV�����H��0-E$��?@]�a��v`�h8a��|�����$�L�Y��r�b=]6��p�Q_�( � (�����j���#���� >�I	�*�� ^rk�'��L�e����s�rx�z;[*T��x�E�0J��%-CҚ�x���e�}��X6Z^��Ϸ�&�����^�i��̑I\�|�rN����>N;��pZ:aJ|����:���]��G��C�xpwfF���nC�h�r�8Y9���/��p���>;|�._� _�Z�Cu��x�dS��x��ӏ��˶lY���mc�;��ySi��3���>{�:�:�� ;�di%��KX�[x0=��vl��}rΚ���f��3|��zݥ<��FB# OP�g�h������+iZp����\�Fc�o]#����� ��:V8�`�-��:��툫�w��v|�)1�qe?"��M!gz(��5��>�݄��j��\�޻�����5�k�/�����Ԯ���t�SB�!k�~������0'�35�z�hj	΀Ё���F�!g2�˞���������`�x�� ���XI���l�g�Z�e5�5/'��S����2�i��Y�r{{R����D�=�cG��09���Sp����]f_��E>we���^�J�^Y]���LU����t�#yYw�0�7�g�exJ� o�:���w��'��|����Юd3d󭅳�ݚ���u��Z�׳a$�f�R���_b�)���ym�@b?<�V����ͯ�4��BZl7�������q��I�{ʨ�߽'S�|:% �F�ׇdW���jQ�šHD���Wɮ^='�*�-r���ξA�L�쐤u�z켤q���Ǯ۪fB�z#�J"䩡�cǽ��;��'�,�I �������l�J�Ǚ��00|[��le-dU�L����P�R^��;�� <O�
h� �H�Q�ѠW`~ce�}�k<{�X�O��{Q*�aK:��s!��P.�#ũS�q���6RC�͎6�h���ߞz���4vTa�T%wt����Ә<~B�Lޫ��J)��-t�N@ʇ�U O"v�rV���d�Qak�x.S�'VFx^���%��Q-�Ѩ%�1�RSM�IB�� '8P�-��L�[��� �.b������j��2���{!(��7�92L�6��)/�"�+���S	�ț_2��5�DC�0xXj��e�)�GK����)�G:������:ɴW�M�N����0������������.�����X���<�F�x�*�,���M-�Қ��k�aUa�9�S�*���х��Uj���=�:<O��ϫ
�b�Nl�pg�	nM-b=UF(я�7%�g�    IDAT�\��`4��'���X��B�}�ܪ&˻#�&P�g����"�����43��S���� +[�5��.T��S{Z_q��x��U|���*��M����le������ʚ��<����\����p���x��1�<<�d4(w�c@EX,�)����g���CT\a�#QYm��L褞�#]�麙�'5�fX�Yo�U� ����c���W�\0�NS-[� 9�>7\��^� Y9��� ��^���h@��̡l�2n�Q��}'kZ�dİ�Eo�4O���Z��]�6o�4�%	���S��(y��) �������`���ml;hp��O�b0��-rΜ����AWu���<YN�db�y6�b���9C�bk���Y���p��9�*9<��F%���z�5� r��]:^Y>� 0@Ͽ���7��T^�G�`}7����FE}gW��t%��[ �`���-%���P�.7��Ǐ*���6�|�`�v��\�$+b���;�9�dga����H7~��[�KF0��6P+�4��N�ѣ�ni,F8��}x��2f�f
G1v�0"��{��/o��n�"Jc��P)cx�y�3�
�'�$D#�`a� x�1Ҿ�F���*�k��KkH�^˰;<0O��5�)y�x	�x(	�tUNm��֨�C�\)p�XS�Y-��A:{��6�&�g��d?|�-�q��t{�z5$������yu�w6�i6k��lq�3�L=,>m�A�B�C�d�e�c%r
}"��!Z��?��g�$>`)׊��Ic���v2B��_Wƃ�`PVM����;��&q��i��V����}�=841���y���i�ҫ�\�]�_;U*fƅ��r�j]EP�X��7K���SM�@��}�stt
I���%4{��@���d��5lJ����v�k�فf����7�AaGh:0<�����������lh:�?�vOIլD"ђ{ei�����ʙ=u��'�g��8v��ʏb�����x8=�j��:��ca��qDQĻ�H$�G9�Ď�O�7_(O0���o�h\��~6�\�*�?�P81�4������e�7�C�=���f����?�uD���c������'_���V�t���Թ�>��݂ |�Ǌ�lf��8����l �	��A�^��Jwp S�.�5Ỳ}�b;y�g��da[��b�	��0"A���b��X'VҴ:u�0N�<* %͔�n��"��bjz��O����r�)��Ξ~�����S��0�BU�&����QJ�u��Q�J[2m�dھd�%��������tp˝�`���䛛�N��<���J���������?%/N��M�c˻T6��f3I�Աr�9�`��� �� ;���yQe4~&Mk-�S��#[5s�4�@���\�Q�~tu&�N7
��%��dq�[�?������caaA�?�ǰe�����=����&+HW��4�B-#9`˿Rht&�Prޏ:}�Q_���K�c-�*�WpX!���6:خ�>�T��O�� ����U�uE����c�@5�DN>Le4�N���w����9��nD�Qv�����0��w�v��eTT�*��h�����W^����A�C~,/?Ó'Kj��=z���� KG� Ý��V~M�~ԗ�$����￧��uƏt&/����۸soJ��|�0��$�����ڗ��p������R^�	�(9����f
��x�R3 o(��ק5Wq�d�Z���9b�Q:�0�ղ��&�J�s�)�h������z�Znbx�Zx�sd�,�L LM<��ҙFl%��k���F�[3.�3F7��D�$�{���lR]�"���&�����h�$�g7��i�#�ޅ���̡�39�S�k§�Z}u[��`M�4tgk����up�xh����d�~�!���F�E�����%�3�Yl�ഇ��A%�����'���3:��מ��ٕ��k�.
��i1�bLɔ�|����g�~%	����lo��ݻ�#(�3RGB����ʲ��F�|J���004(�;��	�Ñ��?v�����Սu4id��73�J ����@޽��xx��sgOb���bI��"�SFF�@���ǘ��G4��脆s=x0��/n��~�.���	KJY/�k�\~��[g�V�d�V��h(�����ƫr�2U��WmV0�H�Z�x7ɨjY����tΧ�y��F H Oձ�x�/$	��V`0�~FR;�@�~��u����|.�]u�c��wpbh!�K][��ߤ�i������qdX� 6�iNҁS�����5��E9�R�R;�mƍJ���P#o�.��G�ѻ�����>nz�Fd�x �3��v��1q�L�G��AN9�A�TFOGⱐTtLaQ�}i{s{��Xw���}�,��,�ٽ�� %�w�FRB��[��r$S��hk�� ������I����nI�#�$f(I6��F
+bD��v@�w��J��a�N?�\��x��N���v �fj�=v,H2TP/����#�k`{s����,R{itĺ�޻�Ǖ��#v�3Y���p����r1���PWb`dC�#f��Nx�>������]z�Y'��*H�*
]�+4$����샆��7j�+b�Ǉ;��Qͧ஖�>W�����h�Cg��N����o.|t��/���+.ǎ��{�Z@2�z� %ƈ�v �q��Յ«��Xa%H o�Hұ�vq#P��.}/F��M$��8��jbgm�3X|8����c\�O1�W]����\�G�������|�Y�W*���Rnbm�����d}�#�C��[z�#��7��kJ�}��!?����p��Β#���^�d��5��ʧQ�X<Ed��@%�rv�kK�8U[H����0��01cE��F�#�����4�j��N�k�U�qiM��hӴ5�ͩw�oEۍG��t�K#6<0 0M;J��ɠ�5��w�o5,g�X�_�#O�-i�� �N%|]�b�X����q˼
�����O��q��'��m$���}�3T�؈9j�?��4�[4� ���4�<����d�V��fZ��waz�w0r���u/�%����7^��㇌���`�-�u/nݟ���*2R���0������F�R$J]�}f��T�x���uS��:�D��KDB���$oK���H�ۻ)]Ӻw��wk����!O�Ɔ����o'<n��5�O��΃�V4xGg��Ǒ�E���Dz{=qĂnLtc�7	���T)΂����b	�{E�|�{��
I���I��sv���"r?��}�`�(j;'%'��8s67gX����V��dQ:C���K�a+A1	�\w�c���K3r^����޴�[ò|��H˳ʤM6
%���b�Y)�O''�Q�� �G;��_���tfGC�u) �������P��&��K���c��t&�uo}p��v���$��2g��k�:h!���&Ih80iN�mJ��"���HHظ+%x��o������PH�`lhgΜ�N	�k��Y�(ݸ~;�����&vovNJfvV�� o��6�ͷ��=���	v���K���D�*X��ul��n�so��ղ$�d���b��m�r�t��,zI4esi2�XT@�$���cL��"�����8�=���ƭ{���[�L �g0�/����-T�9�� �)va��  �3LѮ�2�K<#�h�E�<��~�x�7���.��mTNH����$.�G��8NqgfLLo�]���{)�}==�Jv
������*‏��*:;����pr|D�F׼$s<fx����=
",�Q��%?�Uj��ݬm�{Y@1ˁ��L{gj�Y�T�Ƶ�[�����X<���ՙ�!�g�|k_���3p�\Fu�-2v����LD��)�5�N��R�G���������ͳb����X��B<с]��mXf�#�#C8b��yψ'������h��X'�$�������"�얜�!B�E�9{����Cx�I�.]�nI/�ಚy�������b��7;�~�C�I'mֲz!�fI ^r��0B7��}<_Zē���68v�8.\��gtgs�Ϟ���X~�$��9�T���p@��f�8;���.$��uVe
E��]L��<3�%0�)�H�� ����w��C��[�Z5�w���+���T ���7����_�$�Б�/���ہzŃr�&�"�V�M�e�`�$l%U�4U���j&��~��E. \�&Ȉm�*�᠒!���Lmma��#l��"���b)'��l�`��J���K2�<�5/D��/1\��D�+��~gW���;�{٢ ��n՚�ըm;9�$8�v �M�q��M��B���N�e�bN�K�U9�}oVs��n`k�	�>�4
k���5mA>�)�E��֦�h�i������������~p㒻��93+�h��!�0\\�T����ܘ )��V�&M�}���f���~���)q �-�bک':��5BgYX��\�0�����V�<������w�I��*�[��v��a  O�h�|.������|�lS�������5l|��M��H��^������ۨ ����L��)�����x�|Ś/�3;�7�yW��Ç�X[[���RʩX�g��VB�-�ZÃ�HtDQ.fܟ>}�k;<:.� �- ���ƶ��L(�F�c�m^�R������8��c�{J�K�)��#9���6�vӚ�����7�R �£Y���$"~����\�@W�!�����p��6���,<~���ϰ��7s>?.��N]������]|�6����:� �je1kAe;����G���ϵ �\%��i8��)Ν^��Y��*��r�;�������VR냌�u�	�=��(eҨ3�0���/��0��dd醳���LvWI��YB�6�����9;l|���i=��,�є�m��K�
�e���faַN���病$A.�39�xtl�brV���b���m��-N�3{82>�?���0ԛ���s9�L����r3����cjf�|�V��<]Y���9�}!3,G#�Λ��e�,sKn�km
!�Wӱ`AC�Ы���,$(���@���W<�3���C���~�����?QZ��}�@�������"v�B���g���s15=��~�LFW_?�F�խ����#[!v�i]���H�l�)$��i�戏d�۸�x�b��.�=�8c�e5��l/`��$4�IJ%E�����!�s^G�zntG�V��o�VWF��\:���=%θ%��e�Ir/�w49�A���޸��Ã�k�a�z�"�h�l�&����H?v��\ߒ���Ԍ�<�&`R9��E$�����9�0��ј�d; n;S�$(ԭW����.+�� ���1׆���;~r��We�����
�Wu��8w�.ww7��e�&y�)e�O���Ŋ����N"��R���̜_y�C���=�Vi�{W(f�Š�_j���x�t	�2��8��D(څh�[�]�mj �P� >!�7;�̈`���sϝ"Nא��,��FZ˙*ǅG��Tf��{���[b�	����m�yn�I����������x�[�R�Z�󶳹#I6m[��L��hvw��%Ǭz�3�i�)c���Հ/g�Ѱ��^�$V�V�[&,�e>��C22�� ���(���M�/o�*{��L��(�Yɲ˟	���}]�87���i�J��W��:�������\���Ht��o>o�<m =�#(��Ӏ��֏"C�×�Iu�v��[ӱ>�եTC,�dfP� �!==	��R0�)Dme������V������m1��4��9���6��x�\H�!-�����(��8��]��"j��x5�kL���4������ڱ�k��Fi�p>�� s���綇���p�`���L�~.�H+�3��UϡQHk�+�5���1���ǔվl*��щ�n�����%�E�;�ي�.��9��B�M�֩�q��{0���)���z��HO���!*�#��˂.�e�H)j�Ѻ���5�����+ ���~J��C#xh5<L�J:�bÙ��̩��j��9���4 ��>�mĜ3���w�i#I �<D�vMR���a|��wP���/��G�x�L:e�R~���s�tC��\�C�t`m3��~q��9�d�X��`��	����@�P�'�|�Ǐ$[
<�,�&�f3��\C.�U��A�r)gS��~
1��=#*���|��&Lѡ���*ż���*�rr+ �xo�M�l�f
��Ϩ+B�JH��M�O>B����W/�{！������{K�N�P��{s���A�dh��ƻ��{?�nܛŭ�d�H�v-���'�����; +���;��W�~�����_�h���Z�Zo�Kw�����̾�mv�^L��L� M��a4��.P�gP�e�!P�%/Ox��G���#!��nHB�W��s��se8t�pI�o|�9h�T�[��ܓ=��7ù,���9l41�<b.���@�����Ĕ-�;I�ZSK� �5���8GPHc����O~��G0;u��.N=�cǏ�`pp��߉705�O>�_$���/`����qC���H\�W��6�]:f��m�)Zd��� ��&���@���j��V�PPJ����ʮ��^E>���dDANt¸��o�ur�ȤR�)��5��q��X�`��"�/J.526���I�O�\��t���/�`,��z1��Ύ�X	��t�`<�JJ91�3��GH6���4P!��n�ضo:g�s��g�}k��^��0�=�!O �x��� ��ړ)��F�\Q��`>��g����9���Pq��\DwgWΟ�ѱ!u=�#`�e�aF�}t�f:�0�,U�zvz��ǣ��"�X7��5g�.�fa7��� �U�oHm-�+"O��Y��f��}9��g:�����mXb����O��`ɺ�!�Fo���
��❫�d����,>^PI��z��e�!��Խ���G�#���ϕ����.g�K���O�Q�;[�t��?q����q��<^XD�T��ɱ��[]݃��{�DP��i�S��K+��VM��t�LC%]æ��@��.B�[3$�9���0I��FvK�y.=�F[^�|�G˟�&��|�� �F�my�F5f:;Ĉ��R�� P2�k2a�4��!��뼶!�E��ґǯ%�J��fH�Jx)���!rC�ά��"P4��H�,���ut0��m�kEx*�����_�{���ٱ��?	�v������]-7�>���@#�r�È��(<�a6de�&p�P� �0��i <�5��M��x�i)`e��irOǉ:E.Ƞ�S�x	h�Û���,� ��� 2ΞKC~�����Od�ǈ����9yMƜ,5+p�&y��)�1�p�L;q�q����ik��6�	l�#�d�V)u1,7� ��4�k���Q3H�j�|
���h�X������PC�OU*	�&�xLP
#�'Nf������)\�Z.%��}D];�� ��bqZ@{DI�dBml(}�i�\Ƴ���Ύ��F��;-P+�1&P�!_�#S,#]� Wa� �X&tZVO�M&�䥏ox�|�}�;C��O�uEΌF;��UK- OpO ��￧��_����$�=:����i�MV�$8���D�T��GOװ�]���,o����x��j#��G�����6�,�=u��=�y��j�p�X~�90Z����y�r��d�w2���hr���s8|r�l�f�����J"`rb1jY���A5]b$S�6w������M�\.^�����G3���W��2�r�޼zQ	���dk]`I�.��0X��/� �Xys�O ������������؁�J���ݬ���4[�bkc� �&�������l��M7ά��������p��c�Q�)�>������x8Ӫ��E)��&;u Q_��� T8#���C��|�� &�z�ӫ�2    IDATՍX(���ϫ��Ȭ�fS�v�A>�ViQ3�VVV�M�m�����V�'&&0:4�b�����Zg���dßG�(2�KKKX��4{�����9� _C��E�K+��uu���Oq��f�V&��#Gp����
v�,z�G7����i|ysJ�a�����{����[r�a�JV�� 7�o�?�1���{#1�,�]��b̓`t<�6Ző�7��ة��a�i��[!�+ �����#c���_�~��a�(�����9��B���<\|,~��Q��!���'��_ܼ�4�!z-d��h�JHo�* �F��,E͙$��V� ߇_r��TH"�	�E��l�ֻ�]ϟ�.+?����E�ТZ��1��u�.2���Lg��C��g��F/O�P�2Vh\1>8����2d�6ܨ�@G�b_�Mh���2�4V�-�������5Ð<JY���h V���]&��l���m݉9��t��0\�J]�+̀�>�ʑ�[^;�O�x����|
�t�d�>[*iN�+W�.�L�����W`�9���2�$�aL�##������<�6�����8+V*i�Q�?Ы�qf�<�wOQ,PF�iK�{G������B��'�����$�&=��:t9�3`���� ��5.���������r�}��I��L��v o� ��΍�1�3?�~�m������y
^�P�o�eȯ��<��|Zg�#�������9!�|ċķ���b��G����slTx7υ)�h���=fFL$��@W��sF�>��ZЍ���?��/����ι���������/|���d�S�����8u�"�4C�d��,�
���.X�'sh�� �}�7�І'	m��h� ��$!Oy��[��I�&r���
���*[��ԷW�hоO���y��0 ��Wm1��zv�HMl����p7p=P֫�JF���
+r*Ŧ��u��tE���W���>�- ��V6���1:���ɭ�h�R������Q+����~�f��L���I@@��$~_M@T��c�P��`������Z�V�0\�O8Lc�}[�׺�v�-/J��d1����j�)6�mp	��j���{9���[�<�7�RX|����}�h�����Ӵyk���@�Wsͽr|}ۤ���TS� xn1��J��x+E0(��������Q.�_����������~�C���UD�~�j��Ф����^O_lbu+����LA��k׮���������u������݅幇p7����Q$�8��H���XzJon�afn^_�PF_���o'�M _����������;���^]W�G�	x/���~�[��[x���]�;	��}X~�����Q���Cc8{�8��@�Vс��[,���l&�!����h1j��|�{x���o>�F��k�_������dM����ں=������{����dVXo�W6B̷��샇Ⱥ��x�ɻ�=�(!�I���������QϧQ$�g*��#��s�p��̱8���u�|� �xbo_��c�������˥�i��k<��bkK������f�j>lmm���Xx4�R��b�u�\M����۸|�Z�b�i�Gw*��m����>��~�`yy=�7�|�<C�DZ ���:u��8�]��� ~�g?���a�M����:�F_�$3� ���u�.g%:�E$-��_}���E�Ch�G�"�#kj�sl���0zVs��uG��i 0]%�Ѩ�I�
x~��ٜ�G�&)��0�ş�m�:<��>�%\�"._����lm�#���5���R�|����[X���;���19�|�������X�z��5�S�e�ٳ��<_�>_�^+/��aW�$P���z{W��@u�Ak�w��۝�Z֧��h/�M���@���a����M��&A��V��F��L�	�I;��*���X��$r3`���$Jv������c.A)�'�G��l��"%����F�NQ���*d�rǢm�Ҋc,�c�|͒Hh��;sr�q�K���+�8�M�1�{M �U�`��o]�&������_x��%g/�ݽn|s���8q�$��"��c}}��W�QOŁ��d���L`|t}]��z�8�奧(ʚ�id" ��,|�@���#	즳2& ƃ�t{��g��2K9�q�"&.;iu��g����s0�����Z.5T}P:K4��������>�&�7�E>W� ����sm~��	��)�c��Ay�h����\"9lHG��[S1/Y8�E="vP��tk�s�Y�PP�l/ |�͎���q�]e4
Y4J��p���u������� ࿹����˝l�j��@���;�x�.��:[�u��P�du��7�"��C(��bJb%�d�Baf�RIy-�eK'yz�A���ެS�Q3�M�NukXLi�f)i��c%fs;(�.������H:jk���d�6#�j��&�p���� |KBc|�]����������p��RHo�P:*y�8(��5Q��V�e�!BF���[ O� =�����u�L4�$26���N��G�n^�{��w���'i���A�׭*K7�PC�s�,d. �`��}�:�#��a7�ý�G�_ZF�ސ̉�1�;��+�u��? ��̷�LKTV��?���ʫ �S&���Hh����>��"~��_a��m����v�5\}킆��������5�D�͝,6�3X|��t��dO?�x�Mݟ�?��3S��}���p���I�X\���:zz�qhr�8�aAYX��.���U��ҳI�z��p��?s�j7���z���ai+��:ժ�=��S�U`Њ׃�~��Ocs/��_���V�^��=��06ԏC�c�krؖV~��:N�?{����=�g����;|���y��M���,R����Po�Z�R�[���J[4l����Ѹ�� ���Դ�}G[W���x�/���ܯ�B;�oz^y��������2�{���)D���P�W�t��7�/�����pȏ�]��Ҁ���5Hf[�[��3]�w����R��S��Ŗ�%Ņ�N(t���z_�pG&�Y)����Ӎ���P��~?zz�0<:"���(���_�G�Zf�U�,��Ɠ\�e_��o�v�{�X]~�F�"�@G�³�������:{����?���+�����@>�)+�)�7ǹM�m�s��'-pj���rs^!��x3���8
=�(�oRV����?��M�=q7���b�N��cT>���+-'	6��"��ޛƓ�g�|��d?��+�|0�|͍���'`�����+���zK�}�5u�*��W�	5{;��O�b��%1fӈ0g$�>?���0?����i�7�\K�u�̝��dcC��gp�D���or�^�~�9��v|�$6��&�2J��j�y&Lp��-�}�L��pX��r0�yiAeKӮ�J��&�f?�o�'a���a�b�`�0�N)����ޤ���o�\+���R�?[�~jO��h,�c'Oj�wq�	�M=��؄�/�-��+;�[�sy==\�U��OL�k0�ϟ=�����vPg�k���T'�"��ĉ��@�o�J�
%$���� +���k�����0}]�6����'j�m�¬?�R���<�x�~+fVi�zr^�̵��0��ie��*��oSgf2�@��<���y�&@1W�ʂ�N~�f�;I���L#�4����@��l2瑑둎$��s��{G�_Gҏ��(��2*�t�S�ܛ�Oo���r��T[�|�ٿ)����q;]�Vn,Qߏ�1t'{G%��0�wY^����Yf�&u�n?
�B�J�u��7l��X˝�+��JUde������ r8�7�Y�o�8(h�p���Z�m-t�,�kzz�e�<`b&�btl��x������; ��N n,�s�B���E�<u��װ0wG!9�Pv5J����Mf�&M�s���L�N�N��%K����S4�6J�Z�$r�����R�9�4F���)�g��R�!���l����r�����g����˅��Uf9P���~����I\}�M�ݙ�����(֚
��&�yO��Eg�:��� �h�Ų��lK�; <ݑ$�ɥ���3a�C� ��,�:�;>2��G�
����F��B8މL���f�������[�z��������$�8w�z	,/<��r�!�f[��1��k �O*���݋�<_^W��#э�����	�\��k�R��cd�]q3$����='��C���\7�����>�]�(M��g�0u�����'162 k;e1x�p�bb�x�����IeM�?�~�c\���Bkn�� U����7��E���qFA�e�}�Og�V���[��wM�Z�^����8{��5GB�:��d݌���);d���'Ў����Pz�����ʙ���j,i��˚4\�S�������{o�����K��'cgk[l��>M���7��飥\E���H����{���?�����O�'���Yy���Q�là�bݑܙ�����8�~�}�����裏��I�t�՘{&�iC^Ba�ؾ�D?��{x��5볳��b)�V6;N����V�,DTL������������'Ϟ��]S괉�$m��%j�5�d8O�s�8�k��
[ �J9��(	��n�J6%��+p��i<��+K�G����E��Npʿ���8�^�"��cdt��C�.�������#x65X�A�X��-�>�BC��6�u���^��/�-�t����@�f%��s��v=h?����_k�,=�4�$k�ov�k۲s5�L(6�j7�KY��C���fG�aOF�KU�)�d�l $/�wC���F)���e���Y&��g8]h�����D��P��⽡���7��g+�>�U��G[��K@�-�8ՙ3��n�MF���,x��d��Cs��^ȡ�3��}Ong$�JecY--�׃'KO�x�	�67026�K���T�`zjO�?7���|��;�M�sɽ����OD,��L9&	[�Fh�����dz�c��q��ʄ��"Mb/�G�\��#UԍG�1IK(�N�g	;�
ʢs� �kN�A�{iH^)�Ъd�$6�EHm��^�rXr\��Aj�UTձvܻ����e���s��g�Ŕ�a��T����t�Lf�Cj xa#u)�"�7�K
�hJ�Vї�b�'o�Xm����>��92�����m�?g���/����\�����q+U��P�\�ZF��=Hvt#K�eb�j���k@�I u��
�Tl?q8�<�����p�������
v��*��;=�L6�7��f�䭵X�Y�B7�X�WQ���$�:��Յ���j;�M��q���. �Ц6<�M����NW5�lk��YH��F	?�7��4�����^��$u��n���x�&�F��\,��x7��ìL���v�a��/xh�XǀPᰱe�`�lД�P��2@U*0z>�:(��O�ڴ�n���)��3=ѩ�WxP����I���;r����<�A�.j�tm��(C��S����/���$4<[{\56����z9 ��?� �r}�+,��0�D��1�:~G''���H��)Y��O����+�}px�.^�A ��ζ{�`gΜQ
��y�<{��d��̐,OS�0�
;�Hes�_x���yI�]ݲ�:u�8�һ�2�J�0<دA1J��ђ��۝d�c?=����8w�$Y`�LM+*���.kpuS��%��N'$����'/�/��ݴ�A�����8���9=�o���3��ũ�9�I��i��1��K�ȿ�;�?ޝ=��k���i
�X��b��׹��k劒�����ꀷ�0&�V�awm��(d���˙����ѲS��/=ո�����⹳�{�������Z	"aSV�z�t'�A(܃�w�<hП��gx�ͷ���#|��Wz~�~J?m�"�i����}�V{�+����t���?�)�;!Kď?�Dm{&_*4�L+�:�R��1M�������/�լI�ΔL��l [țA��	���}�'o8�t� �>_��������rZ!��z�0/�Fg��	��s��P�<��x5�J�7��P����e�LZ��Ai��ww] ~�;���&N���R[k�f�����w������'s����ɣ�%�dG��J��7n�ޣ���\��:zM�S���Lb�.4d�5Fi���7b�@d�G)���ɡ��v��|8]�?�y��l]�, )�xxgP�<���u�-	�����;-ޞ��US���deM$4<l�f&�Ǥ�5�J+fBy9���3u��S�x��Q�g��Z����M�^.pf���PggX�6i� _� ߒ���|
�yyXP�A��X�$����E�hV�h���／�XH����{�u���f���w����L1��'O����b��ߟ�����h�@`Z��3ej=�]��do}m�TJ�L!U8�N$�3�,g�)���?v�c�F�w�al�8�US�8�^��PX�A}.��[�AWt�1�^��l$$�HUZqu?�ݖ�3�f;�;�g�)�d%mH��$6(�a��1R!��g�	����rv�X��]�jE|�f]� 8�IS�L�v�P�M
 5:d�:�K��rj�	/��BuO5�ȇ�罱������v���l���?���o����{��պ; �B��~Q��f˺��u�o��-�+�Yg���24��ț�A�!�?��̍v� ż4���LB�9�t!��F&�f4�d��7�8��-�U��Űi�����8���6M�eZ��-2M���S�n&��³��<���re: ^N�z�;����P����i8ѧdR�7ľ��E<�O���M_���L1$H�`�M�%;bSۇ��ץ?-{bp�	�p>�-po.�3׻�[[E�B|r��N"�H 	���fk[ix�"�R����㓭�4:�z����n��E��O���@�_ߺ#�$V���"ny�:��� ��I=}b�mW��&8���k �i�d��c���SO �������ڪ���{}��!��G�XӚ���[{x03����sE� ��������կ~%p����^�x��8��װ����.L��
���D�+���C�#�T:��>���0���g �_���g�#�M���_JS��$z;�E��V;u��t�����Y��>���V�6d%���7p��	��;�o�ȑC��>T����*Tm��U��q�ރ������B �K��3��pI���i�8��d]�e�ej/a� u��1��Oa�u�۝6ڒ9u��I�w���v���	��b��ߪ�?���Fq��	�G�C��Q c�ז�c���΢#�������3�Kt�g��[Y]F)�EOG�==X|4�_��?	����s���/{V>d��h1�!0{*���n��ǎ�ٟ��@�K/i�{�cZ�5���.�+Ȥ����pOg7~���V�uO�>�?��?amu��K�@^ZJF@y��dC�]	����8��>j�*@��8`g�Q%}�Z�.�~ R�,�,��_~���9���k�|�DBǜ��_e� ��*JQ6]H�qJ,�`h��Q6";A:��Mnb�	.}�*w��(4қ�����m�(�8���ʋg&޾� ?��()�';����7��������,n�y�{󏑦�4YK=�}������4C�,�H���
��<�Xtӓ���B�	�A��ӎב(�i���h�ۂ�Z�V˄Z . /Dk#C�5�tj���;	�2YPW�������Y{�縯,K�Hx�	G�'E�.UwuuUO�L��)�e>M�|؞�����ѻ1��*��D�hA�$H�$@x��;���2���f#f��H�������;��sϡ6��G=�+�\X?t�R�3 {��F���q�$��	�� �g��+��}���P��e}.��<�'<4�9���s�,:����˪���ۃ�C���L�"��'�^�	���G�H}.�NG����|vvFZ�Z������K)�7    IDAT�=��/^I���9��������<��gc,�����م[�_ I����DW �18�X�t��b�Tt�>��k��V�?R#�6I��N�./S����gy���0�d���R4.��d�{�	�as��^��� o��3�����&E	\��m���YG(
 >����*�Y�i�,j�1�<pW�x	�*%j���8�1O˘aaJToR6�;jf:0ˑTa(d��atf%��H}�KZj�w��쯪��s���G{[�Ϣ����R,s0�� ��:��(+&!@.m�ƣ����%Uapx$����J�` ~��dx`�X(
��-;F�:&��*�1����=42hi�e]I���������`�1?G��mZ7��Pѕųs#d!@��k����������T���p/�S��3I���%_> 9@ƿ)A��a$b�)�*��E�sU����Ȉ�Sgm��/��4SQ�=u`�[M}���E�gQ�o������v��EK�;���3 ����}GgCd؈1���(���&(�4b�� ��t��R0�ش���F6��D�����/^��F�d����X�A�];�h[X�!�0�č������({2�������Pb�Jh�ϊ+ �b>+>�H��ɇ��M �������>�S� �ӕ�E������-,-�>�T�<!+����ӿ�{ʋ~��_�ӧO���2��ر��\/s��t&��� �m-R@
,�����q1ѱ"\)K���?�_��o$�s��?yB���B�µ˗h�e�FZ?z=:,�l&y���������r�� eQ--|/[�n�۷o˅o���[7˿��O�����˦����2"����%�t�������.�k��|����M�wˍ�d��(y����"vpl�% o��r6��o��ۜe����[A��X�[/3�x�}]9���9��>SJK�\�)�ʧvn�&�?(�bd���F|Ajw�>�[�n�u���h�������!���G��y:�X?��(��dzz��zг�!->؞@Ő6����u�V��g4p��ؚ[\�4��8�j����5:�dT����P2�fH,���~*]2��|���2�z�`� k�o@��r��D+�WE�zFpu`� ���Y�XO����HH:����Y��J��Q�� a`���>���hZ�c����`΁]�:���'X!������;-�X��A,y)$���X#�:*'����Ҍ$ףd��,0����5�&�"!�E*��Z\]����ܺ?,wF��2����{|�� �G��~,���3�٬M],0�^?�����):'e�f�����ٱ�V�o��4Ď��F*B�����u��7�PeQ���������:��~���Of��Ai��P������X�2ȴ4T��IK� �+����{��d��MD7υ��
�EB�u��(5"�w��󭁁��Z��c2�&��<�eSS��0kN�n�t�RB1�$8?,f��^%pʩe�p��L� }�]rp�I�V������4�g�����!$?|(ހ_���/M��L������3�RWW/۷oc��sqn�8ٜ̼~��̥�9����<�.AZ����및L�RQU�l�f2�O�n8+�c��0f1|Id4X]^���;�p�`n@��s^��\F�^��ԵUr�+)+�t��6S�?|��s�i.�5H�m�}��c�WrY��:Ea�uǽ�j�|�n���&'�|��/G�A��jd����Wy����kKC䷎���� ��~� u׹�7�y)�> � tx�:��Va�E�֤��I�[d����ݳ�����W�LɃ&
J�+�%N@f*kkAE<$:�+.���/e�,l,8�B��>o2�v�{�)@h�qC	�gY�0H�6-g���>�� �j��8Ա0�D8G^rɤ$bk����I!��B)�6�NIE$$^�5��d�k�c�+��l��������89g'#��2�C\�`WJ ����`�64�ł�hA��m��MZ�NI3�]�Rqb%9�@K��'�M�&�����ꔃKUm-�$�ZF�M�T:|�}�#x��Q�qgH����IN�|GB�U�����h�Ý�f�ƍ���+;��l
&��T�i��2(
�1`���
�Tdg5��v/��9T&7 lj��Eq&��Tq@ �vw����G�����$��'���r��!n����]ZIm񸄪"L�[�_�?}��=����o@>��_������=^y�wiG�|tD�X<w��J,�N�l�!ڹ���h���/�?�d:G�u��aټm���)�����V���M���);�m�P���;�Ri~0"�����ĤLM��}B���~,6l����_��;y����ג=BW�])<'��r:e~~���k��dC�����˻�$�[���;�r��S�f
��CQ�����uNKZ�]S�*���>[�xfj˟��\� ƍ���on��M�omϾo;}���ȧ�
6�T���9�o��S1�A�+����;�N����{��� Sr��2�H���]RHh{�����O���{�HwG�,-�s�`L��q�{<���}��[�p$�`�H@$�d�P��uJMM��LN�k�i�f��^�,����(�ꦖ��O~&�==Z��"+�ड़H�M`*�����Y��L$D��L�6�I0���U��4`|�J��{��d٭y�P(弯�B-��P�� ��#��{0��$V�?pD��-��+`fEt����\9q����:@b&������B.+�XGJF���5k���Y�Id)�.c��d��KYZ_��ۣ�C|�tR���%�X?�9&O!�Cѭry�|���.����SJJm����nK����eWK�ۡnGY2{.������G����e�V"��f�!�;3܊�ʙ�LF%_��@ч|4̏��:��L^�:ڨs�1奸.@9-	:+����a\1tE<�R`N������0�3kD�j��ZvF�N׹v���)A�x�_��������Aa����`�b-$ ������Z��씵�E���@� z}c�l�Hk�'ϞRz�ճAmN���������RGGk���`~
 ~qfN>�'s�ӒMk�;�R쫐0����$�G�b��7�tn��C����^����6�g��D��l����Tkˠ&�gJ�z�1������-���t�	�c[�!]�J�n@z�3�Uf���ɩ��֟C��IHgXHbG��B��1�Y`��gXS�W0-P��=��σ����/�@٘TsMu���W�����͔�2�y��/���h��I,�	څ�>Cu]g�$؝��6������i��ajXh�Q��~^(l� �y����5�'c言
�Z4`ZX���]����_cmW+h�dTT�z��BXt�)j!�y�����#Z���R1P���ς=�����W���1'�X���wH3Sf	�(�^KveE���__�xb�!<yl��%6^77j��2ú���yC% ��i�ce@���}S�[��ڥ�Z>0`���m����b1g<~y�w�� (H�>z\jkk	j���=ہ�*H�oɅK�()���3�J��F��tM`�zD7F�ܜ�p:�§ab���I��˴rz8�F&]{�3 <��9�xO�3�:�|O��m��|lyQ����Y�
��������d�?��_����F	M9DtP�76�QH� �G�<���U Ѓ���G?��d�9��_�F����3�_N�>C�ǡ[�e��mnZ���|�1~�.�\XI �5N�C����9p��ڻ�]�_��2�h�z�cǎʻ�֖�0$6�?��3�u��
�@�HS[;�����/�}!���T_���mfS`���/0)���	����a>o@"��r��3һi��z(�<�x�)i��q6�-~s��ŀ1���nQ�n���]�=�0��	��ɢ[ o�bgдl�+��.��sI)�N؅����&�*藽;����{du����&���>!���?�2���yih��/_��[�ezfR*��d˶m6�	G���u[�?e��w�N�a�ź����AvC�kkQ�o�c������D�L�*�-���߳O�o�)��'�{�z��o��o._��羐�(�݆�N��G+��2��|~��[��u��ȤI���$[�[�n���n�N)}p�\�nM:H�}���Y�]B3dk$V�ly��lĴ���<�; ,p�@H<�-1T�w
 OY�S�� c�F`V��(�!�4��2������AA/�I=,�բ2��,6�?���\������|��xu�/���i<�ǩ �� ^�w=�kSi���Ot�ݪS�uU���?�0PL	~[�(R&W2�|�t�w�c(�}���H��R��4\/�}�پJq���9h�����j]�젶���3.i�rY���\�  �p�,y����qX�)���Fވ�$��Z�l RY.��BX�����C�J����i���r�(�6Y�,��A� �"��"�KK]U�.��K�������]XZ��.��?��4o����A�=p�Y��b!�3ݧLF��deyQ�kx�����y�E�x�YG�*��^���Q4���/�ƃ�tvvK[{'Ib9��a&�����qf�<eCW ����K�lZ���1�[H��&,6��-����X��ax#�n��Y@�&��6P�C�o�&��gx�7��b-p�����AIg4I[]��H		�>z=9�N7TWH]8 �\b9��_lm������-�#���࿺|�+I��T�Ex�ӊ�XfA;����-[����p�,���-��
WJeu5�F]����"o"�d'�kj�ޖVWdaqI�1T�`�n�װsq������+�������d8,��X;���@��VC�n��x�k��~���:-��6R�c���B癕����RQ�0�����TW)'XZ����O���g���5�[�es)q�p��{#�#-U�$���0:Mn(�zK-ذ�b��*7�o�d�I)���b �v`�%�c�2��N�kl�rЦ۸q3ے���ß556�҅� $��ݸ#�/|+s+���!��9C �ͥ�r��#I�0���hT���di�j"u��P�2}փ²�EM�Ip-2�6�Î$�E<�^�T�.-�/�+��4ĥ��C~��3�ɧ������\�X' pA0k�����1x�re)��r��W��-�|��ӧOKOw�<}$���(��_�B1��HZL�5E�����~�z���x��������A��-Ϟ=����twuH�4����k��� `��	Cwm]�����ljzR�^�*�^�`a�ͦ��w�Q���5��7?�+�;@����<z\�:	�>)�K8���z��wg ���E�[�YK����pv�D������eݚ���:%X;��Ǫ����4�d� �W�<�g�f9yp���������ttT���a�裏����zt���j�8;?#��t�A:�Q#����,���w���39|� |��p J���㲺�Ʒ��/ϟg'E�["+��a�`O�$���G,���/G�Wc������Ƃ`�������eqi� ���U>��KGw�<~:*��sYXX�z� �! <��j�k�5�J��޷��RC�& ���a��&'���%��+�Y�O75�&\��ox�7�TSP*سhlh�,��)�B�d�@��L�v:�<�
�ËA@�+��^�e20��h�Cw�}�L# ����&+�3�y<N��I��6�F��d\�a͵}7��~��$��z?��t#{-lQ�v��,�iC>cl$���b#{Pg'���>
��m��8w)MB�4dt�5۔o��L�pISPd	9K
�\A5�`���dB��-�}R][/�p�d����v�7��E L�t�f��ZI�ژB��ӱ�H�5
�-�h_���M�̮;$p|��p����s�L�	e4 ~maV�ss
P��H�B�=�~���X��5������kE/��pn�@g���Or&a� ����ə��;Y�r8 *	���4X��.T�n�kji��|8)yܜ��E��k�JCB�"�#-�R[���`{�U<�pd�@B��x}�|L��{�%�,`qm�����hҼ�R(�`�K( q��$���`?ï��`���0~LE
��ݹ?,��s��y�a��v������x��1�������ˎ��y�3{ˑ��"R<��!<�������Y�����ί����b�p(�sH<���	XB;%�c��dzj� �V�ܺ}Of0�K�6d�P�x�������3��:�Ze��ݲuۀ l��ܸuG�=}�a7��<3P���p�=���?N����
Cz����:���Ұ�x/��0}�i�a�lZCJ�@��f�3�F,���9.6 Q	L��צ���6�������6�]��h&?75!ܗ;�n���e}iE���D�+[_��O(�?6�b���FN�� ��[����l��w�m_#-ѿ+W�+Ӣ��`*Y�YFҶM�k�m%Z I��HDB�
ц�&ٽo�9xH�l���>;7/	0� ��.��ܢ4��ʙw?�F�¥k2��)
��s���e�y�Iv-��R���*����X��c*��KbR���,�3QB>�2p�lm������k��ʃ��������!ÂK�v`~L��c0����Q��޷Ofgg	�_�z��݋�'O���$[������k���<@1'�/��hC�N	��!�nԃ��p����e&�T0�e:*z?df����
)T�����\�ǵ�U	�p	eHY2U�[R"c�5%�X�@"
��m�&9�G��t� ~%��4�&CJ1�lm�2��gZ�e>����u��6R+��e-�"³>�
`�/��?�� +۱�L%௜�!�2pNɋ	��yٽm�+�.K�S291�b�	m������ŋHf>|����
2e9 ���H`�a!�r�D�Ve��ݔR��`��	t���%9�<O�*@ˎ}nzvF��ڸ�@ {?91E���{��=NM�HKS+�zDݸ{W>�]�ɣ@ol���۟HgO��<.xۡD�AG�?�t�^7��-v�,�7�p���.��a���YYX
�@��R�H���4ڞ�%�!�@qal���u!:=#nr(tX��g'����7�xt��^��n1�G�r�:4��
��D=�<�a��pX�V�� �
�D����6I�x��鐝vN���<��:c��N�΀�9�7�uEAQb<��
�D$�0Ϡ�J4����,Y�$��`EI�6kD�Y|��=�r0�^�d��Θ��{�_�5]�H')��<�3Õ#@�^(�=VU \��?��ÿɤu���́$�1�������#,2�m��E��g�J�Б��5�T�X����l@�;��]���2�8Z��
���$HQ�gr����e�K������TR�IfE�_?gv��t�#�7�;>'��0t��!�޸^�&0�0`��I������=OS�rW"�!zS�X��I��(l�~I�r��b��,���jCg�lh��u��#�*���8��:�C�X���!���B��l͸�����J1�{cc#U&�;� �������JmC=�B,M뉄��g��蘈7��2N��#��Y�C��v>'��a9����޷����$V~���^kjj���پ����7����b,(�)���p���a�����8'K������-��*y�����ƨ�C�� ,<P�ᐸ=Nvd�Qij��-ޖ�[������u�ԥ���0ᯍ����ư+¡�T?z\~�H���' x�@��ֽ�'X�|�.0�Y_^�,����Hsc�465��Z^[�4��1Dه1�>Ȁ�|�p`�*��O�K>�*���e����<?#�ˋ�運�D��
��B#�pMȎ    IDAT��k��X�D:Pj|� +�)g���!-�*�=4JA�Þ�����hQ��8�V�V��ە\�*����ښ45�Ȏ];�Ё��c�n>$�s��O2�����r��5��[���vx�/���1I����:���4CX j*e�~�2���˛���I���2�zn@��o�V Hh�ח	��D!k!�$���:����d��GVVdqq� �@���������<���fW�!�)j��+w��Q[�pX���ǄLp`��pA�Ym=���I���5^AAn�Ʉ���Ǝ�(�K6��RI����x���LJUU� ������M:v��L`s�0��Vy �4���~�`e`;��(s�6�x�2��$��ɣ�qq�#�
��}����f�6BcC�Pc��:��R�*�Z��Z�zx�z�9�>@�
�0��lX���Vؽ���2 ~���\߉��$�ΐM[][��������2??� �ʪ
�4#����`�����K�;�w����AɊ��Z����1 ��t������N�T�n��T2I�= <������չAv������iinП�dh����x�N0�B�7�ɏ�3i�����˹/� cE�^���`��|P��G�V�#:Ni;-V��<s)E�Zn�e�\����ne{�&k�xe��� ��� �UH��g4�"~&;|�b��OZY@�f��`�
Қ�Ϧ�\&^��0�E����4 �0��"k3ӒK�x:�`]��G�YqN�6�� (be2Ɵ?M�Z�(�"�6Yw2k㊇�/v���������_4��AD��b�  $d�g����}B:��)�k�*�MCt*;?���*1��M>�a1�2!PЖ�׎�F1�غ]�����������kaq���n�+�ss�����H�Ng���R�$�wJ$���Fc�:�@����U����q��� �R�83 ȭ6y�T\\9��Z���O�ܿ�?G*��D��H�^/:O��q��s�D�U�,QFc����&����ǽW���i���t��WJ�yα��5����n�����d��R�b	�>����(]�����uYAZu.#�]�����w{�w�����*d��jj�x}𬑵w:%����=Q�r�I0a���
g���	��߁����:ѳ����Qjhj��C�m%���z���E�3��6m�"����-f.M��q䤣�I�k*��K����?Wxr7���!	��_�#���r �<�,F�zDǃ�5�Bp������򊤒��!���F�RU1@�ڨn���	N:S�P/��jI�Sdzf����	҂{�n����p���W��C
,�m�s��UV�M��l#��,0�ٹ�렎0�
�؄�]~T}�$[�� -S��/�C0���ڊ<��:ǁ�����̸=�KN;$��cRWU!-M��3�&�����z�R��5YZ�����`�`QZm���X0S��68����7��*�Fo\���+2�e �Ę��S}Z��+��T���u�ƍ
V�z�=� 6�x:#�x�1��=�o�� �G��;g>`�ȷW����@@<|���PO�,.m8�5X-5��a��5i�o�8ke�t�~7(s[[���<�1��	��m�����˦�����d"%�S�%����Z��������70>�A͑�nhh_ ������Sc���ۼu�D"aʶ�
���}�����@�\+���pQ���'fxȮF���������4��+�G�~_Ue����"�A3���Z�����-j�l�ݝ�Qȩ��;/7\|V��y$��^J4���xVc)I�ݒ�d
�mˢ�n]�U]����o11��ز�.;�L��2���w�ys�|c����R�*>Q��1��w)�3����%{�o���?��$������Dd��#�䣏G8�u�g�՘x�vN0�m�	�|�#��%���=���\[^������J�7�����ŋ�uvw�-����Yd�z��C�f�}~���9|L����$ǉW�PW�{�A�����o/S����S�Ϳ�9dn���Ν���M�et�Z���>�T�
暒�x��_oE��{Ι ��"���L�7_���_�|ô�W�7�tL{K�_�酗?�}!q���� �r�b���C�3eg.���@&�̲����1|%+F~~��ʴ�y!��C����=E� �� ����;�Wp��Q��T�����JmT�^rX�DQ��Ү%I�29^�����۶Ȏ�(��o��;�'�W����~s�����f��H��ųtMB��	](���g�ex�!5ږ���JA|v�����3���8��[��QG��4�s��/-���32��I��`�*� b�k
y	�P�"� ��0@�X_W��}.�յ��F��[ZZ�,�nE��.��E�òZt�@���:�QD�awAv��E�S@fD���0Cx��9�b�����C�ҡ\���� 9�d�G�Q���C;'��lg
U˝後�9" �v �R�3b�������8kP���mm����n �>+Q����e
{c�E�q�'Yv^0C�}�D<�.�u�RS�04\���%) >[ZZ�
��	�,P�1��x<&k���N�<�./�H,絁���`���Ȗ�f���x�ٹ9�kl���V	D*�O�3���/e���$�N����F+எN�]a��D�n��RW%���R:��M6��*��� �/��&�T	7L:L�s��XbTԤS'��O҈tW������Ңģ��)4O�$o:4���Pa����`A�h��n�kmm���n�y�4�6)x��${X[��@��#Y�g%/]<n�5�� �46L���?&��~�����/�dB�f��"(�7��3����iٵ�O�9vX&^>�M�����ȇ �����,Y�HU�����29��%t�6�:@{R:�{a�75��"7s��A>��.�1����0�;�0,T��ë%�&���S����2�>dlx(�tD�i�_]��a �A��e����?����Nr����p�q�(�p��Z��n(���`>Ԗ�:�c�;�03��ۅ����U�3�>
 �M�0ٜ�p�����ih��]�*`h���oe��k~���.ٺu+����Q�٣p�a�υ�g����>(��_�+W�6J�� ��ʅ]6����Ӆ�).�F��޲~8�������ɋW�����-%hd�=^ٸ�_�9$uu����X��q=+**y@���Ņ%�/h��-&б=��S|��{7��1|�9ܜg{�L� $w�?�We9�_�Vrހ�~� �a��XѱՋb�L�&�|��}-b)�l4�b��6��9
3$���jс�-d".�D)ɹ8��?���G����ʦ�"䕽۶��}�e}nJ��Ƙ8Z����%�˭79�
�L{{+�Ǐ�ӽ��A�7�<nYY]��۷8[s��A�L�,��t� A����r��p 	8��~Ǡ9�c0K(&�dhhH�_����/۶ne�* 
�Ύ.�@<�s翦�^ɘ[�ٿ��tuo�[����?����HP�_����+�]꾤�x�W�{�L�q27��q����7����	.��B2cZ���5x����=D���O)�"��˜Yxߋ3���� P�CZI(2����Lp,*��d���8%i�.��`�;��E ?�D� (���@��(x+,&Sb ߜ)||���z�l~�^��1�@�C����&���cr��Q}�X�9��0���>��}{�\>;�����s���3�I:���o�ÑaI%��Ǐ��҃����W_2Q��J�Y�� x��F�C�7\G< #dמ�tcIa߆����s�K2�b��d�g�ڴe3I���E���\766F`f�u[S��}.v� ��C�������<~�\b��q�0���4�U���]�EI&dCO��۽G��eiq�{/ |&��t���/�ϓ9^]]��
vξ��t�B΀�d��Z h�.�r@J��p
FEC.#kP$$�EIIQ�@�(#�a�ȸ���2]��3�oni�@��$Y1����V	Q�}x�G���M���:��#Q�y�ƺ:���H�f/p��B����	~��4OIgk[3�M\��ׯ�i��0��%RI�GE�5)4x� ��#a��xJ]��Z8a�YUS�aw�58��<�����'?��i�T�qP�PNɬK[s��ܲQ6t��;s�K����R�_jooO���}�w�����^�q~��?-��G0�
 ϶�x8����$��k�tT9M�P@��(|`T��H$�	De����$�w����@і>%6Im�)�wd`Fc���@��@%Z��(�P����� b�al�.8�>i	�
	7p}M�`�Q�m�σM�[�R  �xA�oa���5��t4��`�|��%�����ȓ�aٿw�tv�qa��@�!��>�������`{�����R�0y��<�!��eZr��K���ҙ����]j7â��Z�n1�A�'W6F�����K�tpZ���GdU`G��?�����%�g�Vd�ј\�qK^LLI]S��:�.�4��^��w��� %S蚒IU@`���2 �7���G=������P�Bbd@��=JuT� ���"�7S�0�Z�v�K9 @�]�SgN�ᣇdqqY~�����c�VՑJ�(0%,�0���=$2���z8��/^��{�&d���@ ���#����C��F�1�	�9����)�W�˫��_1Cl`��N����μ#�M�F��&�[[W�V>�P0̀��g�ʓ���9�s�����u�g����ɾ�1�-�	��TR���XR.\�&O^MJ����/)�ߝ>zo���>�VRc�,j)�{U$�C�T4�'�t�P��b���-)j���/�u����]���J2��řψ3���_���.����/���˲����cGKG[�<�GJMU��߿_jj��<�B*ٛ����+Ky��ĸ=vP*BA��Ģkd��\��(�s4t�LP[G����8X�2:-����1Ȥ�r��iil"{��������ur��c9��7������)?���Jk[;��s�dn	�j��t���������Z�g?��Ԏ�~ٽH�-��B'�� ��(��в���Ztq!�u
��es��Y�A������au�, E�l�͹C&���+�/�i�s���9�6��u�v.m7�E��e|=e
��h����6��\��$�t���T�L ���d�i踩�biާ�h��MY��g��\/�Mᰜ<yB�'�F���ezr�]B��w�=C��_��@��{�S���w�/\OH�8~�����=�=S`p�냁KXIƅ��8�_�y��ٴe#�r���3X�AB�DcH�H"��_��u��=A��ǏGe}-JY�����( 3�_[S)cO�e~fF��V���7n%p�𱼞���� xJQ�^��?�j���#[gA�y�fٽc��냃2?;'��:�CұuI��H�a����347?C�"X{�\����]�d�{�vAs&G� ,�ul���v���������O:ϤzydW��HyK�>ډ��W%��5�iMs"D{4%EGN����@�	w����P@�{���N"!ttF���D1��=?7�k���-���,�^�����<����d-3$VNM�䒲�`� �� �pV��j�π�u�f���Z$��R�y����bzN�Y���Aʁ�q��~f�$đ^���mr��ٶ�?�s��Dl����}���/�]����Y �}5���+��i))G�S� R<1��/P����Pj��n ۠�f���8�	.k|6M*+��-#c�yП���
�bШ[������{�����:��Q:��-��SĬ�6�_%s
v��ɘ�0�V'��u@�CH�˻�
�c��Dk�-RHq��*����gdu~Zz;Z���=���/d�֍rh���p��x�B�=�gonm%���@�����r��.~l �6�>op�C����c�g��8f�E�\xO,�,�3���0�X{��zM����B����|�C�ю�VI}=7Cx���Y\���;���y=�(u��r��;���!��$��Qn��"���[j*#���#PӞ,/l���\�p>�S>�����,\�a�p�g�}�%4�K��B����&#&>�b��X,J���ɓr��!Y�_�_���2:2�Y�kF�{k�J>L��Q��\�6Ȯ���v��ܹ]Z[����Fꪫ	�т�&lg-�հu�v����K��ʍ[C:��G[P� :7tJGk�6ٴi���/���W� Cɰ�|򉌽� K��<�ۦ�e������_}@�����@]�v�pp�(�:y�غCF�=�ߟ�B��")�yx���WM�Zw��b��q q�p�(��f�A2�˰�B8�!ð��#����[��n0�^2������y�a2-��_�M~�!�Vqq�[�o�g㠕|Fұ5q�R	�@O�l蕅�	�x��i�����ٿou��gg��^�ݽ�-`���"�vn�47�JWg�<z�HnݸN�I�&�e��K>�����a�����AN ��>;Hb �,9X(*C� �g��("���:(���ޥ�7�ҕk��2ס��K�ݿ�9�& �>��3�_^ba�Y�K���̩[	�
\[���M�`x��*����(�d������2�(����NEdh"+�~�Q&(t��\`'>q��� ��U���!���3��k�U�0�"�e�O�L|9X��x�ν..���LZ^�u��
 G,�M8�h!aV���ZeC��ڔ��B��=*#�)/�YD�UV��}@�̃�w	�_�O��ܳge_Ϟ=�/�P P���?�~��Y�����r�"x諯����3��R�  P�ܫTDHF<� ��������E�Ñ���<౏�U�3D����ٲm3�̦�}b�C�L,�6�\���}=|o(�o_�&��ǉu@D:zR**���_���"A(�-���o�h�d
5������-Gbтk�k�l�R'c12�a<�u�RUY)aA`����Y��dSg1T�0d��H\!��d|���� �L�_݊��'#]�ό�F�R!�W���)0#�cw� 1d ��~6�������v�,Q����U:[k����D�TOw7�G ��d�235�rMP�=z<BR���򪬭jכ������|��ڪZ��"� 樭Q�N {��.��]��ei=)�}}IV9I��v#�P%�X��wpEr��RH-�@_��:|P�n�K���K���v'���l٢�����k࿼��������(�&5�V�j9��j�j��~���=Q�A�n�����d�Y��t���\Km[=`P����Hp����Cro�Z,�T]��E}ji�xPT�'b�p7�����G�'�2Xx� �2I���fI+\ ��=���������)���?���l�ٳK��6H*�Gw�db����>n
X H>��34$�n�0�p*�0)<�0��%f�|�3�������]��FT�e����]?%v�85�x�oz�-���c<6l��h�c!4D�#�(8}�K���{r��5x0ﰑDX��o.PB�DA'Y��7JMu%�Cʝ�i������%k�1��[��>�zR�W���Gf���Z.�0�# ���U���
�EJAk�&�oX�567��w�������7�!���	���F}����!�;�����g�������	�0�u�������c�)-!0���w4˩�ǩ���b ���׋V�,x ���Tk:X��:$\���e���\�8d?��oɈ��^ٳsY0�ç<�3��y�Ү,˖�_������)�����=�'�H{O�<x2*�~���r.�{����A2����lX�eȶQ�K�aH�� h��$y�Xvcz�D�    IDAT�����6X��aǿ�����V ����f���`�Ic�Z�ɦn3C���`��MIE�'��u�rF�п�e�PSÔ�Ņ9J���C�K�3��@]������e�~},g?��p���Iʳ����馅g�4�Pt=ε�4g�(���r]�����($a��cf��dṹv����H
LVuKO�F����� f��]���9YZY����ʾ��  {�{Sq�1v���ޒ�3�3/��2jG���L2���E���<{����9�ZL�J;��+^h�LcS� }������/+�A�Fg$�dG��q������lFI��hg� �3�]������>��iw��ryX���Z���ۡs�oJ4����/�v\$�0\}��;r��aJI��1=5EI
~�x�Q�E�1�>���t|Ct�*�� s�0�������t�imo#�Bǈ6ҜqR6�ʮ�Ӻ���'�� ?@���;l���%�&�2�� ��� )��#���s���\�����
	��������N&�F�	�/�Y����CC����'&��q���rj| p��#��4���pI�I@&)�!����
�v�n��(�0�	9�jC莻1H�N} � �8���(��
����?4�
�H��o-:���t؊�Yi�][�V�Cڃ��k�b
��9H��(@�<c$APW`���a� ����x�Tg[�t7�Iow%� ��5=z~�s�(�PȀ=ǹ�6H�p���Fc9:����[=�8��qKE0���^YQA�60�H�Fg	{&�
�MPz��ݺx��L-��'X͙ x;���ފqfץ��I��/;�����l*���ڻ�9�L�j�>�g��v��������bE�*I_þ�@�֕״��`��P�]�9FA�d6q�v	�a�i|�F̼SRY��� �K6��)�l*�4��l�V��2��v\�LJ��x�p1�M}OG�� xL�#���d ��j0�}�J/�LH߆.ٿ{�������ܵ]z�7��~2|_�g�Y⠌TWq#�&��{r���A�<`��$, ��M�l�+jD�0� �wmS[�7]d�s��ʂ��݈̕L*6	[8PWl���`[	t�hC��������$����zT�^�o.��⪴uuˉS����Q���<�a8�
����;w0ZҤ	����Ҫܹ;$k�qٵ�t��q�9tW=yj|���V oT�1̂e���FRą!�U0�KE ��  �� �S}S��8q��� F�������g�S�h\`p��U���{dϮ�:�����;�r�"�buuЍ�2ܞ: ���y���o�����Ɓ~�կ~)W�\�D2U�q�V���~���r���b�����{]�[lm�cG����z�����O����������7���fk�H2���8yL~����P�/�����Ƶ�d��&9����n{��=�������+yoX�
I!�6|&~��WNy&$Cd ���1��@��Y	A�x�d�.B�S��1�-�Ϙ�%i�S���pG���*�ِl��!�?u�&����;n�<��&7�^�BFI��������c��K�� �]]�ܒF�/<�?�g�뵱�VN?,�vo#�����b��p����&����{5����~��A�y�$�ݻ�=��!�75���4��V��9B^�������ـ�{o�&9}�:F`�~v��,��h��E�T��5�{�C�u,�ب
�^�+�⢭di_�C�֐%.�i�76���U<u��0ig<�&�hA����Ca��<n�Z� 1� �@E1�y����9$j�gM
9���~���c���=��v�X��>�Mi�۵��T�J��m�Uic��l���DY��&�����W�F���\��3��yF1����yH:,�{��u���/9(���'�9-�0I��� /��D8k��8B�=>پk��o��kvT�2�`e�{�͛�h����!gN��M}��-��A�k0���ً�2�|\RI��8K��c��a�[Q�e$_ઇp$|^��7ʆ�6�:
�[G#UW�J4&�����f�;@{IB�{���LL�u�8���:~�(��O�����L�#�<R��"a2�0- g��!�zNa�)���<Q�aO "S���)6���>���q�:�@�ܡU x[y�G�7�b+Y�vR�h�܋���˔����a;�<�40����3�T<�ïn>v����P'����^imn��3��6~uu��5�S@�� �XZZ�y�ie%�dXj0���������3	bD��S�	��R�<MH��a}���JT����Ԝ 7"�G�����ZH�xJ����$����[7f���Z�f�cWS���Qf���D�^������6�_�c���,d2: ���5
��0�2-d� k�˴���n���+lĠ)�v�2Y�]}}}k�Q��{-��!������M����!���{�E�M��%┾P"D}���Q;��[ � '�}�Ԅ��I �u�8�i�����.ٵc���׿$�o�V�3S����'��� -�Md���~���у���an&8��M�PM�C�����i[��u�ö`�`���2_oiM� 7ʢ��vJJ�V������I��.&J�r9���'?���*Z� ֚	����XJoߓ�Wn��Ҋ�w�RBS]_/�:/�F�\aS��r��A���%�K����W�.6��KuU�ܹwWfg�e瞽���#�LV�^�A�&����<׍a�h�jb��s��:� ����ԁ��e�Vb�Օ�����}�8,C�ɳ1/�AUv���Ν�y-GFF��ݻl�x5�
�@:-$ <:O`d#!ٷo�:�O�jk�ʕKt�����H�R�m�)�N�#�hB>?��ܹ{O�L�
�1��ρ�~�;���L˵�+�l���U����6������~+Ϟ�iۓ�>:��g˖Mr��	ޓ����7_}I]"F���{wˁ�$��[ȵ[w����"5"��<`<��j��D���+��ؠ��ףI�j�@��*���KV�҇2@M.G�+�3 hY�xlh&XL�w怤��l�0��9���lQ�h�A �`n][	,�r�6�'�h�'`�r���)�bp(A@	�!0V���J(��X_#G�엽�vs`Y ���,��݃�CmXoؤm����
������ߣ�l]��q�⻵���; X:jk�a�ըd1���3Ю��Eڻ:��p��M�5x��h�]	ڎ� $vK3ܟ�����y���AH���b�Ͱ�� 0:vlqE	T��JD�~�P��|XJjѦ���}�G��}� x��[���?����6����e�a��W�><��*�)� qX�LѶ�gQ�����*�".Z��UP_�}��Y��^k�<^�����}=�/�=�̜�`�����(O�p����
)�v��2X�!�pxD�<�Ͻ��~im�P[^S�04
~6˽���g\Sm-��{��|e�s
G���NV�c���L�^�\Ю�ۘ� � L0t�M�-���ܽ��}����65�H*�&�s3�������jbZ�?��hB=�٩�uQ�âӄc�W⢬$�Q�<�Q�=���gerr�{A2�*qX�bR
JC}g��c?�,3��5�>��bQ,[Y�3G-��!�t��	�=���z�E$��qv���IL���UT ΔZ�;J����N2ɡ\qyd� 5�9��3-,~�@p��i�m$��6��Jo[��E"��9k8cyyQ���hN�"-0����]*S� �>30�M��ҝ�A�#��MNOѤ�$��#��2��"� �}!Z΢S[p��2�8��@�����l��+��_˦�������4������˝�af��Qx��]d�p���
["��+��i�p��k4�Կ3"c|�����.p�4��Fk�+N��Y f܌��N��Y�eq�ۯܐʜ#�{�2^Q	����X�U�ap`��9�dlV �x����f˸`#�bu�l���a�ى���.�䏟�N�j��������<~�����= <����<Da�v���Z�v��0]v��逪��%&��������p؃����3>� ([\�����&�]�~Lу�G� �g?����,�`�w ���f�+�V����\�zC^��Ks{���������g��������衃2��%���r��MY��Eb�n�w@��ߗ�C��w�&��EX�ߺ+��n���pK.-�}\v��5Q �[0��Z��@�xO:+'4�5���'���G	�qHܿ��R��R�� �'x��764���	c繑* � �����RLcl�7�ɖ��q����u�2��ganQ�����Icc��<z"/^������TA�������SR�P���CC�¡�c}}�<{�L�>A^��b���x�n�Ť��N��{d�޽\�/]�&{��C�HwO�,��˵[w��	Jg�����!��s�,0��K;O�{Y4�2I$3�ʻ RA�
����Ϧ��n���4�UK6�\��01�TZ���1�ݢ�㣶�����!a�"�G7~:sa��Āk��{�
|�ˑg��yŏs0���2f/����$EvQG�Qs�?�s+e�a��޽;e��m<X��`�d�W,�ՙ|����{Q���S�d9z��ƙ�������D���\����7�ǲ+#��t��5ì
hH&�D;D>S*��M
 v�H��*p4��t)I u�)I�pVX��t-�|��02Ƿ�u����S�+x�s�h?���O�;�H4��e�K�~9�/'U��4ޏq!C�=}��_Ϝw��S�nR.4�3j}�v���O��:�VMd����E�>�(�� �u1��v��z�6ܲ2��7�U�J��Zٷg�D�A���,(
O xXF�|��\$����@����zn~^0�I�δW~5!��\��u�"BY���q��a)�0$f+�|������2��9e�յ��m�v��k��/'���q����n��� #���ݻw�LC���7�N$4W���2!}}�,>�S�o]��Lg
R�� {o0,��\�W�3�`��\��{Lb$���CI
`�c�
��$�o+�t<�-\f ]�����[�����eg�sag� i�s�N�9�;�N]݊>�r=�W���WW��$W��]K�줴/'�x���؃⩤�A�`��d"���4�/�� T 8��N�8����k{#��e�yX�@&3Hw ���"�6�>��?�⚂á�:h�I�&����r�m[�P�Ć;�gϟ�x�^�����;ǋ�벎 B�pi�8W@Itx0��s˖�>9}��w�K6*d�ə-|�?e#�����ܵ���+<�h90�.�BA�ƴBנN�pD�ah��bl�OIf-Uw
D��Wi�3����J#9E�j�~��V�[[��-y��{�z
�&ck�O�Ł���M>rq����`�N,4g�ɴa���� x�������.:Z����Ɔ:9}�z܎�Ƀ{wY-�����m�Ƞ�yE�,, ��,9�V �|���,�{--�/g�ri+I
ʴ��
6�C����O����ˎ����,���sJf&'�8�^d�9����鑇�_ȷ׮���Ein��!Ө��#Ɠ���NM
UpX�����oޔ��Y���=&�7o���_����.�w��Է�ɵ��d��-�Br�.��}�eg�:��u��7ڒox0�~��� �������V���bDeghW w�[��=���`ˡ�䡔�T|�.G��� �^c�kh�]�6�wN��|ZF�<�H�Bz7t�֙�]�]�.>��s+� S����'{��V���#n�ݝ�ic/$�ש����<x$c�_J.���+X+��0�㒎�2�s�����"���F"U���ӳ��$\W/�P�8�~I�����#y�E �Lp�{	v!��u5���9�t�^7�K��x9��h���JV2�$�#�t}��Ǟ���a��y^��3�Y�l&��`A�'�3��곇~t.����vAqA��X��|�����!����s��p���gp�y�?޴��]�ra����@�&.�JjP��M&&a�e9(1�<�W��-c��t|b�]��vTc ���Y��z���A2�4������K��Y�J >��]�hݶ�L�d١�� ��CHi\^�xC!u��T��J�e����oX��=���y������_o��:t��ڭ�5ƾ��,�g���(���ׁ�g�AH �v_�>�^d�	�KZx��O�r ����itx�5Y_��4�!�X��~L>���(O�
���)�H;O � �����0_��V��n�D�cY�s�G��-����<t�.�?t�ϼ/�õ�m�ٲi��U���V�e�6�=~(��g�$�3-��0�'���#T�r��1����W.��GY4��ձ(��~�����{v���4���r?ܵ}�ttm �t��-��=]�������k2=���
|ܽ�	���^%��`�[�;g{�Ql�b�4��4�	��`�q��9
���������wa���ʊ��� �� Z����夺R�H�l�����8ɡɣ�<Ğ���IF�ݣ��E3�9CNv�v��J���x�4(�t)A@T"���B:/
{ɱ�P]�A������þ��H`�10J"�ᐊ@��;��iXv2,�+��U�Ɠ	�8� C¯�4��X��*T-^��TgAM���O �(0�z6ЋL~C}����RF���5�O��)�av�	��p�4��1��E� A�����p�M���(~��H�?{�����zeK��ן�����r���S��	� �7 ��0��Vm$f�ǭ6�K, Ve,�Ҥ�R��)�o��K�\�A��=��[��CL��[A��j�E� x �����KD�Y��&�b�Afd�9�G V&H �
������2ޱ��l���+���.]m�r��yij��t<�g�^?���Uj��|"���O�<�_��{�ԭ�ye�)�b�*g4�Aׇ�|�(�{��K켲O�Q�V�h}E�ʼv�ռ/7S
 �չF�r��0�������3�	�J:!�L��z蕑�1�4xKf�W���[�y�=����K����|���"�ղ{�N��꒙I �[ԵUWD���<080��Y��y�}ij������w� �x��<��oY �!0������6�y�ld����"�������Pȕ%�},ɋ�		E*�����xnD�yb�3�RF71 2D!�$�7=��aQ
F���C��\Ŧ�H� O7=�9���8�~�L�n������Ў�5����*굱���L��.�i�
�(�F�Ӝ&�B�SS#�U!2�6���6���N�����DR�e)����z_� >E��H��H�q�y���[�ƥ��E�V㲸'͡�M����Ok�~i�����J��������tjqY^��3I/�N�	0�8���� ��bl�H��`�l(���A��[`���{��<.MM��¬T�R��(��zev� Ƣ�0?/^0���@�B�[HqrZ���`�/��y�ڡA�%�hw0z�,�yq p�����m&�'�Wx���f�+<cXs���<`�P��K�w�������
�t1��2|6���,��1��	�ć $�(�2�$jO� V�+�)������|1x�8�c��F��3�xp�L&e���y��H?x�Z�0R/���%-��y�*����"�m�BJb�:�m/���a�}�|1T���k�� ^m��c�&����<�)�qH��� d���{��,謫����	���=����;g(�����b�x�T+�w�?x�6��._���s��a>/8�`3���ݻw��c�ء;��Wr���>O���Gѭ�L�    IDAT��%������
<+����=ԅ��,����3�r��=YY�1ͽ��S���-���`$����%�����cy�h�{fC��v�5K�������l�3Ͳ�nzW�Y�
@�<P�}zz��ẘ3�Kc�oP��>H�RP;���%FP��f�fz�ah�F�{��WVz��s�s�|��&&�Q&+��}���{��.��J�\�X*-�HBn?�/W��&2�AwN ��JG�D���z���w�׎%���u���ZxL�a8<�K���$zmnfA�����$_@0��H$2f��P�x �	��{0���IOO�c܍�a�o\�0���r�δ�L
�^.��^���$aw��ٔf;�L�O����xG� �!��B�ft��}X���D�$P�k�Y�����k�y���+y�xR���A��_��aUiD#۸�h(F�������YM�tT/Q�x�<�\��	ABpM�Ĥ�u�헵�6H���q�M߱�$c!Y54 ���dx�O{3/������UO���2���?=���_�b��>^n�(�����&�2pױ����C��MЭ�L�u�[�O���%h��st��ps��:(���/-�S��L%�C�V���n*��d�r=oԶ�;�I<�7�tyC@�@�ڠ���0 �1�K��{��?v�'F�w@���{�fn��|"[��ɖ�1�t����P�bzJ�\��&/����C��b�9m���{��U�k ����ef��I���>����(p/� ���U-L��[��S�;HY=����<A�� �9��l������$�>,th�W��I�X+�@$)7�<��_�#�_�i����Ѐ�8uJn߽Á(y��ee��=�c�F�.\</K�9�$S��۱u���'OK��O��?��5c��ﾐ��\%h`$ {�{B��W:Ԓ t�ߖ�����ٓ9$��3���'����tI �N�����L�`,!C����Mτ�M��k�Q,�J��xT���edhP�f�����L�%�M�Md(*��^�݀�/=���Hz�mӞ���ҴT)��E��Дzx`P���O�>�&k�9&Q�e7k�{��A�����C���Q��؞�U���R�*�^��7�H8��6Xݰ6��HF#����K$���sy��[����RA�*���vl#��t��O��U�d�{�q߸N�����'����L��������	Ǩg�8�&��xf�_���g�)=�ʧ���y0��F@��58d�S�p.D�� �}�u�d��^8|��275��h�ƐP�H� ��.��,Y'�GUR
�AȂￖ�i�O�L+6���V�,�W]:��4��RIi��*��D�,���m4�85#�<�C|��0����@�k����-�K�%��/V-�쩾V5xZ-5��5��=�'�V�w����g��]�n��$�Au>�T8�5�J:R��.�w�
iMT=滲mc:i���Pw�P�
'�s=���\ 27~] ��>�'p�"$43Ҩ @��s��]�k`�}r�4�{��?�ɤtji#�&�A�58��g⳿��gC+��VX���ؙS����S��@<@$�0�/&�BZ��̥ q���m[wH���ܾs��sT�ٌ�l1q�:	8@o4�`"��ޘf�F&z��m�s�6I�d�qMK9�s﮼���j���ڰaS�8�p���NU}��I76��B)����X		���s�w�������A�l�h� �F#'�3U)�ؽS�8vL8G}-�X\ڍ
[�ᐇ}����l'¢�fk ���`H֌���G��� I <��!����>�`�Sp^�r�� ɇ��hĖ�xTw����������61\[м
'+�C<�T���mN0G�u��{ �مE����dJ��`7U��p���΢���Y�3�,<o�+T8y�P����ɡ�)�}�UBH�����o�3aL�Fd��� #Qꇅu"��VX*Rj��A�`J9z�0/d!z���F�'��r�D,(��iɦRҟI����b&���PP���К��� ��gw~|��/
���B���F���T㌋Ĉ�:�0�šT�ZTB��v��"@t���Ć#�<�Qnˏ�7�y��Ӹ;h���8a�`S�"��( R�i:	����9�� >$��i�
� W0+�p����O��}c�T(̦y�愮)�>��w�@�*��ʞ�[d|�j���s28�G���4x�ذ����p��ݴ)������ɓ'��U0�q����zv��Y�������&�a�c���< 	��--��>{l�sp,��� ��R����v�����~� �r \Ӛ5c<Љ^��$��G�f��Wez!/�׭�w�=.#������F`���9v��O ��Ϝa� ���C�ӧ���dptX����K��*�����d� �h`Q��w�\�� �����IRߖJ� ��I��<�y��v�p�ʍ��I���н�.O�Q���jy%	�cM	���}��Az~��<���g�_�	�=�c�'+;v�U#����G�g�n�RV�4��{��$z�{�lٶU��������x� � �۷n�uck�:\�xE�N>�A����x�����;rX~���h#���:-��	HIʍ�|s���_���R=��H#�֎�k`��P�fe�بt�ey��!�;C�ÒH�%��Jn��I�Jx��U�xud�/#�Fe�7��u��\^&�f��lN��U)��ͫ��rML`L �1�%�HK��CB�p��3��(�k�jH2��J9/�XD��I).��䓇�$���K �'���%��܋2T(y�]���ZãWi\��v��\%"/�Pm3�9zx�dT����E$��R���~�(���\CS�̜D1l���c����X�צً6t��A	����c�0��x�:>�Ii��
%x��@���c����f׭	p��{	�v4]��M�5��b���l�V��id�t������z��TaT�������Xti{)�3;lX��������FNq�!4��,MOI�R�.:����fe�p�B*h�V$��#�T/�F� �� T�;�d���|��!��X7�s��[�c?x���`KAX���qX#XJN��D8�q�\V����P0��ψS���7Y�$2=���NNaI�����C`du'�|)O��T �}!�:k���O�8������PΊ���rT�(]Ԟ8���P���X*J	��H� �k�i��s�I�8�\�h�ߡ�"�'� L��5�C�9L�G�F�f����!�d4�{r6�T*F ��Nę%�y�����c�qëx�� ���>��b�\k���B�}l����F��-�7��o��?C��2Nks�3=)ꩄ��Z-##Cl�� ɚ�W�gٰ�}�2"G���f�L��E���x��%�i�`�>cM���A�H2���� �㞂0�]��mۥXn�@L7�D�*�+b�7��M)�d���Į� �PQ1_��w��{������N�H��B ���r�,�-$\������uk�7�#�=�f_&�e:��FF֟��9ѼRBc�B�u�T��Mz^I42�j��Yps�>�p���"Vj�;��^�p��f�~�M� �e��bv!��h��$ms�I���-7T�,�s�X�l���@�.@u���I	l�.����!��{:�z�P8΃��=�C�cz��ݻ$ت���cپe��d���Z�_���ɓ�d$�Cf�I	�=7o*��v��zȘ��%E�:�� �_�����1w;�����1Tf`�6�ߪU���Z�X��#�����'��!�ӷ�C����>���݉r��6�U0|�'M��;�SBs	^�K��n�9r�d39yꔜ>}Fva����J,��3/ю�EH$ZA��,�:Q�MؤNL'慂IB: �/Jia^R`-���"�%:Zq~��`G5��21���.��d����6���}�ҮW٨�`y�ݷd���d|�s��Du�<������W�ON�W�ϱ����s�'�4�q��wޠ^�X���,�����8�#�JUn^�%'O�AN��	M���x�u����Y����+UO76 ��ȍ{w�/�tbq��{��.�98�ՔL"*������R.I�I�?�U[R,T�ϊJ�5�O0�8��Þ��	�W��Jo:�kZX\���\��&�g�֕ �`J����&K��xJe4�.����B>�ׁ�a ��#!�+4��g8h�XX���z��&�4�45+a��C]3Kcdm,2|�{��9�@�R���{'[l�d� �n�>�xoVB�'��=Y�N>��4_����fD�K��[�[��h�MP-�l"�mH��1I����k�A��U\̽���M3�ă�\?��0��O
�=@Ό�u��TTP���/~ƯEfܲ!o��ņe�)O�C,�泀d%�CZ< ��V՘`�}�R��;ݟ���9�h�d�`ۣ��� ��E�FP�Q	�TPM��g0�x2٨����4�I���zT���*IPn9և%v�H��j<N�F��H�9�J ,|!D9�#� �Cu	׃�B8�[�,���3` �� Ir��>����v$\m��xr�P1�u��Pq�Cv�霰���nHrլA��p�4���Sgg�́�$���R��;�qOAH�g5|�:@�
�����e�T���v������0� ��h0,=�!GU4�K__�d~UI��D4*G���[7�����Y�ԟ>��I�%��� 5����l�9��h��2޸aG�>�ꚺ 1r(����{)�D��
�n�OAX>~�d^�\�!��J��A^đ�$dxx��q�dV�[�;�����#O�ߘ	����P5��� ���"�~v�52�j�d�C$fA`�U�sxskֆ��rR�a�"��M�9�'�w� �(��]�v����/ج��A� ��Ɛ ��&�u�Fڎc���l2�����_�[7���6-��� ��|rf�G�/�b�X{������բt�,Uhۇ�ƍf�SC�p��fy�u `R��HP�EWr���>f�xHF8a��0)��{����s,>,F<P4x�Ee�(��И�DvG������<l�4��t�ɯ] ��+Ld��#˓HH:2��ʁ�;�����6.c#r��ٷg���]������\��5�������raߢK�r��u����A}��.�����Y���r,3p[J��O�KM�71�11���U �ɖ�X�f�����~�Sz��}����[��Z�j# �HB��~(_��J��2�a\~��9H���>�[w�Rt���޾:�w7K�Ȁ뵊�f�b�/^����Ds�7d��>2�_Lɍ;w����2��K+h�J�P���E�c��� ������2v�.#�w�k`�عg�r��\���P"d��w�~S<@�z��R*4��h8��!#�-ꥯ��;�p_c��ehՐ�u�]9~�-�w�B��s���cT-��!�9}�+���/ ��A�w�z[~������S'���G�X`��j#��c)Y,����lb��J]B���8 ӣ\��J6���f��G�I4 (q0� Wp`��%��8�d8$��YDB��s��Ō,��R��<�V���5��VKb���j��<�� �`%�5j���������IH�'!�B��q�� ��}1���	��д�+և!k�i�eM��NG�H��B��	K"�'!$WhT��4����
E��Lq�G\y� |S]�B�B��H��'z��k��x�Z�{����U�&��9�0�i��̚��ʈ���D@�I#$���:Яl�V:	�8p�ˎ[��=	&_�[�����>�zX�w���k��w��&3 �����}���I�D�ĪV$7�B*�es7ln� ��$���f;�F�E����J�o�q�_p�"�Յ��3��y
h	��H�zvPf�g�_�h� mMz�UJ��:j�ؖ$%��j��0s�dYf?�3��]�1�%
�	Ϝ��V)�)�N;MH�Ba)Ud��YLrff�Z�Ҵ*�FGZWkB_��^7�K4jw0�H�d�/�T[�b����ᖉO��5��>�� R�O?�����0mV+�AJ�;�8��-�I�^�x4"�j��a|�zY52��ݽ��.`�? '+5�'�.$v��JV��cP�� ��ϊ}��8���S8�{�>��Q�G��3TH�&��s$B����Ie�s��Ge�m/��
B8B
�G��[$��f 1լ�g ����N8�J	�k��ծk.>fR���Q�D�ɸ r$3�.�.��+��ڵ�Y�s�Yzܿ�TO�/	6�xHvl����i�� ��������##c�y~����g���l�B �F`xcP��ԩJE��<�?0�(Qa��z�i��!+�6|�� Nd�5V��tܓNJ4�`���c<�hLG�ss�}C����X�R�%;��jq�0�OM� �m��7vr9z�jI�ł��}b-r`
��Mh�� �,M6t���@_�ܷ�����έ�}�Fy��l۲YFFy]��.^����zbF9��߼�<$6髖u:�]�����\����?m�b���������?-�ud��ɒ��
d� �M#��2 ��M x��zz$�K_��#)iJX��~WN~y^�󘠺^>��X����)�v��&1��K�}�f��d(9 ��i�����GvN�f#k�іB�"?�k�n����o̎N�GG�q䁫��S/�$,�ڐ�(�2 ����l��=O
E ��K4�v��j/�=�>/�J�;�!�v�fE���[\_�x�A����`��h,*ʋ�YN��R/�/��C���!9z옴�m�}.4y2<�8�ۭ:�/��bI�fs<��6a7�)
�f�-���Ⱦ�2?=Ŧ�b)�w����(5c�e'�b; ��aI�H=�J�#ULWEɞCXkL�c�d�9�L�-$3��4����0Q "Z�&th@��*��TP*�kD���8�5��7� ���}��k���P��$' BQM��8%�`Q�9��zM�=�(8���ê����m��� �	���ʷ���}�G,<�g4�!�"�	K3��&�@�O� ���oR��&��7�}|�is�R�k��K"��dke���=S�0a'�`�B��>>����lR�Pell��8����)���k�9�5;�$�ևf[HE�0ɀ���ϕ}[�R�<�L��_�1�.ui�K@��n.X���5�z�c����_�r�E���g��M$�{�y#�3*ظ�Jr"-�L�V����W�
VN�g�.�s �\E���8��1�X�䩑v�;�3�)zI�Sms�n$,��ҹ.yQw+��2)�I@9�Ƚ��rq��Qo }���df�q\c�.]"���>b3���<�%W)!XI�և�4
���[\���4�pI��J}ֱ�Z-��V�J����C������� 33SL�@P�C�u��#������aJp�2��n�<�x�.YQ�lBB�Y|@��u���`�������rw��� T�׀��T����j�4�~1v�����냔U�AV0e��T�{B��x����)H��$pa^p������f ֻh�׳�u@�%T;>�*ޏ9]a�;�ׅw�B�������*�����B�~����C���	�fHS�1 ڑ4��U+ɤ�2�q���<.ٞ��q�����D,��{�F�ltt����������l�z��
uT m�X��Nm�$�9�x��3ܤB�̩^,[���C��7@ ��C:�WK����%y15������7GX�7��������>��b�7��6mX�gc��<�M�T��1�M8|����1�Р��_0�;� ����s/�Ȧ��e��r��5j��a�	S������B�c�v�o �۷�ʉS'���;ڼ�|���>{�������    IDAT��� 7��*d6���j�>w�߱��nL��hA
�"�����1�[�L� �d�z w��I�������������2:�^���xȟ:��\�uS*X�i�8���@�$�!Ԁ��q�HuH�y��+�d����՚,a
e�̒2J�<�0-�Y����r�kF95�;�ۜd	��T �����_^��?�J���|l�%���z��hL��{�-N��@�M��Kni^�|}Q�?Ƥ���dr� ��&�x������D6�	��D�"&��;:���f���-�le�:Xn�'��E`D+ �6���� 9z� i'�1�V0, �J�CҊ$��ʀ����j�y��h�lԽAdfFo)��ڄ�%�	 �	�%L�W���`(��$ z^;�*>�F\h�yX5���q���M�� ��eC�k�1�&F�D�rYf�M�< ������'�貾��z�H����k��~�xHL0�G��N�o���p��*�k� 1@οj�R�>��>�n-����` ���c�C���{�Lb8X��&_N�`���o�h�i�Fz��E����7���^�0)HE�2Y[�;�?DU9PCq0��@R�b<c6�9��@��E�xN�j���v`��m��ׇ|	�'��$_V�.�%Ì�n �(ah�!i�09��5AEb�1�́8��*M�ޯq���z�j���8J�~�_�4b�X4��@ �`&��s�n�1 ����6��'��@&�7s�-j�w�% �`as��0>{V0�?+�L�TR�{�R4~c���'04r�:�%�!jJa������g��I�Ԅת%H��-�˘��麿q��MF��ͅ0y�Y1��@]|j�%�׎���˳���_�]q��k3|��A����.��QMZ3�Z�{�r��7���c�Vz�C�M��1�*W�j�u�m�,P���;8�Q
ׂ� ��[��f��@�R(%��z| �&��
�C��`Q�J	�TȤ�3��Y� ���m���8����<�<�KV��[c�*��ֵ�6����Z�Z �0Y��Y�T���r�>{f��;��L:��H7�Pa�1.�~p���h��h\"Ѹ�)��[R6!c��d󺵒�$%�:��h,��T:��lٲ�����������~1S�����v[��Zզ���7�����"o|����kti�5%���y�C��� �개	 ?2:$�׬e�z69I{E��͋�>�zsx�Y�у��}1'�j�~��i���֮���cZV���%�ù%�j� ezv��F�@��,Š��.�� ����B���d�ݑ�{(�A�u:�"�??7'�3�\d�m��,4�-Pz��m.Zr����|�+�O{���dt�P&Z���(4�p��˖X�i��%[]6ZJ��`�'BI�������o�;~o�bM6o�)�fH�_�FO�����w�����ėg�����;�����^\3z��ƽD C ������g�ʉ�ˬQ�@<}��S�j
	[�-�b�� ���I���&�����w%�������^�@�xN`������H�@�~��VM��E>�Z���EרC/n�o7��;VL�EW6K�|�H�:�pFBnf�������el8��, �,�׃`2�VCC�0�tAN �x��j]ꐨ�3�3�Jj��T8��+5�APK���������1�vL��%����	�R���!M0@���{k��8����(�3dg;��q���9y@�MɵǨϷ����HxBt�i��2���$�^��l���{��s�z�2�x|�=.g�C�u]�U�|�`JrDex�@s�q� �����yx�j�t?��0l<{z���F�SNER�]�ܾ$�����ܴ��0My�����h÷o�C{�H_���% uVW U��bS=�݁0`F�ކ���uD}�Rc���u���z:�8�F���	K��!y=�G�\��׎�H��~7!�+T�Ba�&�~��Q�5�g��)z~S��:d�h�� B�ࢦ�0��:�%>��۽`?M x�N���9�A���d�!mP��+���$�l"��A2]g
�(�#��?Lf����Pq�zPT!��@��q̈ �В���䃓���'��o���9$����>.@w]��m�����D�a��Ť��
�B2�C �&�oW����r��y����_��LM?c��44�Ø F��!���>$8���mz�8�� ���%6`�Q�@�$ �w9U�A�^�:��m�T������Ѹ[k�h�	��FU��PP�Ml-�A�o�-����>K��]�xkI�+%*~�I�Iy(�A�v��:�q�^_ce86]�n�`�u�c��g�7��ֹ�������hϑ�$����Q4�NxϠ����22�+�dTFze�Ρ��fRH�
�H�t���a�֛��v�� �g��w��4�Z	��2�Y�n�@��f���k6�P.�MX"JK�=Ak��P�DpFV	oց��syN`CK���BS^�����T��g,(G�jzv���8k`�ߧ^q��h 4"�׋�e<XWͮ��J@IZ`�R=|pl��G��P�)/ߓ����ߺq����IrSB;�@�5�o xh��db.4�n+O��k�m���db�A���e��g�e����]3���8�T>�x,t<|�d8�]���u	����� <�����e ��<��BYv�9 �P\�]�"S��?���l����Y�q�� �	��\s�"�\����r&��dP��R,$$�W04*��l�������ѿ�P$������|�E7��uw�t�ޫ��{&� �>����f���6t8�c��_�]���"A7'��
�j���d�u�RH��L �4$�=D`y����A�~�H@Z��g�Q.H���$TL�,W�Zp�U���!�������e���<�'K�����m� �����w�<��\A�}��Z-�v��o�W�ˀ+nT�_��k�f ��>�MT�WݼT���i��E�'���i�,�Ԯ��p���;�W;[ҕ��2�-�.�%Na�$�2?&V�I^1ÿ4	���}�"B�a@�k�9� �h���!i��f� ߊ*���i���ޔ�R����'s����]��=��D�� ��pw3M��Jo�1fGL!1sx�X�a|h�\�jD�z�l۸Q:�{a�,�Q݄�^�	��a��'��q��J�L}	�պ^-*��	J�v�|O:�þr�k��0T��&Q�V����MP�v�7�u�)��P'Vk���j�9�-���9#2_C�עhPFS�o��`�=͸:EY� :l�3X�8�2�a4�boC�م2�X+Ի7a>��$�#��Ga�dW�0Ѓ�S7��+i��u_��{� 5I�Q�F�{��F�j�H������KE;� d�HK�E(���8?���J�1f��X�~��ӭ�� ��?��Z��Ү������=�b�����<<�AZ ��a���hL�2YY5<"۷o�'���N9��Q^��[o��� �	�WR�8�:z����W�#�*�;��
�N�A����rU�M7���Tj��� ��>ir��dn%\�
)'t���eb���w	�K���ҔR�A��3b�ŞbV����Z�Z���Z����N
����̱𠉇D����J Έ��7t��z� 9�/�.�(��Dex�_֯�!�'�%�'���e������.3|띻/�돾�����b�\;^n�m�h[�j�,�b�M�`��`�Ҩ�\f��aM-{*��o�ܩl/�����i���<� �C��nt2,�|�-��B``��E% ӛ��k��p�)L�>:�hIͯUP�,��ąM[)�O;.����s	4�`�$�XD3���5�e�Ⱦ		[2����1.۷ʅs�莒�F2�A�����֒[�l�&�����p�������f%�g&�
�8[���`��g���<�0X�BP���p���(-q��Se>���A�������L	�HP`��\�z�ܽwO&��d�������[29� ��V����љ��s��������邁	Cr�6;�V�>�t`�����7Gځ���<ʫ(qP���l���C�x��Cs��G� �z*��*�K�N�	߳&�������N��ge���?�����S�C5H}8�]�V��~P2??O���sx=��'z�R.Uev~^rh�,�(%j�"K"I�N�;��ch���]��¼��_H%���xeƜN0$�����#�vnc�&*J��]���YeT���/��r�&'�]�s�.K;�D��԰��1:ѨW��j>��Ҭ�X�dϡ��S@��/a;ג6��X�AI�M�AXЩk�6�iS���
^4�q~�?�vrs�o`���c����x�sY)����;
���l�%��b��b�wq����9�XN]h�����pM�f%Г�6<±N�۔1�- ��I�o��8 orX�h�P^��
&�Ԇ%���$A�@��.9�J��p@��Z�i�/>�b}{�&�d\�:zH�~����s��*��,Ƀѥ6ڦ�v�<�C, b�& �R���$��>W�N��5�ĉ=�e6�"�j�1[�LL��u�����.�JR�UF�5��J�8�@�~ېͅ01;�T�aCbI6�i�r�?NR�
Mpև%q֍��MKP}H��wI���Q�=T>��S��ʲ�����ב��h)�sc�T�S�q�j�UJաm"�>�"AI�S��#���g)_X�v�d����\�@�R�Fy*Q	�G{��ں�LO��l���t	�K,p/M1�� 1�$�ة�����r��^��|*���V��&�r�D
�7 ���b4&�~Y�zT�m�,�oߔ��o�� ��g?�Cʓ�`�Y�|�qN`���=H�����e�ʍ�]�K�>��2���L�~��:�2W$XM�[ݧ ���5�r��Dq�I���> ��q���>PYOw�d����yik��	�c�m}���UD��n2c���a%bO�y�
��L��Q�$S\=��D]���c&~��k2�P����#�L�%��I�P���d.����ϫ�n��ƍ�/��/�"�F ��/f���J�@�ى�U)��Z*KZ5�f��Q��d���ɴ.p��g@.0;��&���w����Hr g�248z��1/X��ŀ�taa��f��W�R�v-9��i�t(�juQ�FcV�Ug��v�kVm�md�hI�w6��R�)�b�a JoZ���!�/�Ȟ�-2�nL.]<î{4� 8"� .�xzx�b�[$������r��i�~��Ĩ�m+!����VHh�����yo��ҏ���]=�ix_�=f���C���t|��G���i	 ��C7n� �RE&�g�������i���GHiǩ��˕��ށPT:��tl�mVu
reP�e�2:�Z4�h����J�u�8��;�P��69B�TXr��k����e�잛�N��:H�	&�����Sa��� U0sj5*�ۛ��[6ѦtazZ>�O�[���Sɴ���'ܝ��ܽ{_�h���41m.��k����e|�*y��\���'���郱>V5��G�O�g{�ՔM����}G&vmguj~aV�]� _�<���M�9���|A>��y:�(�T�4��` S8�Gu24��L�u}�R xO��M�Xm@�5���i?K[��c��{ښ�  `2�/��{A( p*�4nT�`���@�'��r��!^D�I�RYZ���%�5�h��H�Ufe�6&Ȇ�p^�K�ф��1p��Յ"��G���U�v��
I��W��>)��+���jc���F�BA3�%
�N81�kB��7u���ɓ�H��]^<;��]���;	�����7��RN�������d*�ʞ]��؁��E������3��������bxUEW����^2��+k�sƱ���w�>��N���G����?���Gw�}����XLj�]c}5_���<��4������Xo�/����
J"�+�tZ�p��IP�1XC�7$1�g�w��a,]!��>���0ީ��;s|�޿o�M�C����/8�t��=�ߦ�}1!c�K'"#y ��d��߰j޼e}�>|,w�=���E��@��Դ�(�9���C��d]ViC��|��l�y�w����}9U/� ���ΠW��佷ސ��˓�w���/$��g��: ���HH*�]#���������h��j�db������s�`j�2�WQ�h��%�Jd�c�i��� �v�Ƶa���M`�)̴vuUSs��Oq��3�k��d[��ĀN��GcI ֺ�w�t����5���%C,A��d��v��$�V0"��=3��M�ʰ5�A�+�5���֓�t�xTu@����o�á��`%@�]��������}㦉�}����دx� �9{�����rSB�&�6 �2�\G�g�e�&<;� '���R	%�j#~�[>��s6��������1+�"{Զ@JP�@� `�Cd��Y��t6�l;c��Ǫ�@qd����5��Ӝ�W:�j�M'2t�'Rp��R��;mNY4 �4�\����ANg�<!KK�R���FKsie���{���:l�gϞ���w��7o�z�Q�i��f%�g }~�,_�|=�����2@��<�T�A��AI�K�,ѲM��ɟ����3�8ݿ��@�e�fz�.�%�镫��ʧ����Œl������Ri��>{N.ߺC �F���a��vXo]�JҜ^��ɴ���X;/�t@r���������KR\X�(&���� ~�C���w¬A�4���kb}%��|�c�6��=�o��v�������+r��y��7Y���KHh�����s��o'�1�<�pt� �8��h���2�k����{�ZX������K���Iiw��'@ ʣ�ݥp�ׯY-�{���߷�l2*gS33r���{����>p�>zLF׬g��ե�Rl�o��L���yH��ϱ��֡D��m_�}�z����l���j�CV{X�k�1T�3�x vhj=�-��8�0vdwH(��c�XS,���x��ۘwNE��p�Zʹ��>���Z*�}�DF��;l�����4��~ w\X�/�U�v��G��a$s�!iaJ/�7dX��\� Ȏ���2 O��7	�8<����9�w���!�kb�Ih�ܮr*V��a���p�*SZ�aͨ|��d�Ȉܿu]Ο�R槧i�FB%o�=���5�u�����H2�n?w������%~� ��H�O�Fr�;{I{��H(]�0�4zڜ�Z+	�ai���E��ݖ6'ҁ
RO�q9]1\�RJA�7��c��f{��i��f����&���
悗i�YQ\໯aɈ�͎l/����L�\���"&�����8����HM����9��70({���tpL��~��<~�� ����S^�G��/9`�c���4@���] or�Wr�j�$W��x��].I�����;r��~yx��կ���H���C���$��M���߰N������0^��=!��{�v�pa�}����@1%��lk/�&h�
/׫3y��ij	��~�:�{�Y��$�L�\�������MZ�J9OI��Z{U'C�l9�җU'm�>�'������cB�
㠏�Ģפҿ�mr-z���B�+�J^�zT$$�p�c���u@�x���'M���"!آa#V���V�Z���ٲe�ڷ���[�RSB�FPj���0¶֤fK���%Lf���y����v�Sz��IJ���������EY�f�x}�z0C�����#i��,�e`�ɛZ�6Y��l.Ӄ������Dp�W��
��tՖP�Ӽ: ϲi"%�XJ.�)����=��M�SO���C�dۖq9{椼���\n���?~(ý�7�g�>ٶm*��?��s���1�d��р�\�e��e۾p���    IDAT��= _�A�4�������5
[�����-�����QB�����q�HXз�R\�T#�?��|��)��-ɶ]���P*��|y���![O7�>S��l��F&����&�i2�	�0�3�`�L��a4@� ��٤�}�����-�x����)g{�l֘�>^-k�B{� z �f`-���E������{w�ݷߑ������dvf^��EY;��ҙ�>�T��r��^�L�&�XT�=�БT2!�N��GK_*)S����ŋr��y��9-�ԵAA2ʫ��Ĕ�w�yS���![��^��ܢ���?�.	;w�אhl�&g/\��N��r�#�TVj�B��j�	�ij8����e+8�p��xñ��B+ �s_����ըJ$ؑR~�^�A0��?סb��='0�q�o�t��b�4�VD��&@g33�*]ӕ�����K=��땥%�C���w9�Wi���E���ؤ_l��[�N,)�v�P�d��� �X�F��X_�4 �R)��q��C�`�>�\bH| ������f 5g��H�S	��2d�q��Y�d�m_;�4���i������d `��^�2�K'b�����{��e�}�B�M<g�{�J�>��9)#�̳U%	���j�>���{����!�4�Rϓ��*�xl��m���?���җ�k�F��(U(O�nA V$�Z��5�Uc�꼁<פ�#qu�b�$�˵��*�}:x�`�7�No�:��ժ�}6^��β�+���Hjډ���ON�
��*��,��c�Z�q�R�RCl�9Ye� 
k�R�˚�k)���ʕ��=��x��.e4���+��w���)I��PX�5x>#]rOsUi���[�4�e��R�M�$?������ܐ?��_r�i4�T2I�&H����G/��+_���2�jP�ϙ3�4�`��\��?\�nb�IBP1�W�Y�\Ѥ��@,���˰�9Z1�����%��_4f�e��w��t	 o5������_�o���$���� �\?�'��t!iχ'U����XuF "�Bۯ�5�7\���;��{�k��Z	�D�ULT�q�0g�y�i�:k������44:�o_e%�J �&�ON����q��j��v��n��]Z����N� /i�'w����@(OO�_k�@f�l����6, �x�ph���"�E;�o��kB#[g�>߲��  ߑ�c���s.����Ն��Q>*�DB:є7����@�;�W��O=������������r��u�~�<�z�'&��31�Yi#��7_S/�C��,d�"��.�|!{���zŏ���?�F���a����J o��^�`��!ٳg�?~���l2!��c��"��$SI���ٯ���O~)��9ٸe�|�G?�J�-'�^ ; ��MN��Îx��W�ߕ�Ǻ�)o���X�z0t{%x*w�q�t�NKJ��Tr9��Qe�ƗL(��_�ʸ;��1V�'����=^�Ȗx�3�!���{�#���瓏Yz�w�lߺM��wdúu2�bF�OO��+��'���o�<P�f6�d���7��`��f鷿alL�h8�U�!~��\�qO&�MI�� ���=�e�|�ݷe��r��&n���ׯ����y��p�ܻ��#�w��y���%)�;���`2#�PD�MN7��U]�2��� ��:�6x���D׵�dB�X#�8<	 XZU�b��
K��ƹf�����҃DB��g��J�*�L�ib(�X��$U�j��6t�R��^uiI�_LI ϙ*v]$M��;_n�?�<�' $N��FG�Gp��j����`�G&�+=ٌ�疤�C8Ǥ0	&RR�]_,��Ç�	+թgi7%�끔�x�1�y �X`�G@ză�I�%֓u >��W xO͆}����i\A��V�1)���&	m��������.�f_<�b.'�d��%L &3�<0��?�k��'��Κ0:?w熡:Xzk�#�5���\��+�G	��\3�.��E��3`A0ͱ��5�<�Ut�g��`&�s�lU8I��㬍�ٳ��w�M��m���	��w�ǰ�`�j���nE�Y�����/�������1�>�|�L�z���8W!�==s��S6�����߳`����i#��I��z�hK���^�#���[w�H~�(�J���8z`��R�UI���6�ɦk�����#�X�0�Iw(���f�&�RQ��KR��9��g�ُ���G��ͫ��~����K%b���$\1�\����֭��k�ʵ�Wd�������=�9�5EO"*��&a�܌J���˛oYmw�ڒ\���U���I�%�����\&{�� �����>���ɱ�2^2lg������'��ԓĘ˓�L�ۤM�x�v@]KHc�M:ƺ�v@��O#���TK)PǞ���:?��Iw�I_�nK�V$���7��*�vm����Hh �?>}�OJ���V Tn�{�!�"2����Ny�1����g�I�I�4���J݄����ެ�*��p9��š��<c�:F0��,y�CvpX�� TJR��%Ш����<G�uEU �Ch��%��pBm�\l�{��C�%h��{2<��w�8&}��>��#�r�vϣ���c6�ё�i]GwxA���k]p��Rn(��]v����X�e�/H�7�C?�G��=c?x���z��*Y�k������*׉����`1�Ȏ�� 6�s"���g�������?�r�E ��=ibt%i0�B��3u�A��{_������|��~��~r� �x1� ����XCek�U��xVp<�n�PUJμ��%�dQ>�x�0�&"�LJ�}�uy�cR,��\��c?��Od��n��3&�X_���s�p�6�b%a��G�O���� �f�I�I%tR�5���r��]���	����`4�����u˦M���+;wȥ���׿�5K����u�6�Z]|&����!�r�=sN���P�K,�+�x�DRiMTb8| ���u��\"�fw�����%Q�� ?��ƀH�,CBV��8Pc�؈��%��`�"�<+��3,�r���co@:-������'��>���fG�<��\���� ��V��N@���|Ɣۨ�l��V /�-�b�������U�|�~�u�~�`r࿿ztX���$�J���3yx�T`��ɴ�uA�	�T*%���H8��㒫V��H�V��ϧ�;�p�ׂI���E���3VQ�� �)��tV����2@�򗟜���.�Z�U[E�pi���
ż��R�e|L6�]'��Q�Z�d"�tըT�l���D��<���4Q ��l������-��j}��&T-ҦhJ�N�#���\ə���#?(o s�T2�<@�w�;�����k ��AH'p�~�pG�kй+i��Nl V����=���M�h���i�I���8�+~����7�j��~8�;B��']p �a�>3)񹐘�#�R XA�:4���1t��G�$"YUG��F0���T�d�	�DB�Œ,��T���X���8d��t�wn`wis���v'��A�|�ѳ�5�u�a244�.�3���'r��a�y]<9z���"�tǘ\�aMp�ٴy�����;�e)� �tR�l�׏�L���w�;2�	'��#9=c�Q�1�̗���gF%+Jz�+�RP�7�I`��H��*\~�j9�у�Y�����Z�z�����ܝ4!�^u��.Y�����=dS���$���g�-Թ��N�E%�|�A80�����În��T˂����?۸m�G�@@�V|�^� |���"�J�xz�x�@e�uIP��~�$EKc�i �Ә:1ͲM�l��Ϫ4S����,��Ԇ�	Z���>�l`=�T���e�t�iJ�\�F� �z��":0�5����[ S��F�&{�O�;Z������ɛGJ$ؔ��$����{���ܹOr�y�@�Uop�=4�`������p@P��ǹ�tq7�{Y��B���3�ָb�k{}L��=�b`^�Q����7�� ����^���a+�������S�q��9���y��_�-;v��/՚r��y�q��4�Wx�ݶ�+6�u�w�0��~�Z@j�ҵѕ� NbM�`r-��h�%���ӵ#�x���l𕼒�%�z���[�% ?	F�#�E²w߄�y�0�������{�vl�LL�"p��R��ѣGY"����7��
��+�Lq��!9v오2i�R1OpחM�}���z�A����r��WR�de4�g�TBAٹc����1:$����o�����u��!�`�z�@�Z��'�|"�/_%P/��"��K�%���0�\����eQ�a"d��~R���4ۡ�4!�@��M��AX�/��~y��ò}��&"2��|��_˃��9Gy��N�t`#��t���ؽG��^ ;q��<}1�T�6ְ'8�����2$$m�G�T*��ԴĐ4��d
���"�[§qJ�. C�s1���+ǎ��TLΟ9#g�<ͩ�����M�h�j69�xp�y�J�Ȩ�:"��<�g/�B����pD*��,�x�
\t��9ݿx�߶33p<�+&��{LB��,���>&G�  �<m�K�M��]��`oZ6��$��R���m�`1s�bmx�F�h83A�&p���Fq��j�I1��j_0v���Y<4�a3,��x���U��Q��t@6�5���̂>��N`�����$��\Z� �$@��&���cZ���2��j�#��YJ���R��uRj�*a�7�j���:�Dh4��4x q2�p�s����<�~���B78��d�ɩ��)oq���y��%�������j�Y=K�L�E� >��g�:�p���+��?6�{y��e`B9��p�8+�Q�\^�K9)�/��iM�h���Gr���q��ş��Tk%I'S����cػ�C�dt|�z����{���D��Go������2��g���uF�7qM�z~w{�ٚ��G�
��w���q�^Ǐ9<���͊�Y�C���צ�g��C�H_Ʉ���ʁ�?��w=n�s�=��
h��C%�����=Q��G���&�	��r�>/J�5�� ��%A�:b�Ih��b_��i΋�(���p2��lپ��@ �:�����/�r��_,VZ����
�!��Hqj�aw����"[#��t�fN�/{C��,�q�i9�@�6�x8m�� ֺ�f=lA��2(66 �m�JQ��� ^��A��s�6��xR�h�C`�\�Ւ�#��������+�~l�L���1��y��  T�1�.-.����ܵ�R,�R)q�v�;�Ԏ6�{A��Ň�/c�-�Y!/�A��1�3)��$�T��}xh��%�v��5k����Z	�0u�%�vG.\�*�/}#/f�d�}�����o�{$�`L0��?s�)�s�6��G�\������bk
u�ao���G�:� ��b�K�����(�u�;l��5힙��A���2�@s��6��߿I}����сd��U�k��0��.ţ#C�>ߺqSn߾̈́�wޑ|�� x��@ p�òn���,܂�o�LOR�(�>��2��B^�>�XZ�a�2��n��{&(��ͦ���ɓ�%��Sz���p��W03��ɗW�]g����da�Bw'8��{z芓��*ك� �ې��ʞ��Z�QW(8(#R�`� �_u2�|� K��TMO{�r^֮�~�;2�y�$#���E�fi������\`�����H,"�|��Ɖ=�eh�Z�(���|$wOJ�=�:���m@���<5��g��$-}E|��U45�
�[&c0�"�f�t���Ss H*�Ŝ����#y������<-�OJ6��t��	���N	ptAO
zPv>*��z8"W�ܗ�>�Bf����_��$7='Q4w�� ��Ɏox������� ���1�]-(0���� �ސF�� &�����qr/�� >ј��D�V� �L�a��_4h��	ʭ���YAa�8I_��%�+���Գ�����&�nO��k��F݆Nr$�@�s�;LO� $ D�
�jؒ*� (�|̻6������}�gc�����������)��;���p?�g�5�
��]7�?��&�<��U4d�LҜO8���nG�Y4�B��P�@C� �N��4��|��35W�S�Tn��T�lXY���SZ�0IVL8�"����tPm�wr j��w?@a��g<z�KyV�P��>Ger��}9z�ܽwS~��_q0_*��L��� �0.�fS�~�cᓧ�������w�ϑ�)F�j?0N&՘��i��U�q]"ɮ��*���7��]|���x�i���^ǰ�#p�J��4�zNlm�]'&qjř*}�z�����i������:���#�yڛ�����꼞1<�m��
�=�|M�s�*U޵���sk�^P	����J�7���H$z�'���6���i �Ɖ��z���WZ��WZz�BB�F���қ�[H�X�0��VJ�š�&i�� ��	��$��4� ��#�E ��K��:�H�_�Gͅ��'�&-�C ߁�� |�ZR _kH�MgE di��h�^k	�oz��'t�:6(J��������8*�p��(��5��
K�*�t�	�& $ Ex�F�&��%�P+s�zm�'c�<l!ٽ3��ϰW~ς���������{�k$2�HK*�����l6+�}�:>��e����^jo��5�H��Ǐ�ʍ��<�֛���@
Ն�:{�|'W���,uo>�ŵ�^{��6}�ˈ��W���n2��4hmc�s��G�&�a���L�J<��8��3��c���w�Z
ų�< �|��_��S��z%��g�Ƙ�<28${����}vj����^`�Fdp`Xʕ"�֡�����᜙�&H�S��dn1'�r��]��#C�y�5��Q�T���? �~ ��,sK�(� v��5���Jn�DM~ %�����عKv��'#�Fu� ���{�x��C3�!^�
Ys�Ssr�������s<ԡ�4j�nd@>|�-ٶn�ϯ��Jffd���lK�z����1"��Y�0]�&g�d��zY�Q�K��_��<x:�!oX���H�=/�2I8�����H"�D	6rK�S�F=�3��K �bz��])zA�� ���?���@�m���ܺv��۷n�t*��QE\/qz%�T�bA>?u�����?�P2-�<��|vR�
O���	r�^)�'����Y̹e��,����fG��ݙ�{��V��sM`ԒSY�jv@b R��B��zMj%4�?������0��V��09�	`�����t�6[á�y��β�&}��|�wH�(I1��/�����?��%jN+���L���͓֘��wp����`��N�gu[�u�����U?�XLGN���V�����V�$ ���\��]�ﮦ�,՞U%�\WZ��lSm?�sX+v��4햔�o(��]��� <�i��;�>��6�^�׶X(2Ơ��MԨ�#�����.4��Q�@�������qM�2�MVu �"k��*�"�_!��U@LZm�_�T���O^?z������ϯcb5=�.`�dU$�����߰� ����%����έ��{�9���}�Zi!���[��i���|E��2o��0Sp��J��c���hkB����@��*l��{����T]�d�}VoFR���Ҧn35�_^
�$o�]z�
�i�o�14�'�uO�C5��P]��>���x_'A mֳ��ᙀ�^Jg����'>�j�x%���~sj�g_]���r���F'Tm�T�M���Ҫ�H� ��u�P�|���`Ti����� ۔��q�p(}a�ҳ��e��L�톌�5X�=r�b��Q�Oj��Z&�5X��@��    IDAT�q�5;!�W�|`�0��a,�V[��5�$�nQB�
�q��VB(=������C%R�v�"��F���o�P_F�ܸ.�st0A@�G)�RVI�dR.Sfb���r�X�R9�߉GUW��l�A��pˤK�\�?LV4Yr�q�h������v�%�	���seQcO�!���o�6�q�?0�Nd��pA����9d$��j�E0�ddd͘lݹ[����9��ܾs_�����M��g�*SX�ʃ�E �<X�U��M2 .(�qG�7S�i�Xm����fM~h��y��a`�ٽdAw�u�[9��7���d��������{�懎��~(��m���p*���P���jfM8`�ՠ�i��qY=�F�}6g����+ynnF߿��e�ƍr`�^����Հ\�vS�>�'S3���H�������~!��~%�T����0�{���
K^e����g�����;H�0�֖�wM����I��0A`$������l��ׄ��9��F�g��%����|v�Ky��	$#��l� +@Կ���21�N:�%yp�<yx���œjF0Q(�@�ޝ���{OK2�'�v�B�#���\��H*2&�a��r�&��<{�#�zSғ�K����,�M�~0�`�}�هw�D0h�D�5ɵ��(I�V�5��_�?�UC2��ܿu[֌S�yN�V�w�ʤ{%��˯��_K8���Gߔ����_�9'�"1)�d21��� �]��7 ,�״��� u�H�"�	���C��2�8��W<�ǹd(�[�S	L�1TJ[���Cm��t��b�v�M�9�p,�>
��XS��Gti��}��/8�z9�+fn��^B��x���8�c>m�hUI��w���_s/4���J�%l֝�>\-�����a>
�(��j��M�[�k�F�U�i�-Y\������D}�XQ� ��f�iC�d�R���G�j�@o?���̬VO]����I��}���A�(�5�����Fm7� N�YM� Wa\H���\n��GGз�]����d�風��١ái��Æ���`�2�ްI%��t�``L�_\��RN-kq_�49n8,�J�dʏ~�r��a^�����Z����T�B�!���$c1N�Z�'�ͦ������q���P%�.�}�*�nP�o�w�
�wƺd��}�	�6ǽ��B��Y<d�a|�����X�)��M�h����ML���Yx���{�˂P�4��D����G�9{��L�<�۴�Egc�uO9<k�N+q!$�糽�Ն�'�ΓX����b�ɋW�t��|�ؔ0lݠy��U�I�<�ge�;F5GB�m�a�((�D�����!�P�^�E��d0��mi�2������m����+!�<�!��.-H2���< Be�0�����-��R^BtU@��ͬ�⬣��hX"�c�'����QSǢ��`�ay���etd��6t��a�V�Nw�#�����4�:t�d�23=)��y���^���!��j���	��ι X��;P�h.r�gyt��֯���� ��L��U��S�,Orp���[%��/��|Z�FrV��$,<}��P`�#Q�@�x\={&�\�.Sӳ@�|�����dJT��C�-=�	�]c	�B��j"��_�i�l�RKi�D'6Jc��.�=�F�l��[�ַٽ�c��L�^|���J O���W��ZׁyId� ת�&�ٮa��f���}�{�dY1�J��Խ���Y�v2Û�>���������j7=fg���g�;�K��D�~�ȅP$�$I� � �%W���=�=���wy﫲һ�!�sߍ�2�zvf%P�YU��޻��s�=�t���6P��O059�_{�y��)ِ�ZkE|z�^}�gr:z�0����
P���/����Q��8�`&4�~�ps�2.�t/?iM�3�k9gh�j�l/z�G�����9x�q3��yM�����H2���{05��D?�]��rU��.����~�86=���2���wo��́Y���W�G���r6	fs,���ŋHfz1s�$Z�^�������5�FLH/��K/7Ta�"$�Φ��h
��S����50��S����jUN��a���1I{V�jE4�L���O��a׎Qܼv7/]¾�=8�����Fa�j�����aaq���՝z�y��ă����GXX.�\k`�PR#�����~t�zc7�b�P� ��&_qYZS��v ҚQ��A��*
���T7��{ѓM�Y� �"ȫ��!�ri�9dXB�������2�؉'�o�L�,�\=i!	�!Le@��(�00��wɾ�aĉ'm��"9�Q>�DTnAtb��&���a�l&�#�,gS\��}�3�H�I�F�FE��%
�g��&����595TX_���-?;L�nĀ��M�J��4��b5�|�}�Zr�ƭ_�S�waߝ��DgT=�,L��z�8;��Kɫ% IU�8��I����MYA��g�
�c �</:�F@$�]^K4U��u��փ����R�b��6��$�crN�O��7�Z�<�&_���ƁÇp��9�����-O�\똕�F�XS��!H���)��<��~攘}���U8(��f�{�J��l�).oifv�i;p=9A^md��	_/�=׃��s��d.C�m��m��k��?gT	l�"LR�ȼ����;�5��%����^���mDۮ8)���u{��㾱�cc܎$���MO����{���` b���o/����w>�'��ol�[�*a��F���a���n��xԤ1�q]K��n��#KfV�����;�*bq���R���姄 �&<��6�0�tw\�JL��b�YIeՂ�B�$��m���M�˦��8���ZXCum�ͦPf�B{��G���oT��3�e��c�xPM���@oO'����l�ȈR�[.T:7�SK͜� � ��26֗���������Z)H|�s�+��燚/`~�[@p�����و�u��.Ͼ��-���qpM���$� N ?�k����p�\�J�tYpw-xi�8�$������U|r��ݟՐ:�"f��؜f�_,������`Gm�6�,��P�q�`.]��F����7� g�8C�H&t< ��8���_�ɢ��_�0 ���fZI>H��&�eu�Y��T:�Ě��V�P9�+ס6�.,�r=޾}��^A2���#�1=���>n^��C�f���amig>� K�=�'{R�����8{�&�~�;���~��	�.�Sc�R2�	�n�Q������5�J��X�֦IV��?!k�!S@���رL �`�l _����]صw/N<yc�x���酋f!V����N������pdz�����]ܾqO�~�v�Ǿ�z�Ixɮҹ4W����3�S��+ۏ���H �ޝF+�BmS�ѪN�œ� k"�JHO)P��������%[���];+��\� ?��A�j��zm#����}S�ø|�,�߾��O>��3��덒t����e{z1��������;ؽ�0�&�Q����o���
6�U�jl0�DZ��?���6�3 �'����x��S���c�$A[M�7u��ݑK%0ԛA.C:��7d`�\rVCK֒���� J�TZs�*b��+�j�3xX{9�,'�6/��\���s���$$��{v�p&������j^e��U� c�]g�� �q�I�a|^x&�����а�1Nt��%ݏ���w%�4ـ9��b�}:��E��ʬ �I����,�;��\S�0�+Q`e)HbH��KCM�IK�����12>���7��c��f�ު�������H�3��z�8����P�$2Ȣ3��*�s�M F��W9\Љ"� ���U��'��cF�DYx??�C�_V���8/�@�-Kb�|T
0�L&���|K1����{�g�$&f�I���a��Jy]M�<���8���019���8�/<����f$$��%�VA��S�w��OI����z;`��gl�&-}��r�1�!��}+.i��ۚ$]6���g�·IuD�o�M�c��{�������?'R좵�0��z� 	��ؾ��y%�	U=���W���D���ῷk���ۯ����5�?zs���>��+��o���
Pf�ejK��Q*�<�rs��ÅH�)���b���Ə-v���Q��� vNM��znqA�97?7t�F��< �#`5��v����|qqAA�͒C#���2juB�L�TE�&=f2�O0���@u}�FC��]���� �;�@*�C<��!M�-�(�*-˱u�a�.��S
J��Y�Y��d0��j��~�"ƈL<y��2��c/��d��� ~w�_��D :�����������&��&�+�ԕ�'�/���\2�E�;)�Β5�TVs�����v��q��#�Xd��)Y~�N���{���cP���#F&�t��hӅ�|guŃ�S�~,eI��2x8�C3���dO��6Z?�_�F��|�1<l� �eU��n�������Q�-g�������Ռ�B@l6��A>� �ѯ�_s�}�8��I|������x�7q��]w�tdϞ�,FV��������'�埼���9=����Vx���;���������ܾy���Sܽsi hLY_yNK�j��t�J:����<v�٩��LǆrE֒��Y2٣�.:V~d�3�]�cѥ�q~y��>{�4�''���6S��"JhʫK8<���ͯ���]�,���o��k8��i��=-}=	<1Jt����G#�����}����|��ҽ�Jd�7��رB���m��`r��8�j�֖"E�L �\Qb�"�U�h^5�?ȅ�O��Z� ~lx���!���ֵ+(�����GR�<}��٘�Q�v��C��G??<>�]{ �4�ß���K�ң,����5�~�陔�1md��Ѯ�9u�"y�=V�����M`��U����׈�9�0�6��ǾlcC}�Sa5�I������M��RO��g���A�<o���Ȇ���$;lnd�u�3Y�I��/`h�K�WD�������Y���t�qS�('���(�� ��&�;�yV�dc�\���g�S����a��/UK��Y04�'����O6+��5B�]��>�H���U#hfU��j�{9n�9V�l�&��kj�A�j����jE=n�{�0�bL��)���&���rZ��d�~��qؑUR�$� ��h�9$)��c�!��f�R�&6货��U��|ó�R"�?R+�	8\O�C��K%k	9芉W��������dZ�L��lH��0�sY=~D��ڵ��L;�&%�YZ����/]��WWШ�	�y�{2�3O�³�>-��x�Q �>K"�4������[0F�Ms`-w�m�,��	�<�$2	.�w�m �%K���ygz�{�.?����s�]�~��|V���=����c �M:jh��f"�|}xt��ܹ��'�2��W?��ޗ�����ך��Qi$���O�����جV���k�6=����d'']O�)o�E�+2X�DN=~_�ҳ�ǧ�������{�b��LP*׵٩i� �O��j�jS�PW��ʲ>��vMM�;������!�d���l���Co�m'�/����Z��ҔW�K7A /ge�TZ嵮d�eձ��� �S)������ �fS2�\�bxȵ��Y�q�ZkHG�lJY�X�S2,d�S��#���W�
�� �h7Z0�	���#������?G���>g�����lX����w��J�L�]g��fd���ܩ�*�d�\^Zw2��A=����'8M'��c�_kk 	_�����]�2���w���z�R�J�A�V��P�k��R�l��D��1E�Di[�<�/��xI�p��a��6��p��\��%����M��8u�q|緾�7�㧯��5j�	�)?I�Z����ӧpt�~ܽy�|������q��Q%�м��+8q����ϝÇ��*��Ș�F�ł�
�"ʥM�˴�,cueA{��)��@3{�5�deu��]��TO��MT�����~5E��8�F��//�����ڿǟx#S��^���� (�Xő=��_�MO��Z��3b��=;yL �=�JQ�u�R;����ҪlOٰ�c� �x������@�G �xSw�b�le�jd����9$Y�#Q�2�`�Wg��,��6�� UQ��@~bt_���7�47+����kh��J��j�kH=������/U�؉щ)�S���?��J�l�ɬ��gF:�}���X����%�Ey��b)$zrAϪ�r��v�h��l���6x��+����T�Mwc��R�b�udR�<u����nY��iA>����GC�?�fOo�L^	�f#*[�gu6	�����do�%x��DM�ab0`���B��A$�# �?�����'�[�d"��i���D�i���N�� �	1�ɔ��sHK�++�A�B6��_�v�wIeH�"��42&[X��]��N҆���5T�|svE<���>)l
����3%F|��m������e}(|���Y���#1C@����<7$�����ښ�l�Nkm�P(�1�����֐H�����IB��āf��YP�����ܯM�
�w��X]���DWK�S�?�W�8|,�BO�I�����С���{�f<�_^X���CT��E��Hg���=���c'%e�'j�e6�����&
%��g���=�Xd 7
�� ^R��٤^�N�-�u�v
�@�:�]�wҲ[�M�w]y{�|G��ݾy{��@ޥAVH�q���n{r����II|�	>)�b�d:���Ď�j|׾s�{��>}���~�����O7��(7�&�H�hcyU�Gd���264�}33j�[]]�իWq��=�T>+W�27fw���ܨt=��r.r��#��W�WɈ�G�|�m��ps�P��"���TrK�9eB�)_���4��y�
똽���E���*�߾�r/5n>���.��������z�T��VY���)�Nbivy ���6���Cޝ��C֐l�jkMsIـ����5X���mֆ.&)R c d5�4Bh��������CA���ȫ��eu�3�ntX��}�y��/~N^go�h/����7f����s��2�Ϥf� �`�PӤl.	�m�6'�*�6˿�33fV#�1��2��.�29kx�&��Y�V�mjh�������rk$5��M��B����
�:�Mg�{[�ٙ�g%����יv��&Vm�m��6� Pۇ7R�{�w-n{ ����aR2��"^�
�]@>��ɓ�4������O^���+��]Q����5�'O�Ф�&�l⫷�Jg����_ū���cǎ�o��o���Oq��u�8z��|R��r�.�Ǎ��4�&KB��ԫ%�Ҝ@6��l&��|V,<����NI �qp&�����;(�:�=gXSu�-ŔW^{��2��z
��v�O>�n�T����:r_�4&�-�ƕ��W9t� �wL���zfE� ��kqqi|�)j�n��ُޑI���7p��"�A4������V�e`�$��$^q�$�&�8�T�l�Z���m���4R�AK�je�c���׾���"�k�X9x@C��L7���p�r�u{��m|��?@��D���.:x�p��5���Hg)���f��9����%*�c*�m�4�.9���g+�QU\k�e �,ڄF-�&�.{Z��0~oVJ�$����Rd��L��J2�1d)�I�u�}MxI5Z@�@?����f,c���{��H3��US�JH~W\�=e ���m�
�Pt�� Uа;�ɵ�S�LԻ"��%�6�*lt#qRD��p�څfB����P�c�ksoPS��� �rI>�7��9��K~=���`��Ym5�.	�8�#�Gy-V7i�9F �8��?��.�q�x��CB�l    IDAT��w�а�*��guI��"!a�W�bY�7�gƉJ��M,.�`qu�k%<x8�5K	���l͡�\��2S�=R�������[p3� vZ��t�G���
�	3ٌ��wtl� ��ځr�U�U�,/j�����޾�۷oj@Yc�b=x�8v��)�>}�	�����&V�C�txcu�a���
�G���?G�����%�׫��-G#$�vɈ��<��K��v��m����H��	ޭ�x+���ul}�=���m=���z�S*qQ/��~���d���%�����_�윹�+���Ww�����\�~��]w<m�Zn����P ���ظ6�(�޽�b��T6#`Vn���w��gr�c�� ����DC����p��uܸ~�RMl��L��J ��af���I�1><$��kƆ��aM ���..�Tm�q��	zζ�p���uLO�ߛz��VL6�Z�c���b �Zj��қ6���<,���LlL�b���b����2��r���u'��A�ИJ��!�Ƈ�~Xm�&;��ˇ%h3�u��P�c�%�WnӱD�(xm�P�
	��|3�:�tЙS��d(5��i��	�4�Øq9&'�n+�rc�_A�,Nڋ�UZU�R�)�dQ��Vf�Z���+,#G&�Z[��g.H��Ծ~V��i��Fow�R�[��-g?�o��9<�-��&����+�;��ބG�P�P⥎<C�8XzKF��� :�>]�zr	<�O����x��w�B{�tV���#l�*bo���Y�	����l�R	/��c���8q�8������75���������P.�G�駟���[Ht��	O�T��T�R��[�b6�:Y��R��JZ}34B&�H�!��k��7�=�v��K+(�X]/�G?y	��2�?�'v��O�����G��x��!|�KO�?х��p�����ߏ��Q� �)�\$	������*�ڃ����^��z��F����%a��P��H��$4aS����/>?��=a�3� 9��19�_��s�L&GGp��A��&����F�a�Ք���_B��x��z�K����d�Hf4�S��X�_��枡*�*I>�&��� x�|��+R#�S+��U5�6�%d�1���"��!��wN(&�$4�JJ�ĕS,	�)��%�4)hУ�w�Ij��Abp�p�'�.����D�a;��������{DL�~��a�֔���  HBb!$ֈ�q�l
�Ӓ����a^ϵh�����
�C�����h����|�%���2ɬ�n1���$��J�����K�����e����'K"�����a667ے#��柁g��d*��F<�]�bE����q��9ܟ������%JA+j*��ǜ����fZ��aJ���f�/�,+9��-9�p��7�ݧ�~Rཧ'�&(��,���M�s�._��F���n��J��+��=u{��FCø�1�<��a�G# �}f��[��4:@�R=jw��g��u`�#N4�.x��e�?)���6jg�x��ɒd�H��>�~�(�-��U�����J���� ���D-ѣ��݉6��$6<�j�Ļc�J*�������fl��������^�}���t_����ht|��R�B9���o
3^��4�٤�';�!	e�h�P+/#��BOO��&T����ǃ�e�H��t�a�'� jת���.���kK��}p��
ƻ�����:��֕5��p�N&�=����i��
ժ�+�x��2~F�0,���7�I���(g��>�A�gTܖP�����X@ɚի�ɒ��K�=�ɐ�灱a�f�|�beZy���s����:��,��J�%�M���C+xmx�$�2��'?�J��&"x�`�>e�d�����A�c�l��`5:f��c�����n�����O?��s�Z��{����AG�
\!�p���5������͸.`�Fg���D+4���J����'/��u|�P8"�������
xM4�	dhN
��̜�A���x�|�O?}
_��Wp�����k�;� �|��di���D��!�B6��\1�����u��a�����+/�������G���e,�?ĵK�p��~1�Ã����p��@<���C�8r��z�b����<$LG�k)��l"%�j��t���!4�RhƳ(V�X\Y��f��~��ll�s��}������p���;�|�k�n[bS�b}~O�8�����ob��<�s]L�ѣG�74�f/	�XE��5S����Opgv��3�ۉ����P��;Ӈ�$��'�I�m�EcE���ue�>R]�BC+IU�XQ����{朤�k�� {h���sO�Bi}YM�GА�.��4Zu6�ט1E ���be�(�wz�ߛ]V54��E,�B<�Q5�<�B�cЮj��x�0�;켳�I����3�
�P�Ě�!㮑#b��R�� |�z��J�M�1ܗG&C&�@O#��tqn	�o7�rYU~G��$��NY�'-9h���n;�ˇ�c�LBglnes���ߙd��s;�9���[��ț��Y��A>������X���;c)+{��o,����D\px���*��$���t#acS�MWe��w�'"���+1Q�!Q�l���&z��КQ9����W�|����y�c=�1��"�c2�b��4� �71C�ҩ�X�D�,")3s�a��<�%l"y��d|�K�#:�$��J��~9����^��?�w���F��fwe^�	�4�!R�������L�����E���4|� >��t�"!Ş��O��c����ڪL9�\O��j��h����,/���k��7T�O��TD�D����)ɪ����G�#j��d�s |�(����f��|� ���Г�D��e�M*$��-$�.uW#�����9�v�(�MG��	�����M��$)μ?B�U >�����H��h�ф� _Lg2�a�Ν����̝�����ǵR�[-�3G��c'NJKX)l��a��R�,ɠ��ZU�I�|�Xؔͪ�#�N�����f�D�҆�ᜲ���R��b�޲	�+�%G����]ئo�����N��\F���bIjݺ�V(h|z7�.h��h�G�:�]� ��f�&�ѧ;��28�P�̰�!9+�"���k�&���������_,5�ʰ5��'��F��p������qT��Ș^�=w�_�5�n�N��'�y	�Y -dפ�;���v��`7��� ��Ĥ�J&E���ky]?Mj��%	��6h�8x����(�.2f�d
��;��~�:�����ò�,���0��ј��.ϓʠ��b�4gi���e��yb�f��%ʦ���v�s�!|����ޒ�NĊ2�hu�gH�s;o�)z	0���LC�x���#�:��38|h����@�T��}��sshu%���>�i+�pg`jb�''���-ܹv��u;zG���tԗ^�)>��#B_����ݿ���㘞����]bB�ݿ�k׮�y������*�jV��8w���Mv���v5b��S'��1�B�Z�\V�
jt�ב��1�c'6
%�o�p��~���P���ɧ���Шxx��f�������o��%���n^9���Q�8q��&)�暞��]���n/��:�>\�Ι�H���/���e���UM;v�S��
��gU��e��������lfM�1M�6�n��:�\�{ɉ[k��F��Rq����3O����F��}�����O���G.-$C��ł��I\�v?y�%,.�#���Z����f�]Og����zP(UTȲ��eAܛ[[T�`Q�����sڮ����3ȇ	�L3�U�-��\hX!�_�]��Bӓ��qs���#t�f��d5��\��y���tNe`^��s"",�%�f�GJ~�5�8V�����>HGx~q�-%�����'��}�9���P�R���e�H3��ͩ�U�XdoVl���D�~PRa;^R67l ���ʛL#oq�c{�6����͊{�(��X�3�V\k��	��14i���h��Kr�+���P�� ��1�C�u6b�	%�jN	�m:��-b�n�\�
F �\�L��h��H��h��v��ܬS��ą���TFY,�Q�o�����p��e�-�"��U���<�ei���h�� fh)Y&������4��<ĺ�.� �3���q ӗ��b�n�?�E�T��� fv��5|8{ׯ_���)?�ÇP�D2N?M�ľ}��ĉ�n�ʃ¹���9�m���lR���U.��V2���}�m3�py���߹�B��뚊}o�6V�l�^<n�-��>6�ͽɟo�=%)HLhR�P���]߷ѳ����#,�]B㕶G��Ϙ�h?D*����5��{�+T�8gޣ�Q2C���z&��7c#��pxj�������<�����j����fh4:���/������
�^�33Ц���>"���ԡR|�toк �����p���o/l�XE�X�����3̒�m��'���DR�Q%d�#,
H�ްL��iZ���j#H�C@�r"*��+�Q����t��LzcVT����*4�@!�<Kx�]9��M��orq�2���Lo`�մ�C% x2�V-ʹ�1��B������"m�F���IL^��`�d�l�& �`=F`#�����.�\1RJ`�HhTs�a�S`�|�������M����k>|X=7n�Ƌ/�w�=DC_B��,>���ZoA���2��)ψ�0 MW����Gv�-�d��2��4������/ ���� >ڣ��
���d��k5��nHc���#�cX+l�,�GFt=?��CܽyGē'��nu������#P�`�^{�u\�v�?q��گ���{G}2�n�����C��9�t��3{�18�#7NA]��TKnԨ��e�.�HZ6���K���cau�/_�����ۏ�{fdK�hva~q?|�(T[8~�i����'g4�d�Fa���ݯ�)`��ܾv�cC8�fO6�Ǩ�� ;J�l�%���?��f�16=�����$��х��W���ғ� �������*Jk����`cg��Ņ��$����k���F���~	��:*�uqz��	��IB��d�bU�y��Naie?y�e��x	=}C��M _m �\?ɜ <��	������.Y���GTW�O"��EW.�bg��E����}�C)��w��������@>�\�ң� �����%p�����a>g ~��e��b;��N�}�q��~жe3d4�CK��`BQ`�-��a`�$-�����>��IO�Dvx��۱�����Ҩ�s�V�<�U��Mw�qެ�u��|ϚT�4��I�y�0� sw�����U��Y���V��6_lz����� �E����2�%�v�:��O�4�{�[~��ܪh�s׭0�x6�XyhrX�	��w�����鹋X-�4�Lßx�S����f\k��r}i�KsȰ��NGzߛJ����ż�ً���ҹ3�<r�${���irv7n����g�4?'[��&$��3�S�'{c����������c-kJvL%�~ �>{"ɀ���^)�
���V7��p��E��pA���w&3L<(�d_��e2�t*%L�Ǩ��I���sO4�"%	S�� B1nX�CV��.L6X�ے8�D�Xd��v`������~��>���A����A�aB�_o_۾gE�}p��˙l�_��Gcc{�~e ��~���?{�X/V~+��f9]���#��x�����F�6\j����`	�̚1+���.�2}1{"ޅT�ن�f�	��?�����t�Ųɝ�����y�{��HĺP/U42�Ʉ;���t�,�J���0s��:󧵁 t�1Ь!�gb���F��K�4�c�7QHnB�  xY��16A���I�55g7��Zi��c�XδɆ���wpg��l#�yѽ{��3�A�C�l}j(P`�|��5��W �� �ode<~	��}!L��7���m�	� �rQ�b��z�Iwl��Pa	�������y<��x0��7��w��*�'!�"�7	�1Cm�����1w�a��� K�պ���������pP�Ft����䲚��5�����!�;�.4Ѡ����b��R`�f��s�„	c��/j���ⱓO������S�u��p�.^��{7o�?��Ǐ�о=K��1���������
���8|� ��o~s��w<�HHz74�/л8?'��J��ݻ��fZ~��-2Iu,�=@�RPsb�^E&��ôђ����19�lԛ��<w�"�QB7<" ?<6���!l���/b�����O#78.� ^v��*���;���/"�]���Wp��UYl�YSb�i6�Ly��81���A\�v���܅��)����+%��ъg���-�P��0����`4(8^}�zpx�u�h��H:��c{śG���]��W�����-/�_����4�b���u耓f}|g.\Do�0�
%\�~_�*s=�H�rH�s�*#��?��Bc{��Dx9zؤs'K"A��&�Jh$���m#=��.��<�M�6+��
Hǻ0:ԏ�t]��d^;��%���fbd��&02�/�Q�ww�WoT�N��<��l����Ki|z�qá�l)EdU���s�߼f^� c�&l��ܨD�A,ߖ��?/c�{��n�V�7���J�����:��M&��é��}j��z�sw|��o�]a�J�x�EKO��0֫Ӽ�����s�H����� ���v �:;��Ke#KI�Mj�F�@ިa�$�v���g��b��%�ń�X��q�VÍ����Wob��PUl������a�{�4�4�b�!���d��I�o��v��<��3��7hY+c?'cON���;jbՈJb��+��[o�Ν[��I�$�ٷ{��۫Am##C���z�������f���������W_�B?���x�`�u��Q\s�7o����s����9W��0�D��DҤ�.���XV������Snw��9��TF��(��D���n�iG��+Q��%���a�S�_��E����*9��b2�cGs/�ףW(Ce��U��L.�/�G�����[�ȯ������w������T�/���f����;�0� ���_�$K8�f4�J���4�|j�%��O`�����lXK&���{-V��3�o���:#�wd�Yf�M������,��t(�-5���E"����AU5�$�i�[� K�Ը(o�:�Y������i�1��3؂�N�A7�&{��E%.���`���@����S9E�l��fW2��5��Cp��&����Z�`�b�H_~>OLz4��JK�����mkT��!{��Z �v(�֑K���k�Rd�rh	7�X.��Y
��������O=22��{�O�������Yܹ?o�$BɌiI�����@���Pz�����t!{R�ir.%b�4ʪ���#�RC�g|f��6 ����@e�����_���У �	B�b~��:z���kzCcc�����ZW�]�+�����[�I&p��>B��|�gggq��M�m�J>7�o7��7w�����w��e�{r}��W��ݑ�l�Z�����3���A�4@���ŇjJds"��|�:\�"�2��W�V�70���3g��ƭ�bv'&wbz�~��� ~����Tm��S�!?<��?=�+7oim$��<0��~�K�M n\ƽ;��'vL�C�Ӵ8�p�jY��==9�}8�
W�001���(��'�`���x�]�,jM&�I%��B�|�)���&J��XYB��>���&�E}������������۳_�ڗ1w�����c"b�
�u�s��{�bc�`?.\���w�apx\�Ʌ�7�K��7, ���B��8M�D����O������hc*���<��5 �FN&ܔ��Q ^qÛX�� =~ʅu�1G�z1��JNU iّ�    IDATlh@L���Ν��t!I�HSJ���%KA6y��9'�D,����2V��-0q�>;hgܒ	B�ޖ�8c��& ���P�ױ�@ :�mꥭ��՞��̦�_�9�����ݹ�&�L����{#D�Ds�ű���]�@��籝͸<�ݥͫ!0E��>G���fTY
�ɯ�9��F ٹ�\A�jR����	�	�.\�|-��9a��&��7�U���Gx�M�% �F��<�B��f[Jc3IToge��-l,�cciYxZnr�e����~�<v��xōu�?|�T2���
�޾yw��F�hL<j^�+�.�ƍkX\Z@_�O=�v�������bhx �-���|p{��m ޯ�/��q���6���=�U�bq}��w������l���*:Hgݔ�k^x�gy��֛�srm�������68�ۿ��lU���
��l6������uv�k��!����װ	�Θٟ;��.3�uI3�g�V�2"��i�:���H��2��?�1:��{'.�� �_����k���OK����[]=Ãr�yp�&� ,@ӿ�-=%/%���&�Z�����z���Sp����_� ICb��g�b�uml3�2x��+��2�ʧr�t�a)XY����=�������1�`f#�h�a ��Zz��U��(8nO��м#�����Y��nR��o��zm�<��|�����!hf!��:����E�o�:�������>�6薬���'����A��6�?�s*����pK�t=BR�Ó	K��Ni��/J��Q���t~G������paopF�TM6�܉�&��u�JJO���6-����z-fv��*֗Q�X�`/��34�EiOCj�2*�^���z��߶y�Km��#r]��$��vPE���,�pp��m��W"q,+�g�3z�z�;8(��4,=v�!��]4�E���ۘ��.N:�WP,�m�r03���{��kW/���[8��<�J�<��ݽ-����9��cϞi��	�=5iE�[kr�`S�f����fW����ws�SW��ć$� ~l|'��?��=���J��cO�����'�~�ٲ�P,�᱃��[��2�sI,<�����P,�cjz
C��e�ի�R*n �Lax�_T���Urj$���.5ض�\�ָ��o7�O���I�z֖�����%�}��O�����X6չT\������o�&�߹�K�Ϩ��K�=�ݻ�umK���V��Ľ8>9�X*�W_{wg���p�Μ��j����$�Yt�1�^�2��" ހ|���A�Cm ߓd#i�7U�qMr�p�9�a ަ�W�E֙�墚��{Ҙ�G*������{|l���`���Xy�?6n��� �L����:�vK;���쭑S2x_��*��Ep���9���QP�!�����]f�ȬV���:�����;�=��8;��v�G1�ԝ����i�!����v܊���u`81���7��NZ�J�\ƀ��\x�sB` _�L`9u���p�.O~����	����Ǔ%6���奒��6�׽���Jrn�~�l.�z�ݒb)\�~/���_��F+vJ�d%,��`��}�6`�����6��es��ɦ�V��c8���8|� �bcu}�y왞R�Е�eذ��h�N�Dl�m���=\�rE$�O<���^��?~�Fǆ%	55��3 �yf;>�uM�M�=�}bg/���|�7�z�n��ß�zq'�owǅ-���R)V����Nߛ�I�P_d�Ds��X8I���k�;����(H�3��q��;���)V�/�*�?{R�{g\�R�/T�5��,���K��MZ��f���yrp�_�MM-o	Q��y?�g?|u�����R�w�Z_.��f���{�ѨWt�0���p1�܅���3��L�j�`MY��A��{��1��ρ-���=2�Ĳ��Y�`�UX_C�VK\ �bA8m�7Q%2l���4����t�bi-��q�>l��v��s������(8v�����'AM��n|% ���3�D6�͛�T�h��#!��QS�lQV� �v"(�wf���w�K����x���Vl�/t"ZYYQs2�Q�&�7�W��!�}##gU��~s�s����r�[��;�W!�X��v%3�H�ʠJٓ�q{'�􅨂��%�

�+�����O�<̃W
f��pњ�Q�:��Hb���};�����Փ6������z{���w��v��m�{�E�>��J搰N	P��� ���\��#](o1��.��"������&B� �YI�h���݅�������q���<zT�flz�L��(�ƽ{w��>66"F�R Ƙ��<�d�٬�X�<���c��``xL����5\�t	gΝ��F�CØ�5�=��c|��*M���WP��p��3H����>ƭ��fY*�������;_��|�+�X_�������z��U�[��(�!����R�3g��ar��ׁ�������T��� �l��"����uz��ZX_]����,]Z��lU�_��l�1�X\ơ3����Xxx����þ��32$`����ڪ�`s�LMO�.y?y��9q��x�=|��e�p�����-����_��l �!%�����3 ^R	�]s;1b�*�j�^!*�$)��K�nh	��G&Սdk�L
���8�o/�>��|FC��Y��N�M�-��HLbx~Hwܧ��q��Ӷ��%t�z� >� Xu����g%�������e��\�����c��~�{�3�{�������Ă����l�uuƄ���Z�(�o���O��?@B�CD��﬿����2L���~�(�6�St�z"L�E)q��g�u6|��Ā�ƈ�~�@��M�e��jC�A�jV�`qu/���x�CU���i�l�yM��^窚�����f<��RʡuU���G��SO���X\����C��];w`b|\���>��t�$����)+��__Y�͖\h�9u##�f�Ạ����܆��������g���XE��(�׽�f�̿�N��d��~��p��YܺuK�smmC��8����$��v�6\;��I���%1����\硷M�J���:�YmG1��I`���m��I�F^K��N#���ǔ¶���2����u�(��>mRzL��c�A| ��\>�O'������_��c�����_[��4[} B=*�Ў�0E��Ĭ��0�T�2��8�]͖s7����R
n�0��]>hg"��x�ie�^;�l���X�eJ1�Ҋ����]b&�f�4�Xvo�X��5�`��_����+/C��	+mH'ZR��� 5q)�\wڕ��^?
��3o�eI�L����p�I����=$�I�OJ����c�F�M�#�5��mّ���fZ����� �-c��	=����L�׀��2KN�74b���L��$E���,e�D;~Y����	0�b#�	��k�=q˫E���9ܛ[�W)>I׏M�g�.��l �P�ײf.�!����d�E �h��i�
�rKhT~�؏�m��l�����Q���o��a��].4Gw���w?
?��g��\߼��JUm��<]:�!��f��{4�� 0�YE6ӤKM�L&4��Z�j�Ɲ�ڵ����[7��퟿�\*��V��B�`sM�����ܼyT��7�e5s�I�SO���d&�=}���ȸ4؜K�0����E�^��O`trF�'���Ã�e���k��bx��s�g{������گ|��5�S��W���p�*�(�����֫�T`��F�r���&8޾{OS�G��`��¿��c�XG����T5i�Kh�%;dB��T:����eMj�wm"Ê��C镙m�G�"v?H��F\��TZ���S�����(Wp�㏱4�Ps�B��j�*��V������dzr���y�����/��s�Kf���R����UQ�"sM�e��Hc��I�슡A	��|��>1�$4�M >�/b���X-�^͒�*�P�Rwߪ��ߓ�̎1d�q��}�eRx��>tH>�ݭ�,4����qI 0�$#�5��ty�k���Q`/���Q���L��aГ~��4k[!Z����zg���i7g B���N�� f��ɚ��1�I�PE���� �����ݝd��:皤Q$���@�6�Z�j;5�|���;��s�����p
X��ͼ�g'T>����� ޯ��ĉ ^�cx��ϱ�P���@�;�dUY!AIQ'�K���z�C��ڛ�/��,7Ow�.c�CC6�S�� �����c�YMi֨���� ���8rx?*�޻��\��*LyO�gϞ�;�#;K8LM�V)�I*Ѹz��\N���8q�(���L�^ �[z��a�*+o~uI�\7�3�7��Vt�E����5����bsUQ8�]����յ5i�)Z_/h����:�=�;Nu'���AxN�g��6M�5�$O���7�a��Ax��d�DNc�Hc���}Lև�/[�a(ZH@��$hh�12:$g���A�1�����M��Խl.��'������G]k����� �{�]�X��d<֗�d�|m+�s(�6�Mˉ%!fX-l��/c���@���]]�ܺy��<��^��<g����o�0�Jh@�J0��!LM�¬���:h����ޛp;C5��� M���L{��U�tn��W��#��@3��}�y`��͎H�6��4wd�5Zӏ-6]onR�t�/1�=��E���zc���]�1�2	�[2�^�A��cb��p��T���Q�L�<+5w�.�0c�^�fr3i�g�T1MɴM��Ueo����'�\(����]zT���LA)AA���kc�*�AW������'�\�
���V�be�
y��Pwp O�+����7�O_��Q ^/Y��4i�����A�U������e���"�{�v�	F�d18��	'�#eH}C�����9�+��,�fT�{:(Л�	t����U*��Se���;&����aa~���Q%`j��r9|�k_�ӧ�#A�D�&:*\9Q�7U5ǳ�W���a ���ݹ;��108�R��%>1�\�}�������Ս��x��o����3_���wq�ެ>3E��5�م�=����Г�B>���{(�
�@2�A��)�%�cw��g�&6��b`l'�H����,mT�@�h�ͱLH��:�)�	&��p�W$��JQ��&V6S����w�K }�`v��˰kGɩ�1��5�����q��e9p�>����d2پ{�r==��������*������x��fd��JZHƸ������h�M>Cy���&m�ؔ�b�\�D&Vʽ҃Y��[�(���<���K��=�%�QZg"�DO&�ǎ��=�5�6��)�g�"2���)�w �o�����H���]�:1��>���O��8p�g��u7���=��e���0M����`LB*0��0�4����q�1,du�����h������]����	ܝ	7ݰ�c<�q��+�!kCHn콚�S�B��	5:����J����ʌ��<	rYl�x��6^}򜢛��&��]�	4����9���x8�"I_�-�1Vig�VF���)~y��ˋ�-�L ?�߇g�>��G	���0��)ɬqU�2~r���%��}%a�s�ݷ����F����ӧe=�s�D�XՃۑ��	S�� >ʪ�" ���>�أ\�gb:�D�I�f��:6��RRE�Q�s@��P(�R�����>������{���Cx>��ʪ@?MXE�K�D���ו�K�H���	�wW���5��o�&Yֹ��Y�z��δb���D��/Ůn����?�v��#:WI&D��6�O$�d��490����a�#�>�SB���o��fc�{S���z+�K��.��qa����S��Un~���CZ�p�`	YBpq^�@�|+�	�r�l���x̼	��%ۗ��kp���7��D��y����Vgp����ۆ�t:�Cb(��1�l��j�ԐT��*��s�A+ݠ����`_l�?; ���,�X_���L
g~�>)�"71U�,���$0j�u��N.�ʣ,>7`��br�+ٌ���8T7���㜀�JJn�	�}v��x=�� �+H��*V=�?�=������by��W���.r�G��	m���N�Z�`�7�d%���3\���jeWVQ+��,<�s���/�	3�_�~@��ց�}��m%ɭ�Θu{�h��B��}���ߟ�����H�	�O��J6P�ojH��|_?zG�Q�Rj����+s�ҦgY��LB��k&��岒�ё!����;���[o��|��T6�S.CIeԤU���,=���ս;weO+�Dӆ�driMz%?69��;w
��Ũ՚
��t�PR�F��l��7������8����[]Ë?�n�{�ɾ�j	��039��|���9ԋ��6+E5w����7��V�RuJ�(�h4�Xă�Xm`j�>�M���{��O^��F�Z�L�ZS�Z��&J%�!9�C���G�{2(�.����i�ɸU��R���[��qj+��;DQ�v�jQV�����&�^8�	�\>�Ǐ��_x���������p����B��X:�����������yd�����\�*	w,O*� O}&}�~� +��Q�#��'{�Ѡ���;S?� ����SX䲚o�P-m(i��	N4q���5��S'�w�.xs��B^��s�w.��1�=��k�o̴cն*��K��o)� p8!]����/�a�e���t�ř�6X���.g�=	��N4�{p�d�ϐ�����>�&s57��ͮ�2�s?��"S���vm�k L�ؠ��-"�q\Y�0�J�<�r"̙Y'��I��g�`��賄*7ߚ�ԜӍ�����_��^z�nޕ��G<k�ܙ���.�j��T�K󨬭h]RBg�O�.II�	=}�)�ځW��Z*��ozj���)�y���N�GFp��!��%<s��U\:�,E��W��%�<~�lJ�T����W߷�����j�-Й�����6!z;��}�uJ��$�Na�+ټIk�6_�=O�s�"�
%1�j*M%���HB����9=���"#x�g�?V)���z�L&�	6���#��h\"���QҚ�d��׉#�s̈́&����C��$	H�q�'��=�ٳc#��5'�E�M\������ߏ�����3k= �ƻ�jԿ�sr�7�Y�;�����
�����%z*��A����V��)��Cc(�,���ogĭ7����t��A-�T)�Q`n��)��qSCZ�F&�"@�20Ϯm@��c	���,�Rz`�� H0���X�v 
�L�A޻���,��|<l���x�F�x�p�9H����΃�p��p+e�{tΘI�џ|v�C��j?g��ʃ����O:�t� ;��l�����.YM�3����oq,��t�r��w5Jt�V5/�l� &vN��c�c�\�[��͹t�3�Rn���tT�f�3�
�OA$ '��g<���c��)�h�ʨ���RZGrS��0�)��� --�� ���� ��R�]hNc@�}���1u�h�aLlq:׋��1TZԚ���(�����Hl60�ρw�����R���q�fK�˿���{�Nˇ�6h,���&	b���)� �}������|�._���:Qz�*5l&}��4\��T~q2���|<�p��o�+�7����l�]�����.f,&shL���;G��/?��|���(�.�R)��w��jb-� ���1�$2�� ��}�T]����u���S����Ʈ�Gh}��F~�q���ɡ/��4�`4E֕�|H��TlnU�Rk�R"ȵnO&Mdg1�	��L���o����ܹ}�woa��8N?�8��F�Z0?�`���;�)�#���t�:�Ϳ�31�i��h	91��,��j�C� x5���)�B���|?�!��c\d��6U�"Vn"��u��DecMv�=�4zsȯ作    IDAT�b�ͧћMa��O?��w��r ��ɘM��s�p_(�u�kQ��c��O�[bp wl�<���Xh��]S:l����oN������q���2���ud��qrII_� ���ߝ�K����̿�{����ێ1��W�D�5���>s�T
d�=�����Փ�(������g���z��C ��%�RX$4���f	$29\�q/���\��b��,��$�l��b��n�l�Wݛ�X[�Gy}I4��� �<���o~뛒m-�'�n�&+w��ƙ3g����������c��6q��Y\8{3K���_�2N9�\>-a��E{:{P1|Ư����Q �ݶ��h��	$ч��G���c���:���^,HEA��R�d�����Ab	�9�������fk-a��"k5%��Z����5�3"+�_q&$]HyՋ����J�J��EC�F�O<�e��u�.�sx��g����݈���l ^ׇ���L�f��������Ȉ�]��%4����?lԫ��kr�7׽�)���s�d�H��t<��Ի�}�
@ j�3���@�VG��Z�� 4 x^p�P�2����w���$�A������+�����,\ئ��dm�H����N��z8��X9��*��?w�R�и鹣 _׆�=x��5s��(���h;��&�!�y�n�9��H)�Q4�F<I�`���YC�5�����SS�޸I� du��D*�Nv�Ǭѣ�_��6i��uw�RnH�A~db��8��x���m�0�*$:
�aІ�d8������ix�T�+(/�j<5<���]��[~y =l۲�_���׋�Ƕ�ݷK(�F�1���`���;��{�a�4� �Dn` =��ҽ��%6�������x�����$l����	���ZCC����}{gv�)�b&�)�W�;���^�������2�}�m\�pQ�8&�d/6JE����q5h8p@k���zaC�%g~NZ#�:���ӗ[1:FıR(��z�,�TjU$�8�g'���gЗ�aq�6�C�T���i>zD�T��>��Y��J	�s�r=�܃�D�\�����T@����V���V{�i�\�L�Hƀrq��:b������&���S���f35��աk�3
�GG�����5��4�������9��V�ZY	�����{}r����\ >���ϻ����ɷlY;��mG�6�w	]�ȮY?C�$h�cQ�.f"�cI���F���RI�f	Nb-���$z2	dSq����R�ó�Oa׎I�4I�|<��lzCG��ǫ(+���4EA|�G㢽� i
�s�)���7nEQ٫��<����?[����s�y;h�>��e8��\^��I)'`���(��g�%�`E�[4!�~�(Y�Qbږu*���>?W���_g��!w;�n*��T�hzY	K�� �����W^_&F��F]��i��h �BS�U��b�Ǻl��"H��?�C9tX�2hW��0��O&Y���{{���8z������ipI�$F��k_��ڏL6�>�������9X�Ԋ��lmK���kj;��G*�PaҠ7:,�Y������u����5�{�Ggyu]��|���3>ҡNz�Z�}�������e��{�3������hPo��`iKK�$�V	oܾe����M�Q�ZU�� c�����bg��v=4X��zh�>d�Gc�T���C�������{����?-D��k�y?���w������N���Kv�������h���{�捑^,x��A| PA}�{�D&Ǖ��ra:W��ݻ,�W��r�o/$�c6�dܶ�C�)��
�E"��4ޡ�D�ˈ����,Ԟfi�q���(8��Mg4\R��s2�P-�gp`@<�zP�d(z��P�x��|��}i���G:�5Զoj�~���~O ��_�&��Z�N���YyOr�{|,KJ~d"�����z�O�l��SU�]�4P��D�o��8p�,�>�|�������d⥇W��5 j�n`��$�
���T1j��'��' ߖ.�ۼ]B��{k�%$���Re�jSL|:�G�А��:ͤlT|qcM)]�*�8�d�)e�6��L���|6���>5	2�����eHw���e@�22!��W�X^XT�(�
��r0m�J��z�L�7�3y�YN����`I۴�����Z�*V>�`���FJ+8���Ϝ�@:���L�#9�?~L��bq��+eY��5xx�
�:��w�����;x�7�R��X�Dw<��f��q�.��ĩ�M��U(�PŧQ+I_-�K����b�ݭĶ'�Ӟ+����)- ��^$�`���Z����>|�7����V�瑊ua��܏�<m�l*5�F��}
�
�q��I||�<��_��.im�fOp�BKd&?����Z��`62�����"�o�z��)����DG��r�	���b���&�=c,˒3�x޿��YY�U�UY�{߮��g���bg8�b�K�� �$Jrw��S�� jA�Xؑ4����]��{�Io������UM�R�	2�{߽�D|��p��2��1+���N��/��� )˼��<�w�,�[��
Ћ`t�O4n��z\id�5(r)%
>��
�j���K�q��t(��=T��M��1��i���.�W � ����Ȼ�U}���N���;yӠ��&`����<�a֌g��\@Q����x��:���y>p�܋L|��}N_���~�������+�� (x�H5f�
 ѡ�
�
w)�S��f&9� �!Bt�d�#�Ѿ];e��͜0��e)e;99N_�4������PC�a���D�~Y��-Ͽ�O֮��v�61k�Ia��!ճ�����릳U8��)��b��Y����3T��I+C� ~j&#�C��xhPjU�����{"������F��,�[�)�cǎ5�4�-```@�o�(K�,f�^>�e����ν��ks"y355-�<�G���G��,�Bݞn�o�K��j�L��Z8 �wl�$R�,h��@��/t3��򧩎Eo���d) ���c�~4�hAkk�/��Q~����\���i41��L�w�z��� TSꅳ���	F�au�-�l�,6y�t`--4���S�dh����!t�WНo����ͨ�1�q8|��f�[c�9 �� N�V90�]p��xhj���O�ڢ�I�{Ԁנ}��*�`�6���N���fhv@3����)����o3��󳜯偺( x�^��Fd��a=xc�Ay�ͥ׈jB>�,D��DC JT �8��h�C�W�,�DJں��途�!9��3sP!�7!�eY)����VL���}g��7|�Ƽ�f��mfi��;�V��_�o�)�� ]e �視y3�~t��7�Z��N-��^�㭭��9e�L���ԄL��P�<
�}d=8,��AK�$���5���2�Vh:&�NI̓��Q�]���Q���	��Q�1�N�G�WQ�	K���D�R��F@�5#	F(�E�@,��9�5��o�eqO��ټVZ��~"C��Q�y����n�Z�Ad���"5��
�?~<(�|Y�zI�����[�L
g�C��t �X�a�ԇ\ d߳9P@J�|�TG�n�P��%�*~T��mƖ���\kӃd�T+iO�e���y;��Ě^�f�l޴Ab����T���|쏩�9{�B1y�hP�:|\�&2��I=C� ��}��:jJ�fT��%T���i����HH=�AN����i+��u��t�g5�x��(�#� ��X�'qi�����}ҷ��*S체��P�AS�'3kv�p��fV�7��^�+C�6���*�㍕�ϩ��g�ۤ�(�W�V3�sQ�y�/�4(pA�����t�zm�u���ש���7�=g=�:���	!��V� ʽ�n��~?���wh�l&�� 2{<�0�|v2���dQ�<{醼��'T����k3�
��P'3Q��*�q�����c,lW��D�\{�����d`�b��� ک�29N�-0 ��#T�x�@	� � �WB�C�́~ʬ�07W�S!6��ۥ��hw�_�b�&П-+���=��L5��`� x(�MLʝ�����	�!J T�.H&S�����LH�.�B�ՏG��k
�kw��!7����)yx����P�s�Ν�;P���p�%͵`�f������T
�}Fڜt
;������*�t�Z�R6mX3�BC;�p�/t�o��4پ���^����������O���׭hK�D�ǆdjxXFG�%�R�� �̈+���Uۜi� ��F�Jc$��:X}��ݻ��eGFc��E#b?��p��a3���� ����J�u��Bid�����^'8�P�p���4r^�&�����)�.�u37暠,l2�
�՘�o�`)������������˥�иis�+!f�'���4 ����jJ�oD��D�(0<�v�YkGm�0 x� t��3%oS,��GE�Ѹ��둥˖3�y���?<� ��x_(��q�{��xgx�&�i <���( 6�=�Bc3a�&mǫ��
�3d��͌�-�􋊔�8���#km�Ь@$,�R�G3�2:���=^,�X!�Z����P��Fh(�}G��{IP�&o��@U�}2�� ȠBi]ꥊ�Y)�&ۄ�LF¶_��/bԵ��\�z$�P�
q!X� <>�T�I$�$h�V{�*246nOYy�@�*��ʎ�%����zxW�a��۳[V�djA�1M���aB�#c2>����^�#r���Ň� ��^sMp�,:�\Np�k� �U)fȁ��G��U|Қj����'�>c�<s�;�o3�[��ihy	�|�̤�N��jo!�ߺy��C�ќaC;%b��a��L� �>�\.^�&��Yy�dX*5H�HB39t���l��h�;���$�W�YP��� �CxLa\!Ԉ�1+g�=��Z��F�d <��R���b����%�T,"mɘx~?���Lc�Ip]�)�ʁW�9��.]d�ć���Y�\��]P���$\��>C����t?��M.�V�����,��=h�ι��R>]Pmq����o*�z�q�9h�R|\����A�I�E�'�T@��Vm]~�~��=�~�\��p�&��a� <�0p�T:�fm��@(B ��M���I�G����2|�c���F_\����3�	HC���y3���[}��~�G*��D�4&4��l����&�edhX&&�����p�WPd�����e�ڕ̿P���t{{ި��0Ȇp~�!Cf�4�:� �i��i��9�P�XQ��MT��h[�]�!�c���m4�lx:���!��5�����@����hmk�¢�U%+������s��c6|��c�|�ܾy�x���.�~ Q�j4���D��*��R,�ب~<|�P�ܸ����{2
R��j��"�JDɁG"%FR�°� ����W�-�J�����gT"�� ���_�I,��uk�⾊�>��.D&oJ[�qc���F���&o�{�d(*UL&d6���v�k�?p�5��	^T�F���'PP0S��M����d+�C)@�m�73�Im�<��aҩ��GT��5�jL�D��Q��}#��p��k�FM���)�k�{�Pg�L�����t�:X׀���g��Ƶ�{�p6 po�H�XX� ��,X�.u��s,M�� 8����84���n��"8h �e�`D�:�BJ���ۏ��Ȥ��	)��C�Ag8Tf�� �%*�%�����+�����Խ��P�����l�f#o^?�ی�i�͞����9Z�M>AL�4{�P����4�g8�`fj.�P� ~��yp�.O�Op�����d<&����R$M߂��w�^Y�z3 J�瘺�5ǵ���e����d�A����f X�4��U���H���k����Vr�5C�u��q�K���P�&_�I�T�K��ˍ��X%m" ���#��H�m�̌JwG��ؾY��7Af����en�V���I�q���$,�@DO���	��9$����AE�_6M��*&��H@�C������R��
�/�S���?4���ؾ���S�OԚ�LOL���(����ݸn�����á1p����V%�/0[�
>��3y��9kM�h��2H�ˏ�_&8�+٦��:��,K����%���Q��c⇊l6$�8��/�+HĨ�-�2�ΔI��AO)��:��$6#��J:�t,"�����tuJ~f��8)>�i�G�)w9�
z5�V#]`���Q}��a}��k<� W���&5���tAr�� ]A4-�gڨ���+(�/70P��O�_���
R.��\�������s�V��pG�gt��^p�t�����5w�{�XF<A�M�+m@�h�A{���������gQh��O}��H{F�J� �83#�H��=���t�O$�5�W���u/�V|T�����̆�L���V�D� >��U����������x��Te�x���y���@'���a��̹(�A�Ѐ!5�8����9�����I8�d���RIҭ�
6�o8=:+`~X���F����������eY�b�\�pQ?|$�HP�����K�F321� �o�bI�[���û����5�r��9q�ܺu�G��B��(3�앨��ͤ�6�+�D.����ђH�A_���:��{����y�~q�_��?ھiC{����G����ش�vZ�P3 ޔ� ��4�e8Tlf� 5D��Q��v9�
V���d3mvр�J�	(W��6�9�g2w�Ȼ��ޘ�7�7��� 1�h�t5Tj�4�>W6C��N��f!�Er8��@�a��Y�Q��gCCž��lR�eX7 p'������ �f[�r������J���i�:1�Ѿ �.ө}t�x �r�@?�T��2����B���dZ��\%і.�58.����I��Qx�� ��4�)���p ��a[��|�3�B�r��> ���7{T�J ����F,4�FdAw�,Y��%ZR	N��yOg�r��mVG]�m��3>��K�����J 3��9�i�M�` ?�S�NQ���^��{��Ij�1�[0�L4oc&�l�DU�`Ta�C��Ȉd��y��xBV�^-6�'`U���1J	G"���RD�X���^I�u���������V-IgKRz�ۤ����Ԙ�EY�r����>ioK�|%O�?����12:!'N��'�Ӓ��Lkr�ѐ�))� ����2�Cvը,`XT~fT҉��t�K�Iղ����C�.!�f��Z&��?���A9��Ψa��imI�s9��<�[f�ƙ�޶e���o�&K�,�p��<l.*��x�3;*�|}����ߐL�$�hBj����(	��}/�K��#줭����*�:�!ar2�
��O�(#IyWx#��y����g_�f�A����~ �$K�uIEÔ��lIɫ^����$� �6t�#؀�N�T���>�n�I}V�w9���тid� X�'���#��!pU ��T��n�F}��]V@��9.��qݬ���C}��C��J�*׸��o�Y��z�g�ɩ�55�=���������)^?�kN��Yծ�l��"�C�
8� �?sI����<4A	劥�Q��f�ͼ?�vY��`�Q��1�� ���Y�G�����kd��r��u���LMMP?�E�,dsl�G�%���8��U( ��iٶy��%��Z)29�,�W-��?vƋw-��wc��jHM̨�,���t=�7�B��k1�S�!��)�O��ҕ����#)W��)ܧd�eVe�ə�-R4�d|�j���"���'�x��_��sK�]�*gN����Q�����W�;��*_9,sZ�eK�����T!kfuvt������Ί��G��ٳ���z��{�~!�B6;$��ˆ�� kN/	^�    IDAT<(4�\l�l��E�з|ys��?�B �����UK*�-�׶��9ɌQ�Q x��И�f�l6ϋ�f8�\,�c��K�3����C�G�e�S�sw�".~˅Ս�LS�'�㳆p4kM���,�`P�K��ke��6���܈�����V��f<f7t5j4�6ӯD'��}�F������\�V^�݄������9͡4�A�1�H��Ns��������j�7@^�� ����v`6�e���dی�2�2��ѩ.a�M�/\�/���;2%w�J5�0� �Y� h@���j�9��B8�� �;0�B�mb�浰�u�NG��ѱ�S�[%/��L�Nߖ���^�iO5�T�92�X�P�!���
y�;�Iwg�}af���W�ܸ)#r��m�5v��)����~���r��q�FB��Ee���c�����e� �����W�7�X����Q[�ʊ�OF�|���8���@	 ����e��c�N^�/��R._�Dc�� ˁJ�Rv���a	@\�H$���[�����ܥKr��O�ũ� բ` N@��&0f3�"�����%;�od��4�:p��dD�G'�/��+��Rִ�,�?*�
���;{؜n�
y����'d��u�:����C�b���H(j*SU��ML��������3�pC�(\���r�qHx��4��Y���ܿsSV�X&��o�����4%�r�Ni4�,�ׅ�3 ��0��81�F;of�C	��3��X�������[z�Y�^q:M-mj-�Qe�P�v I_�m��GY�ZI��,HH�!�������ґN���;�ϩ�(S5�Z*Ѡ����(tm�k���v�UO-J�����ٯ���T�auRu����Zj�(+%j)���
r�:�����^�'���i��}��q?݄�����L�I)W�h�$>G�\��lS��"&�1jv`��̵(h� �a�Y���	����(�|��<�e�BR�AYfM�{U8�{ �r���$�`m3q��4�WJ%R:֮Y-c����P>�اVy�j�%��P40�,��O�e������Ʌ��LO��ql<M�[��{u�j潱V���o�b��`�q�8���&��{�k�<Q��8����Ŋ���˵7��A�AYA�,3���8& � 0���V �{	���@ ��s��ټq��������r��I�b�����?��۷ɇ����pM-�룍42�%~~W�<b���{�(@��̙3O��=0��X�
\�H$(�V��ukW6 �b	�c��>����G�W��|k�D�9~�
���g�u}|�ԿlM�{˦5�JN2���#CC����z]�<�f)�������Ci��nj�Jm�%3��=·*�n@lP#���-a	��21�xSB��V
�8L�9b���f��n����q2�� ��kC��{��ê�
�\g�Y�^7��kР��f(�	� �&��Hpc���𫟥��b�E�\�#�������Z@�*�Yl<uH��Jmtd���aQf"3{�In.3�b'�#�H�ʂ�K$��+�3r�ш��\��� �L"���t���`  x�Р�Qe$��x�Cj��� �yl����=z��]g�@jG[��ؾU� ��r��-�}���M��o�L�L�՛��������XHnߺ/���=�|_�|پm�l\��MR��!�̭[��k�Y�dB.]�,o���}"����iI�^  ���a�����]6�\,�~�5����Ǭ��,G1��`�%S)�R5#�6��ƚF�Tku�$Ҳs�^9�ʫr��y���2<:"�t�T jUNKĴ�RvJ*��?�'�~�
��*�c`���%#HS���'r��%�ʕ8}����{ cڵ�ǀ24ia���rnZ�c~y~�v������ݤ� ���4zu��G�����r��Cr��9��Ѓ���m�u�6��z��F{kZ-\ �BVn\��L�w����&R.�%D��6�L��>��25���FPq�����s���È��P�'@�)t9� ��%�%�����I�Z���m�Mar�*G&�Y����*�&�zYJ�,+B+�IM�3R�~v��i��mm�s�&Y�@�H�"+�AY��F����l/��c7�/�����x��y�(���9����2 �PUݤ��'hf[�4��I���=/��ǽ���ޡ�����.�p�
�{���67���n���:k�Y�c�=��t�w�_�^�2R�	��"�6�1 #l~���S��/���9��� ���T����tg����djl� �C�EPg0,� ~���e``����J�ݹK�^ߚH�xp�A�)P��Qڶ�5){v�/�X�V������3�u�����vݽk���4] _2J4C#c2<:&=���q5��pX�Ͳ\��:���UX��Q]+����� �X��_�o�@��'N��ӧ�����������;�r.�ǝ�晡_�A, �%���-�����`���.���� Y	XY�0Ѱn�Y�z����U*6����S],>����}?��|��:��3�����3����Vv�r�29�Xʹ,3r�F� r`��}C�7& o �u\�7�gS6����ƣ\�ܸ����f�?���NE����F*��D,�@6��f��d�zE�6��C�q3 MCk)5PͰ5�1�RT��
���o����r��Qq�� �N@�]ш]��^'f�,-�y�ArFo� �|C� ��x�B,l,\�;�7 b�AD
#��w��g)Wz?�;
�� ��@�R�&��&.�t�y2]�[��TPa���mJ"��se�	൉�( ��H4����K-��?�f���vJ��B��T�$m��y�8��I���%�2C�w�.�O9,�N�&w}��M��k�I(�s�.�b\wwW�ܻsK>��?z����@_��x��u��1�՗_��˗��}{������S*W���҈�n�vWȒ���q)���$�'��G�}����ꫯ���8'�<~��f��nVy��? c0+jT�ZD�����b�e�Ny��+r��5y��������%��@�9��RVRѠ����%+�!s�QFQ� s(��#�x�=���q��΋�TU��2�l� �fU� I��}%ya�Nf��-^�c'�!6�b�YOQM���֝�����DK�T�D���vٵk��X�����ǎ���K���wwv��Ĉ����m�&���W�V͛a|d�@"3��_pO�=xH&�2TF�f���ޔ���R�����A�� �f���l,�Bi�,1s �eG��C� S	 �Lbw��c]׫��LJ:�5�V��56�X�:���5�t".;�lf��"��Z�x��Ra_�up�KW�}#?��Ֆ�MT��R+ݪ�|����*Z�7q�rM��j��='���������T�?
�Y1u|�����M��[��n�^�s�n�L]��U�$�����w}��G=Os��k� ��� �'�a�Gb�+U���s��WGel2#���RRU(�[�5R���!N�b����D�B�)�`��lߺYV�Z�>�/���:��A�r��lM��{�R	�x�8o4��߻G^zq���t1������lb�֭������o�H6{1̽�D[3���t�k���f�ל��r�s1 �P-�(O�F(g;4<"����@*����i�U���U^
$ؠ�xÊx0`�>ؗ%Kˆ5+�Cp���p��yY�r�������_�@~����r��&L�iǜ&�JȮ�
� ) x@M�V޿_R-m\7Hd��,��&�x��%����+e�򥔼��?�֬dѕp z����'�m���>S�>�?�/:�Z~{�����Q�z �b��x�9�b�� o�F�i�r�1a�df+��fҍÅeK1��32H*�h��p�p��'�<�2��,H�l2.�L����y_� xw1z<���J6��ǽ���ܳ�FQ��7�`l���k�ۭh�����ո5�	���:��z<��0�lC���::���:0�E3�:' �y�[d;̹�.l�:i�*'��.1/(��i���^RhO��/��T�A��¦�u�A��j*�
� �����(��6I\5�!�ubC��|���r�?��1�vC�/� �����%���O�đ�\C�,����k�`I�?u�����l߲U&GG䣃ʑÇ)��ũ�`֣��,���ʁ��h�2j�^�xQ��]��b��F������`j�E%MH�5�����F�� �V�&����#��!�����Q��=2@hi�y]=��@�ȱc�@Y'��-[�ɾ^��W��[o�%��?�b�h��i�d��R+�=�?��kY�f��Q��B��7�h,.��G������3�Έ?� H-VLc6���:>\����e���������K�Z�|b�rpR����z����r��9��/@}{�}���b�*�p�|��WF(��=�w�@�H�,��iY�n%<
��J��r�B �N�����g��߼�_ �`���D�U�A������k��� ��!R�GA[�?�ʑ��(zd̐�2}�&�nG�S��S�K�BE	?�'@z�+�-�{? P_���j�ӎ�[daO��n9�P� 8�
�鿱S���"���o��j�
�UMnx�2�w�\��J��݄�f���\���|k=�{,׆y}��ʽ��}��j�5M4������(�	�w�7�ag�8�#Ļ�4�\���\���s�g3��c�1��� ���C�&S(�	YU���M� �}n�6���8� ~tTj�3���<��R�^�[�o�.+W,���9z��ܻ{���s�je�=35-�|�8��=-�vl'�_��C@iJ�Fʒ��Q�5ЙIR'��pE�hZmV��k��8Ϻ�M�47Ԝ�% $r�������Af����t��%��FT�����$i+� �l<��^�@��h+&	Y�f��_���Ӆ��9ͶZ)�֭[��c��c�wޖ��/I�XbZ���#��uqq�ړÇ��)#o\�K(���v2F�\�T:.kV�����%����� �
Ət�k�I�ҍ_:��>����}�u�ė�����5+�u�&�dztP��
#F^LhtSs��̊�m�y�M����7X9bj �i>��?&R��d��X� �c;9=-�c#63�!3^vS!�r3��w6#�d\��0v!+�E?�`4t�φ�����J�iz[�jd�g������l���x�:Lר�u�u�)��h���o�sx�ŉxOS��dbԡ����kF����zQ����]|��kh�5c��$^ xd�ۺz��{�t�̗p�]�f���A��Ę%�ǆ@	r|^ �F�ư��ANA��X��犬J��Khl� �c��2�f��Cx�Ymh��YiMV�FeDuN8��XX���A ?=1.'������-��m�wJG�<9z��9|L���#;�nc���_�-_}񹴷�6Ԇ�5S�S	f��-��H�GF��e���r��5���OdÆ���K/2�
z���ed|��� _�`D�ݹ-S����˦OP���~���`$O�
�ysf"* {�#G���������$S-�i�vy���z톼��/�ν{�)�SG���C��
ґJ����T�۽]bQ�p4��9���������7�������ū�0�/ܯ�G�����,^�$�\Vvn�,��w(�ׯ_�(!�:Ѩ"��~X�Wnܒ��������/(��"��L�"�f�:�\?z���7H]���%K��QV�-��m�6Igk)4���%��l�H8*�����{�@�;!������6�|�&C���'kg��~6�! 'Ӭ�a��Л����U�!fߑ!��xp|1|	�J��/a��M8 �g��_4��LOpT= LwG+���ٱCz�uс�^bԩ�{`�T�kW�,ʧk?���`{_���7��_3{�,���9�r� �Q���N+�V���>��^���X���u�]?��pk-@�1t��J�Q�� �]�k��}�签Y��� ��3�_��&��s���i���0C�Ò-�ɁW �7o(4��H|�B �" x�_���q������ǻ:��޽;�� �H�ʨ Q�I�b����2��Q6�>��,[�g��<�Z�i��H�ه���س׹ P��a/������8���\+�{�ӿ1uC��=x$�n��	̉�JR,���
v��l83��Ġ��&"�C1J�����S)��زa-Y gϜ��׮K$��{N~��QB�g?�k�u�6���Ɲ3�0nҭ������� a	<�%H��媴�&Ɂ_�l�}��'��FB�/ۻ�����_�?��}�=�;���k��=Rh�h�@Gt�̋Ɔ�����ANeۜj�����.jlh�6�ݜ���m�Y�R��w�F'�gO��djz�)�5�J)i#L�ut����5
���r��R���>��g�dT�Q?_�~Ө4;^� ����u��������]5�������5��uq�S��*�gww `&��fce���㽸� d0P}�v���`n��( 8��Af��RhZ;��{A�tt�@�P��d4S�2���<�փ�78�0r��aY?Jz�@��̕�wu���U�?6�WJ�;i��c�dR�X>�АGC!ټa����^*�?�j�˼���g��L�˩3����m�Vٷs7�%o��:�� ͸���H]z�����9��5��x,"COebdX��/b9���ҥK(�՚N���(A����ˢ�>)�d��ׇe�ɠ���d����LߋYg�@������_���!�P��MVv�.gΜ���P4�aN�xB6o�!/���\�vM�x��}���*΃�@�&!��+ߑW_zN:;R��a�h�!���/6��}�q�z��M�T�$�yp~5d�ͤE ���*�;����ʫd׮�ґJ�T�� [C}	�d�/\�&��/���SFn1$ Fv>�j�l���+����r��56caP���(�	 _��d��U���4SIU6�:������/dl|J���D�iR_��jBbÙ��0dgs��Ҋs��$�J4�"��Q�B֝4�P����QN�%�~�jɨG!��������hZE��N&�%�d�1 |ƥ���}��lZ����kY3xZ�UA{l+�.�U��~���^�i�@���ךk6m�@%�;	��s1�9l�&� �S��^z��Dr��S}�&��c7�o*V�Z��f�]������`�
5��:8Έ���7 �^U����\+�A�W؞u���?q��|��1��!�R�1��n)4n�U=�,efbB�X!�7=.Є�H�T�L$D9�!���v�Ķx�b�l���|��2��h<����JK�e�ޝ�rY�D#؟�>���W�}�B��:3�NX������y��7���� o�}�ǉɌܾwW��}H;
���&�k�٠�o����1�˲�	k �f8L��4׽�"�u���eK���$�˗��ի�D �|�\�����r��U��Tk&X��P����Ԋ���}��	��D�I�+Bx ��-E���^��va�<w�	�?����K֜�� ��}����>;��}��,�v�޻�&�@�L�º�\����j�[����-�����Q�1,fS�=x�Q4�p�U`װ�Wc3��\M�bI<z�E��d0�����\7c��Ai�xxj�l啚��¬��Z��~֐���I�\�v��<M84��f#u�PD�f�Y�ª@�gk�R�-�\Z�w��l�`����NN3Z\ءPC�	 � �\6 ˪>�Ln�V��Z��P `�3�*��R-���']=���hFd��{D*Ȗ���58��!(���5N�C�w� ^�X1���rj�    IDAT���`�{����U�M�4 ߸M6���x��\�o��h��N�ARf�b��A���h0 �xD6�[+^x��BJ���M�1��*�Sr��)�~�HW,�}��p��/^� ��J�#9���*Ӭ[���l��[��c��G�}/��,�]@#=:1�5�� ܿ��3�����h!�5�@��1���j�jy�WȻ�t�Pf�ڼz��?q�j: ��d��_< �\�7�|S�?x@#�5L}�2u��\{:Zd�����{E�Γh���U��A�����o�+o�{P�ǧ�\���:���`����@i�~t�t�w���dݪٽs�,Y$�b���u�*οR���7�o�zG��<��l�B�xP�-ZB����)�" Ԇ#	��R�gdx��/Y$;�m����fI>1��Z�` D �o��?#�G>�JI4��@$΀��H�X of��x��1���I0b3���T��B�����k;\	�?$=SIiO�5o���5c�Y��G�?T�l�u�C��
�����e���"�,�>�*3j���1b혗��ث�j�1/(n�s4���1���2��!Rm���gU��~k2D�&N�租�����a�lUZ�׬��W\���H+K�Ht�u�Oό�}�\����}��Hyo�]��\U|� �F�)+9�!�
����oQ���iNb�6�RJ��HI,�rI2���+Ux$c��+��h��R,��U�T*)K�-����0A��ɓG���ce�? ��_�W��r$ ��ze��]�~�j�E�l�����+�}.�HGh�):�����G׻�!w}κ�v�a�ւ���i�����*)|B
�?k�M�g:����!^�C��+��;�ӆ�8���Blb]�z9�PNݳ�/ʎ;���D����r��ڊ�y]Lp 0H�S\�C##л l��'4�A���Q	������A� ���E�/���k��ѯJ}Uի������z~2��K�6��?O�� ��������b�c��=����جZ5�~�&�ۜ���S#JoLz�]�эH�Iv��f��y"�`hh���M)��~l|R�>�/�C#�i}��43�, o���V0��Y�;���mF���N$T��0�n�ƣj�ܗ���0^3�1gk�t͟Y��fklF��iJP�=�S:{��Q�ׁ%;�,���p�k�Q��R�;��`��J�Q��Ὄ�+Ћư���FP�G+!����t��y�=R�d��b="�p�SNǃ�6��1@&m֟i22x3'�M~\���&�����04�N2��w����\f5�*@�~�M�����3M�5+q��oN�C��I��3�W�5��m[6Ȟ�;h̆є^��P�hm�Kׯʡ/>��O��۷��_�۽W����Ϳ�9u�t��[��Җ�޻y�d��5૿���ҿ���Es��s��/?c&x�ڵ���N�"�L�h �B~��ݛ���g�D"Q6afrY�<�NKO�<f�/\8'ӓ3�{�.ٳg��Sq9}�,�L�.7nݖ���J$�P4Jc�e�ٽw��9wA�~�|�U��ѳ�����z�u��=�?��,�cv�� 藇���a��:��;����~ cYj���:����$QP����f{��댉|h:۲i3g��Q�t����7�ț�/'N���kƐ����-��������I�ʅB��X����<|pG֭Y%/���-\ �,���?1�	��kx��	�����UfrhF�H��6	�RTy� ̘�XJ���m� �s�D�O����PݪK���_t���p)/m���]�/+�,�zX�V� 	�b�đѷF2=�
l]��0y�1d�[RR��d��%���o`°mf��0���`���1W����U��f�ݿ]���Z� ]�������S��U��f9]��&D�q}��n'q��l���i�^��>��{��(�	�4X��s���q~J�l���X��7I����v�O}�V�7�p���.��sEu�(����R�@݅�7U�b	�9yN>���_4N�3����7Q��5G��  �擓(A)JJK �H.*��b���O8�n�����"�S�28��ͬ��f����Z�Q�ǊCP�/�7�[^xn��_����r�T���+�i���<��@:�H�C�uב7�r���:E�x��J%����Ƚ{��P,��)Od���l���=I �n�0^*c�E�x$Mpܶ�V�j�0�#�O-�c+�'�o]����{�.��~��Y?����ʵ���B�����	�uP��w����  ���or�`�(�A�9�e����p�ݧ%lU�H4�N��t-\v}��n|*���~�v���g��ޮ�߫s��� �줌�����@��A�1Q�M�t놤C�\b�-�k4��d�a�̈́N�����C`*'##c,�*��s���%��o�|�A��h���Eo 1�c��~�Y��9���v��3�����7Po��ó���z�
��XnD�8�cP���T��([6���Z����22�T�B�M��
Q�)��l�;���{�L*2SK5�`$F]^�x�� B�QG���&9%��P���kF��q|T*�����D����TV3k�k��\�,糙o�(�Vv��/�o���u�Xhl�����*6��D�Af�S�lݲEv�����~���R~p���M%����r��Eimi�͛7˲��251)_~��|���R.�e�~ٱm��L����ؑ?�a$"��]r��y��7���k�6I���n!h`.J"����y,;��λtT�V�1��8_"��i/��\� ��\�{wP�~��}�\}��6�o�����a�r���')ٲm��Ϝ?'�|r��LDct���K̒�Q7�߀����Pvl����@9�1#D`�ɮ������嗇edt\�h����Za���0/�ic8�G�V,Z8_֮Y%۶n���J1��J	Y&h��HW�>�|����ˉ�gŇ?��,�8�m-�.�9���xHr��#Ti����_��,]�fcd��-B_H$�B�(������+)�˜���$�j�@$F.�ʾ�M�� ܏@�*%$!��DK���q�C�A�R`����Y��M�_�zaF���|��~ٱa��sST��DJP���U{��R�N�?x-�qG��S��Ẵ����  0��R�w��f��Z���1�e�i��9$���IoR���n�K��A�&��W�d���x?s��'sx7��� �ӵ�Yr�N,�`Em�7(p���_o�\�����4R�nx�f����1�5��~���
�U���4����5��S��"�K��\oV�G"Q9}�|p�y4<f��V�I�"%�d)?	o����`�t�$�H�����`WT%� ؼi�l߾Uz�u�\�qUΞ=m�!���|22:���j[�P�
�e��Rٳk��/�D�Sش�
�6��/��^+�q���������'7/q�����}����Q��� `�J6�������ܼyK�'�ȉ�MI$`��/���j	��n��&�<���N�K�5��^�R6oXK;���ɝ;w��o�<��>y����͛���t�RRo߸̈́	�I2i���PTV�]C����'dtl��b#���/�6����W6n\/��$P��B�]�	?�A�B(y������-�5ll<���O����̹��������L[ef� >73.�#��ňaʣY��6�8G�� s3�!����H#y�G��j8
����e-H���c�2��Bb����!�D�$� ��|�Bv�\7b�E�����{x�����@_o�$��N�)��uz�fA�4�f>T����m�	�;>>��x�!#���N��������	I�[ņi�U9� #O��;S(sk�P?j�#9� !��c�3� ��|F"�à�#�
"_ ��� �B��_��]C��~�jcK��c���&�K�nI��M�e��M�v������+4([�m�U��P����{�'e͚U���\>^���S�w�&������;e��U4�<�{���W_}%�m�k�yx��|��Avޯ[�Jb��[.Z-�yB�����gF��� �BV��V��X#��[���m۶����g��q g ��L��� �x���[6ˎ]������������$�I�vTa���싡*��Ɂ矓;�HWg���fz0*� �JEFF&����r������HWb�Ԑ��:�jMV� u����ŋd��U�q�fi�u��s�T���"iA��H.\�De�-��g8�3����١p�\[8�t*!}}�غd�bIDu�R�Pr��ezfF>��Ky�w�X�I$�$������E�M�p�hp�7`d�±G��ꃾ\�r��I���Ěa^�	��IQ~��s�s�:��r3F���)4��@��,�稄1�f�0�:�Z�� ��Ye�w
��*(Ԋ�>��֭�x�,��� x̀{|�ƛf}��ߤ*���N��X?��<ח���X���fpi2�����J�ּ`�����2�kJ���韚Yy����fx�^�1t(	��cz>x�o� :�\r�1t �jR���ȉS��O>�ѩ��"Q��� �߇�U��l�:����IA&�~2Q%ڼq�lٲ�=J>a�Ν;Gi&4�#��35��(�0�����ǽ��S�l��x2�Nߊ��&U垁N��?��;zt_xף�9����*H�Ü ��޿/CC����elbZ&���S��h��GЃL��m S��� ��b&	��Y3HjEH�ܶa�9N\E� ~��=���/��[������et|�� ]]�2=e�*V�����,#=�0�X'x�G�	
�{4f�������NN���G՘XϏ��Z>������/���ߝ76��Ӟ��?}���K����_���Z�"�����0b�
����\`�FŽ����(�%9�=Z��ͤ¨ߔe&�c�1d��и��i���|6��}�������uV����w�X<�:?��{��]q+�c<�}��#�ʹx���n ��5+䞫6iS ;΅ #a��ѠrBee;gp��g!�a6 ��-Z�J��V������d|&+�H�<]d�5ɗJ�����PV ��b,��g&� �6���Q�1�n3��0~�����=g|�o5�t�΃N��z���~0���Ȯ��VHa����P��$�/[j��.Ï�Ջ��������N���H�#4��o^�0�U+Wȯ��d��C���we^W�lݶ�M��l>xp�}+����!Ź|�ᇍfu�r��޸a�Q�p��#X�z�2���_x����!�Q�
�5����>�x,%164�d󶭤ݜ9sJ}��d�'9��.�!)�	���)�r��/���%�F�u�
�Q)*IB�}f&#�|��{r:C�k�śc����^�C�p�|fgP%�5�ǡ8��0��L&/��?$��)���h���Fv�@S[.3�@�:e��iooe�BϼnRM���E5�:��W���R�b�,&^'%OK%%T�`�%���5sHD���FE�k�Md����Rcv�:7����H~ZR�*��uk����bv����8l�A�B���_�1mDV�[��������^\s���ש�q��k���x��5�ͮ�5��ٗ.���/j��O�x�Hk�]���ѵ��/U{�VR��Rv���~����U���q��{�z�\0�穾W7��� 7(sLz��}
��<q��_.6�Ee���٭:+(��E��?+�}�������I	*Q��$��y� �t�\V��F$T��A?3R.	�X�]�R֯_GE%4�^�tA�=��� <�+ ���m3��X�h���򋲸o�Qp�*x=Mͭ��w]3��Հ��IP����|���y�l�k��dU5&@�'�����23�㐭���с��ͬ����"�?ۀ{�L���������a���P�)���c�:`�z�nܸ&���w^��_~�~�/���drx����;_F�G�t�}�42Thp<T���<u��c�Ҳ��'�q�[P׭['�;�_/q�$˸o1Ư&�h4��������^��]��_��h�~$��4)4�3�R�T>,|,B[�w��{��q���j8�ɮ�&�r$^���� ��M����ѐ\f�v�y�*�Nltm�1͍��T�{�Ε�x�B�O��{�:ҷ�/��7\C��K��n���5��i͔����?ב0�d\�}0��2 E6b�o�ϊ'R�l�Rټm��޴����ސ�����Ԍ*u|(��p0��PchlE�#�1�'�. xppI�)d%���+`i��3�^ ߐ� Oo�'�4��^�g���-���Fv��=���>e�TX0��q��_�I=�'�$SqՒp8Hm�i ��!��s��d	�?�π�����fg�8��kߓ'�ȡC1c��w^�\���!��}G�,d�, <4tQ�\�h�C�(B�t9�7/�t����l�J�������h��1�y���!_��t,!�w��ɉ�G�ࡃ���  >X�H�Xf|ݪ�����^�H�*G�*J�B^��dsy<8,����pF(�*x0{��$xOBA:jp[��,F@��ϑ� ��#��Gbq�fr�dxH=���Q���El� ��5�p��|B���z�X>.�\WW��^���1L�-�XM0�Q��~�d�C���*rQ�*!u��&(�A�X��o�����u� P�	d�)�G(�:�LfT
�!�߶v�T�9��(�7f�X)0 >�1S3��a���7t�"�;�]ڗ���ˁ/6+� O�0�W��q+��Y7���s�>���&��}^�4</0�@̦&�]v��'�{�kNכ&��`E߫6ۭt��u�����7��|��n�`���n�*��&��zmB��H�,�z,^����`�tTqf�!ϡ?5(�hGq^XS��i	�#'��ǟ�D� �`�%�{3D~6��9|T�b6� �hbż	 x��������dŊN^�r���q&(A����G<'���������iV>QY�Z��C�TA���/0_)���5�o��3I�38���V�\?��!&�b�������A6� Oe�b�cSr���d�,��Ђ���^#�`N��2��5�����N�����Q�aQ��$�	R5��z��{����K��߿O8 gϟ��_�Jhjؒn���o�j��	���VQ��Ҏ^�tY�9����
�O-��G/ <hR�F���e�~��������4�?�^���3��Ӟ��_?�q���?�H��^~b�u��]�O�Q!!_�S�'��N�n4�<���=Fx����r��l��L��F`n��l⦁urs[iI��Ch���m g��н |.`��b���c ��gn b�c(�=�|���iu��f�Z��]e��C��7���Z�aG߇���}"I�ZdI�"پ{�lز]Z;z$S(ˣ�a�|󎜻xI��'���!���́<4�BQ ���G�n6��bB(e5��Z&�	T�a��f���� ��(\�=��խþ� ̫a�$E[�gIQ��t��jHD
��d�D�H4�� ��#��Y���	Ɍ�JHꒊD���rd��j�1L����O)��=�	��޾I�-�7�s������s�6�d&��eْ~Nu�xCd����!��~	f�������}��{����s�p�"QR��=|D�P8�`$,���=��ʱ�Ɂ��2�y�fhz�Fx8B-`�>�+E�#c�kN�Q~���X�?�!�>99m�\Hc�f!>M��'�t�e`�Q���Mff�%�ό�.�*�J��d�R� �`��w�L�6�]�]�� �pL���C��iG��|F�
; �ࡂ�	*�h$ �DZ����Of�T��t3���1i5F
CU��A)c�a�mD�z��a�H\s�O�R��a42    IDATOKG<@ �e�r���~�� o~��x?�>��ޫ>6l�*� 9�p?����]�r\KWE��ֺv\��p��R��b^ �]j@���F�cJ�qm����
��.�.��W޿���S ���j����{��/�q�Z�8 7�Ev�#}�^O=~��5;5|�M� Y�3�wb�zy�f5Y�eE��_��{\�3��Р�����g_H�P�Z �e����f<y�v� <�p�̌L�|������zE��"V�!��pa/U�p����'�|b6��w������|��a����s�>��MW|�>���U��5��g�S^ﳛ��x��u��`+p��=:2:I �˗��C_��]c����A��C�M�f��	�4�7�f́[5��۶�����@���	��7C�m������G��K�,adpp���x�MI�����%==�<��KW��G��$J$��y�'�y xPh��u���8T9�M��j-	E�H���i��ڛ���OM��_8��������ZGܖ��(G}+Ex\h�s�K����W��Q��H�>.�n<Nγ�D� z&�#�F��ĳ��i�u'���x�.�x'	7��ꊧI���� 8@ǿ����x�\���Fr��7�p���\ѵ�p��jp��X*�i@ M��BX/f�C����JZ��{����m�w����c��
��2>������������_h����ѱvA � ��&�B���j9/Q����if'����T�, �����Q������ɾ�1���Vr0rFƠJ�h�3=	uP�� \�J�����[[%�r�Ѥ�����=y"�zM��X[�j�[��G�ebbL���.����.�S����ꯨu�q�����B�],�΃���6��niMK>�#pŽ�y��⟂5T���'�7m��FF�t���3b�\^"�$������۷��G��>�
���N�D�Ä�e�r��(��c7�h3H.��J6���ESb*4<͘m�F�ą}>8��Ӥ��6`ŵ�`T@�3yI���[�Q�;�6`�R+����s�<�J���ר����,��R.�=�s�7�$M�c�PB��dr%��Z�,LG
�/t�C��QRg���?(���Q�x?�\om�C��hU�MIO*,����y� <��ԬW-�߿	��Qy�SWe2 6c3L5� $M(�4 �9�����؛��տ��.�q�� ���9.������>vsR�~�7�������y���w��µQ��^\;קz��\�J߫����ߛr�&��\�	!�]�Yb<��n\:��O���~_�\��nHƨQ'�� ๦������ɗ_��!��l ��� ��u��T�8�%���ꒊǨr�~+���Jgg�,Z�G�v$M �@�ܻM|�Rf RBs:�oM�*���S��,Y"^�/kV�`w_�ˠ���A�����=�5���n��{lZq6d�����]���$> M����r��-R�D69��9�# VL�� ������1�	(iֶ��S�#�[��~ ���sV�Ǜ�O��p�q��W1��@����h�@>�j�o;�"+$�|����<�1�:�J�[�V:�[$�
�Ƈ�A?S���"o���=��/�Q"�g�ё��w�I,2��g���Md�x]�ޠ�6���.���\,^�Z����(S
3Q2�s���G��0���Enh�\ߧ����^��~����u�P7��\�3t��gbc`N�ᬩ~֦t�~�ˁ׆:�?$ )�`L�,P�k4~ �b�����aSZG�lܴEv��CJMQv "!�BQ��{$'Μ�'#��]@�&�r "�r��xRt,�uF<3�ղ��rt� �Gc��Թ�|�f�h�{�i��e;���ʧ>̻fGлk��w�>�A&�����\'�t����ju
`zBpq@H8,S##21<$��r�N�4~�M����S*�eb|T���)��믑����?��g�0ۊu N3� 3�^�\;��
j���-@C����G��*8�����C���A3���)� ��q�zX*�Ϝ��rG�DD�q:;\/?t��dh<��j! o�3��q�� �{o2� ��L�6���~��vdT�D��f�c��7�(�Tw����(j(^8y34) �9�ӁW�t{���JPM�&�Q�/�I�P����̆AF�2���"B_K�rޡ.�;��X���30��������j6C ���_}�ٰb)��pphңm���q��9p�pܤX���T��{��nAyӞ���:�6ҥ��:m޿onM����*;������v�Q��j&�������J��3q�צ{��c)�W �x<�t�{}Is0�9/����\���T���u�0����ք��^O�����r{z�� 
k���\�㣰�#��TA��H�X&���G8kfv.��*���dz|��C�3m˘�,2��K���_Db��5��
~7t�QA�ZF0Q��A����e�*�.����_^9�^��h�[ �ٞ��Q�*����9ʻ����rZs�P ñ ����2e"�QY��&Eqd|B�&�@j�A��E���M���ݎ����� (��G{hV,��[��@�R���TC Qؒ��	&�I��Rb�v�� ��㇬p���t��C���D<.1P31#�眊e��Ia��!$�EB�bZ __&��,���KVm�3׵l��=�?���ĕ�G~ojh�m���W�R�����8�G(ߠ\�Rh�ƫ�po�n\�5�<܍����6>jf �3Y4��&w#� )w���p�̏C�q�ˉ�v��� �qK9�j��9���{�wK�^�^C�si��w>����1�j�԰�����<�rD���B�f����Ӭے�f��&�s��F�`K�p� w�:���5M}�v�0C�-����r��9y08"c�9����%%[�K�d�h ���gFG�V)H�.1D�ANP��vnO������� ^�/{3��3�T F@��i�# �>ʑ�M�� �����<�q(����˒���	����&|R*��3'/x^^���)�x��m�y���Yso�U�L�ȪL��4![\���	���y��0��N���or]��Ƣ+V�{�L\(h$n12�h�k͂��==���"/������ؐd��I�A��`\'� τ��+J��[0�sd�Zb�:��KVB�Z\og丹5�(�Ff� �gd�`�	�m���J;HAW�Tvҙ;�kЧx�����$fe��B`_��Ϯ�J� ���wA�	�`����|Aii�Z0$�B�I_4�� ��������+������E�P�"Y�b�Y�С��AR�z~�0��1䁍�%c�?���ǆ�1`<��4�:�ժ��sN�,��bz$_���`|k��uϻ�=v���W(�{Ͻ�}�^�[k�[���ꥃkH!{m�r	��z�*�ҭ-I�Q��3e��?p�~7�F]���Pj�>VWc=B�ık��t�J���  ��.>{n�0��{���G�*o3�]�sc6�6�΃^Ok�z�oGҧ��MO�2&�p-�;�J>�a<��&��{�.�1��x�GFx?��>�l����}��U>@ �gV~��|���6���q�N���������^�~]�H��x��j��GQ���M𠻠�p]�W���K���[�(u6PC)��-�iVwqeY-2@��ד�Z]�
�Y�4;-S�e������/~Nu�;ʁG�5��>aK$�	ɹ2�����(L��|���wa��Bt�F�Ԕ��e����2���I���K����s�
���G&��S�!M�͚unk:v�ob�/|�|���/{��U�ȅ���c�!��@a�z�6RY�/��5
�u��&|�V��pH���$�y�xR/��s:x�.A �M���؇y�۪[�R,W�m�P��;��hݱ�& �K���v%���K3�s2h�5<��`�,裀�zq+�%'3#K�u��c�@N�c��Q` ~�뱾�E�L*|#�t?j�����ҕ��Q`ُ�xX7?du����!���z����7�u���
�����k��1�`�=d�aƹ,3h� P�ǅX��ULU'����=�+�RAF3�4 zIN��(?y�99{�t�E���:"��J���!&� �ۮ+��5Ɨ �M�<�_�L��:Y�ለCh3a�k4F�����cl����Id5-|��c#��ʩ�	2��s���L+�Ga�d�,�TJ�]����%��I]Q��L����j�t�ɗ��9ٶe�f��0��X�kX?���5emq�lt.'/��w�}W��Q:,�̺:�BA��͢ ���Ma�zw�,��S�!�f�\�pN�{�--��#h�f�@u��M�S�c`5�=�`�N�Z{M��e�1vt�n���Z\�� ���(<�F�04f�2�
���w��5pѷϣ�+�z������Fӵ%aAY�P�V����%�-K��lQ���d+Ӓ.���A!kJe"5����yG[�\�S+��ےt�)��l��_���~kUR��T�%��P�� 8�V
tR�Y\XV�� ��`d��;���+�`��'o��r-я$N�&m!�'������u~��[�����]dKrXFџ�I/��Ǳ>cN��$
�N^�_cW��f��Z�v��k��k�c�������\%�	��T���x��]{ܯ���_�<����Z��U�'�U�M���/�K��%����y���h$b�^9�Ь����|��'���Z��4d���y睲��$++K���W�]���ռ(�����Gՠ}���R����$di����*��x��Q6p����sJ��5��o_>_>&,aa���S
5;�xn4-�t�悜=w^<�4�����W\�R� �{}]�P��� 㺫���"�.�nj`��^@+���1 ���OQ�&��a7�v{�p�Bx��A��׈.P��������w��H6��F�.�d�w;�P2+��Ŀ�NT��]��8
D�eܛ��?9����I)��������V��ִ������K���El�^r��	�"V<\x�Ɂ���2i\d��cG;��ꁳ��_�v�gԽ�z?i����8���}��G�cD&��4�ttޑ�5�H�y������6�7�(*����p��3k3S�r��ʑ#GtA�.��g
�#C�3S,(���7ߖW�9&�-ʠ4!�;�&���%��" |�U�d�[uU���#^O*���N��|��M�X��VZ�}�yb�_�'�R�]��$��� <�;�reQ�X�׍�G3ӪB�g� ��ܜ�&���QC��V�B�����r����{�5�*9�V*���a���S��p�o�І?}��r*��̌��:W�B��D��"ۂ-T yd�u��Q�%��t�y��m2QA��;���9y"���88Cm�� /p�] ݞ�5�3 \Bkv\#2�
��?]@�Vd�<C�]W#�Z˴��L(�2�:l�Q��]Q�kl��ꥠ��V�h��T��Ѐ�,~��S��M��lY�9�JUI勒*N+
F}���*3�K
NE�v���<:o��I!�k.ˎ��xPh�0ũR.X̷���*�H��Կ����Yx8f�}P��C��¿8+@ �Lr|0���p����ɢ�br}���|�Q������X���k��׬�� �Q2$�߼/��s��}�Q����� �g���Y��҇0;�qL�V"3�v�y�qm��jTJ�h��+0��jQ"�"m���F�/?}�Ey��7��<:��#���j��ߑ�j]V@�AC��e�a�KR�g���Ν�%��J�Y���_��u'L�F֔�0�Z�с��23+۶�����t�o��\R�PJ�i �qL���^����G~L9����y[��%����s���ea	�������S�K%k�A.� ����u��H � Y�[�dB�h�ԛf3��S6o�e0:��3Y��5Y��ģ���C�v�U�Zd^v�ة��w�٭E��,�]�{b�tzH��VJ����)���_�������N����L��-\�<[�ix4$@�[8|]�ʯ6\������&�ψ@F��a3��Y�$�g͡�p�g�����M%����� �(#���ɱU��A�������sE��|o�i`�k�%FsA�W~/@"��8�ء�<Ȣhvt0PI<��������C���M�I��E��A3(MLʅ+��Wߒ��9&�LAj��dʓ*?��?� �r�C��b%	 ��_���i�� ��n��!u;D뭇Q�ߟ���=�`DŬ����U���>_��̴+U�Z9/b ~Rb��P`�d4۫ ; Y�o@V�\�nt,��~g�EX���=�54� B̾�a�3Y���FM���/86�}�N���*����=���ez�('� ���\�rQz �˔eS�� x�;���Khgţ�Ȋ2Z���� �	v���M��8*`t5tv�هZ�R�⎈t����1 �(2E�=���	�f�uG���f���n/%��@:����e)V��01%td�M��{7�wԬ"So�w�m6@c�[�-��`g����5�d� ���޻����2Y)�T�����/�ӝ����*?��<sdضlަ �2bF�A���4`�7�3	��
Ɲ`!����I&/b���'m7�k�;��	N1ǒ���d�'�6������`����?��Q2��=�J�����6���y�]��i����?o�x|����琉����c�Dv�4�[�����p�R ����Ϟ}i�7�V��-�tW��]�^[���u)�
౳��::u���<۱c��������S"��M]s�RQ���Q��$�T�*۷m��GP �DE�Y����]�9�`o���~�毷a���_�;8ƴM\s�Y�/� ;W�������r����Ҩ�9�H�X�m�"���~�S�
�ְ*d���P�B-S����:�*V��͠��J���ĵ2�A�vT��H *��v`y.�&(mU�U]C�ĭ�g59V)�Vb�Ԕ��(�K���9�g��ݻ|�.>�& �����v9S����˳���C ^�u��L��N�w�L.��.f�{� �7�I �9���i�'d�\�L'J�Ck�:X=����QFz�$�����ā�0�O�a�8JS8�b���s�
���g|��Q�>�hx->�.�)g�c��EFXp,t����l۽��'�>��lٲ9 l���a��ld�ڃ���#��+oȇ��W�H7m���iS� �_�>'��,���V�!�z� ޏ�8 ;�X�t��?���s�3;�����)L������� 8�S}���]�J&-e �P��PA@6��p�B�R�m-b5Ko�@��2�!���c�[��Z-zBkތ�f�9udȐh�և�HG3%��7P��~>�Xe3r��~��cG%������ ��\1��t������%r���Gz�F����,�:�@���  ���R*��Da��@x<��J������Ȩ��V<.��c�NQ�����u.�qψ�C�Z�A���N�t���� #�REJӳ�+O�v?U��R��?SZ��t
:�\�L��@�t=�\���!�֊�.�׿�9�������DEf�'Q��N���uݕ�v���sd��/��{n�C)3+:hA��4w1wp�Ԗ��s�[�} ���/��c�z�=����k�o����I�J��8#?�D�O���Sh��Ю{��m�=���QcB��1L�_�D��?�� ?�P��|,;�u�"v�E@׉�Z`^����R�Ӡ���O�~A^~���R)�QH��     IDAT]4�'�r��!۬�F ���qnQȚ��jmI���m���4rK�z�)Q�}��\HJԕ#�����Νz%2Q*ʦ�Iy�����'�۷H�(4�c#��٣�#� �����ϊM�o�DE�$�C�k����։�+�6���N�%����`GU�U�M��4��N���ū87�`at���v�Bץ�$.~}s�ڽ��k6c��d��!�O�9�fںF@�چR*4��Z��w�)G|@�4��>��L� 	H]��եB��tө�g�����>�qo*���o���o-]�� �Dd�[�1 >����eֻ8J�q�{ 1�<u����2����XtW�\�N� >p��Y���8����m�6���2��a�KG�y�~�)��q1���Q�
����E�}YZ���؂�w����i��fm1�M�Lj38nݶMe��ms(��񐉄e(�e�ޕg_{[�|�UI�����K�P�2��K���\�R*-Y-�1xu$#2�P!�gZJ��;�c=(�e��P��Q��f�<
�"�##y����8&ڶMiadq��T���X�P���#n\�"��.K	҇(��Xf�����B�6WT9O"dn�)&�8PE~w90�W00	�#�{'��B�-u~dԁ��b�Yc 44�@ ?0�
�����ב�{v���A�)o����=}\�-�J[�B ��1נꔩ^`na��h�cȐ�X��:5�\�)	x�N �3>x\�����Am&��$;a�1&F�1 ��D3ʥ@�*(l�mA�x�����vS������ݴ*��'��45#�/kT��3I�0��0����x��L�Qo #vY�:��9�k
�Q�z�{d���j�$3S9d�/]� ���|x��*Dt���v
U 8�%�6mQn13kx��E�2��	t1��$}��ÿ۸LtG�?P�x}�
��� �(�l�{ �sq���g&�,,� ��p������=�d��'�9F�6��ǜ�~ǀ���fl��<�|�5�J�D�Xp��
��c���s��K�6po���v��ß<-��� ���"�P� ��G�=� C��5���M��k�!K���n���!{��.�wmׂ~�u��@��x�R�&�EN.�V�:Q���329Q����W?_.夯��0qk�>A|L�ӵ��y�Z��N��c�X$��-cc��Z���Uԁ$�� �պ� �Qg���c����I﷩�e5N�3��3`�=�4���q�W�3A�+��aG�b��C�ۨ����<tF4����G�(CAv��)SS��i����}r��Y���@�q���#Y ��b�������;]��7���'�t��s����5�+���i
2�$x�F��xo<F}� �[& E��$ ���z ^'��L�&� ��z��{�ߍ�{t>7�����a���7���U8y�F���#���զ7h��r�i���Z� �N��V(����9(�LLT�Fs�}��#G-�Ũ)��E��6А�x����u����?)�^Z�=�LyF�Hf�V�J _�I	ך�G�XuL@IHPhL{�d���rx���sx�����չ3Ò ��Ī��d��sR��� ����{r��%��|Q��
A�����vo-W'�\��t�����B�DAh���ȲZ�	��ЈFB�u���s��"2 �쪬"�1���!4��5`�@)�#
|�+���*�s@�횼��r��S�R�����Ȗ3Y��S��$m��8Ptwŵ�ʣ�V=��b\f6o��ofwI*�̙z��� �Ieтa�!d�9��.��`��b�v[�7�SN7��L���32=;v�
�ѕ��Ϛ"�( �m]li�:��	�BU|*鬀>���-�_�qȬ'�uq\;=p�	
��[I��c�$_~�r�òs�T��Pȩ�$5׮\�&_�>�Pk$P��{Ǝ����m��.�g��GX��v���d^�Qî�8����6ā'΁� }@�gx�Sw=��q�*��$�����y�������<�7^q���&}��	jWî�k��^���l��\���������ˢ���c��9��y�E#&�Ӱ7-�ϥҶ��hؚN#�e�ޒ��͏����覬���r��� �+�BS��*U4 Um�A_չ,��T˲g�vy�dǎ�r��I9y�x�sp�a��H�͖LLVe�̴LOU���;��ˮm[�TD2*�8O�Q�|���k�(.��{�6���D�H>[,�)tYGR�+��3g���s����hh'Vh�+`�i^� Q1[H,�LIB2� ��9l�΁��������G�Kr�yۈ�|v]�����.��53PǙ���-�6k=ئ�)������e����oz-Ƈ�d> ��B��/2����m߾k�ჱ����L���;RJ��<w5����k4� <���7y�_���P0��׌R (�PJ�Q������B׼#.*���pCQ�����E�k�Q���5�)�ػ�9����y�wI��Nz���Q|^yj�-Ί<���Wyg����7���n�����LX'5t5��	 �L2��䧥Z-Kc��n��|���p��Alu
e�8�,?�������J��+I[L�����k� >��R�"�j���DV�h�=��0j���W`�2Zø?�#�	x:l _�67&�f� >l���S��J�:_���*U͔��_��xH���Y�i��R�*�Ӓ/�5��C�,�$��$n`
��Vd����7<2#�c�ќ8�*�Wl$m�`�Tl�RW����B3� ��c�?�P���F�L���i �U�w�|MN��@j�%iw�J���*�^�h#'-��|'�K�<�\kP_p��|ɺ�6��2����v*`V��JgZ�� �-�i�<����:���(��!EW(hd�NOn.,h�)�MkP���6�z����aM.��ڈ��=���.2�a>k�(���a�D�U���' ��ҋ�I�m}�]��x��^d��w�k�3�����i)��JK�M��G����/�����鶛r���r��eYZ�7�k���ogΞ5���+~��*5�{�n9|�pT��G������g5M������69���X�� �e��u���X�~
s=�z~΃�$�gQ�>���Gv�!p�i˓�Ex�I����z���}st
���M\����sѸ��&�y�����}y\DΠÏ# ,�Z�8h�B��{ȗe�֐?���7ߕ~�(�ipk��o�
�=C������R*x��x]�۶m�l.���ѭ����Դ�8qB�{�m]�[7mV ��o7[Z�_�eU�����c������ J���%���;�z��]�/mjP�)�
�u�9�G�7ʴ�;P���s�ɋ/������W�+���`	�}iC"2k6�Wq�������pN����>6tC��kW��=�����a�K�y�Es�o�{6E`�7o��]۷��}w��;dr���V�vgɁ��P./���9���u�λo��ƽ	
�����v.�����k���G#�v]{���mjs����X���`����s�B�
��x�e�'�Rl�	K��-󞜐j0�YI�و�.:s`����� m�9�B�Y[\����|F���('���Ҝ���MMp��ZIc>��ٌun�" �
�Rc>�*�ٲe���?��Q}^7�_�V}Uf��ezbBJ��d2n��d��:�ȋo~ ��K��5�͖D�� R��UY�v5��0��G ��*k��[A<eUE�~܍F
I����0�Ff���' 3`q�P�< <x~
4S}�y�܄
MF�{i/dU�%;�:9����|;@F6��6�K�(b7C5�C^�H�\�>��Ŭ������$�6�U	��L-�@(9�X�P��ݧ0�ˁ�w����~o������Y]]t*E��y!�֬���P�Ϫ?�mvh��E�d�1�ՠ��׼w�^�޸67�9D慙^�O���{B���w[$�	զ�3��sW.kUHgB�feu�_cF�)�%�w�&g� ߳u�6��������Zħ$Nk`��(�{/%-���J9�BY�����%I�˒��H*���do�阬��K�k�J���ȠݔT�%�lO6W�r��ٿ{�f�o߽[�nʩ�ˉ�Ǵ�9:��  <���G���!h�
Yy�	 ��ѭ�
�ˑ�-�E�DI����~��彲���c���}�x��G/h���~���t��൒��9e�Ԋ�p&Ch��N�Q6��������~� ��0*���B^C2p珆��8S��+���{|�T_�F�[��P�w y~��  �a������jk:W�A%���5�c
8ha"����@F��"K�� �A�]�>��!=9|�ٺe�\�rI�tFJ���eؙ+�?�g&�t��&�U�h�ة���j�O�1ٱe�d3�u�!o�lk �I�'�H�c�C�;���؈*]~��w�$�[d����s�=�	 m��ν H 6�#���(d�_� j�4O�ot���Y��tq` �mS[���,���W�_�p�s^�7~�8�os�!� [�Dʶ�[��]Tm�uV0�J��RQH��f��R���Z����w���_��{��?�gS���K�j�/�|�i��_l�;8�L�C���v��^���Q$'X�F��plm�a�k�����8"_+!p��<��'���kG�%�=*�H�sC$_���Hj���q��/��I����@���~��h� r(����bQ���T|V#�ō��2�N�p��OV(�����)�259!���Aա�.�٢��sr���ۧ_��7�eP�TjMG�
Ү�2�ҬKY��(�Gït���� �se4���R��=���K�mso햦����Nn���1�%�%h�O�@�=Li>[�HybF��bh���V]Y�yS�oܐB*�E���@�![�H	��i��r��T�VT]�����;�^�RkU��lU[�fq�x�j�2�A5㮗 $0��PL�Rh�:�v����\��,P;hքyF
���T���!�8d��i��h8�҂Y��kW���и��,s׮Y�#mu!��c�v�Ix�B�y̵���YCk �P���u�V�7p4����~����{����m[w�Ν;�w
�ks��nԐ�\� ���BrM�����luJ��XO��w�B�}��tG6�J�; x섡�M�#C�^Uxz�B3h5�����MUٷk�l���rv w��++Kr���r���ZĊ�Bq����/*�m��`�a�Rէ?�iݲƸr���p-�/�NPെ)F��{�m�ϒ �Yw�0�������}LX<�����y������nB��� ��Ŝ%��1<'��|��c��Q�1[N��{f�JM��`�󟀚�G���/��;�����+���6s̚�.����S@ ��(�W� ;�ۍZj�5���H&_�|uZV�BS?�����:7�k�������J���Q�k ��� ��w�cG�K�/�믿*�.}l`4��s�[���:���G!}�ħ��{Xvn�,�h-�If^d��qsT���a�}{������qS_�`�̾XQ9���^����_7%������'ȹ��]H�h'�ЗYw>&wtmdbJ��ޏ6h3l�'�BFkgp�'��E�:l�\����]�c�r��Q�R�!�@3J �t6w#_(������u����yo�������L�:����߿v�����%u|�)(��CX��ڲ�� �V<��G���Ee,��P�� ���E��D ���7��aol�@�У�-�����@wY/IR�(�]_2r��	��p� �p�\�\h�"�y���3���p2k <w�}��w�!ٹm��{]݉i7�j�P��xPФh�-K;S������:/�lY:�h@��`n��5�	l�#y�Ŗ��)�_�y�z�ď�'7V�'�w0��G����w�R ����@��: �Ne@��Rח����%%m�H^UF�%W,)�VC4��ҵ�r�RQ@QJw�P5S�J~jRJSS��d���V ���(�h�gz�0��`��+ף �G�m@� ?i�� ��!�A�T[�'�L*���������'�YC���~� �s�ϥ� �ՠm����� � ]�y�6�6�x�^3�M*�m� t"%��܆�� (�ڀn9A΃L���^Y���:���{ӳS<�� H���K_���k8�̌I�"��}l_Bb#�k �v�!Z��\uZ�h)�+� S�>$�R࿣��h ��=�{XN*��Z��m���RJw�B�{˴l��J%'J!�--���9��@>R��;w�A6��ɓ���ok�=l���=��c��O(u	�Rwy�]�AyM�M�;�9��'$�*�+ <��]M��L�a����6��^�(u}������6�u�%��N��[�e*mה�������GP�g�~��~�;��?���O���Ee���<�'�y_īv��=8��
%��>$`��2�9��[�Xk�_|����H*[�|uR�eZC�b� �m�ިs 𰝫K�Jլj� �;ݺ���[�s�>yⓟ��7���W_���SY^�ęz���БT���JK���_�ԧ�qPh6o�:0�*���I�֣A�dkm~�i�۱X���3>9;\���0U��{D�^}E�{�e�%�X<���V�Y�*�4d4�:�7w�1��Bg��9aT26�db�����㞒��y��{����A�"$�|���ڌU��Q�(
n3詑�����펽��+��k�䘟u���>�v.���Տ�m"��V�F�+N�V�� ���s���'?��N?0���pP��	��x.~�/?	���&9��8�����r�����1�@�( �A�F ���q`{��N$	(y��T�_����3Q�����h��P�T1Q�H�� ��3�ѧS��c�Sm�{?�Y7�m��nI��Ԫo�h� 0��H?W���5y���Gפ1�J7SR:���#�jH���Fk��Z��5�}��~\`?l�/�q���ܼ���(������ �����Z]��PH��k ��~G<2��.ck�ݓ.�X�*ũ)��lV<�'��jE� �]-�뺫�:%Sf�#@ow���+aG/2�>�c�+吁?z�!Iu����Ϙ
M|�i��Qԙ��*����;m�[wl�9�L7�fjfZ��x�=���۷O�+�K:���<���F��b�:~�Z!���}�s])&'UF �{��!���m8/|@߇��yDN�0��M� ��mz� ?m >]�N�Z�� <>�v6<Gݥ��
dݮ��q�  _���S�u��x��,/,���4V���Wk˺��
��jE����ԩSr��y��ۺUw-`o�@�<8�GN_�.->��B��� ��I��uH;��4�����%g�BpA�H��$�av���/�'y{�k���o���=U�� ��� 3�qp�� \`w=`����|��G��l2��O�Q�|��L>Kr�ն>>�
�%AvbՂ񠈥���V��D^|�M�SwqB$WR�!3� z�P��|mqA�h�T,��P��5�C ��7^��_Ѐ�E���V9¶�{ƷF�������|�ӟ��yH6�N�;� .'	��'h�=�B�k�S��؉Kέa �`6U�8���e�o��]��j+���i�;c \���F����ԃ'��;�p�$��}&�{�͝�����w�����{�ā!h���x���^m%RP����������t����J��w4�g]�N���T��W.lZ�qEe$�x=ċ-)C��xV$A!)4T�I�dԔ��ٙ�-	������A�G�?(�(��H��DZ��nYۜ'i������s$�E���"H6�̸�I���J���\���q�[Y�&KkaI    IDAT�~�۲��}��'�>�
�0��%ٓ|ֺ�j�f�$�BU./5�;{Q9��|E���4�@��5I#8��g����(�ƍ��!�5��
��s�c�_�:[��){�������:� �Z��
���_�qM���
����r��R����Դ�9��tBQ�	�+�?��V)A���+��"�� �,"�;	�#�*'C���阐��������{�t�%�����=yL�92��3�Z�\��ɣpt��-�͆~v�M�^C��sx$��������u  �u��952�q ژ�8����T.,�&e��;΍���o\2f�/�	�\@/ q�`�5��X�ځx4?KW�<�z ��4 �ss�m�}P�M���2�DQ�o��͓%���2��Z?�؆;��.w�u@��߯� ��}���?��x��R��bI���������-r^O��m����b>�`]2��$}���<3ᴝ���0��<��>�`ƛ��Y�]Ҋ�7�/��}"�J��?/��+q>��wJ�u�=���A����8��N���v��� 	���u������������,#�㕁4���r]9���	Yn�TF�! x�q�87�wtW

Y! _�䤪Ji��4��S������K���%��� �����nAR@��Q�D`	�Ub)a)ix�>3�?��9s���u�f�S���e[����p���2}�9��$�G�y1ӮB�\�W��=�.��:� >[a+J���3be�X�1��x���m(:�'����jn�r�ܜ��BN ��ŽDwQ?��q"$lM�.��<�95mmn�TJ��R�EC�V�[NŇ��1 _D��pMn)5`�geHK%h�2�q�z�T2�.BQ�����\#��'H�F��p�A�����ˍ���Q����ܭ��>Waf��N�G���+!cXϣM���-M�0�n�_��uh*�=~��^4�W�����5�w ��{�(�Y-6^���QU������b�K���.����4?+���f�����1�����i�W��8�U�,�g	1W����_8��o������ؐ����3S����>v��~?[�P3�6=~0��=m��Qɲr$�������(r�i �̭��.Q�u����a��,Ex����f�]y�z���"�D����˾Ń����^��X���l�@OY)($+2�����#���"���2���=�"W��3E �g�ԟ!��ס�1��B���5���&�6�s���&�.}8�j$�5��T�϶�/7/r��%��Ԕ���U��b�+7}߭XqM�m�kN����1m2�=�|jj&�SGVԙ����w& ��&�4rK�Nƍ�gK�k��!�QY6"�]F6�a�Q�#�Q=�F�l���oWs5��k�D9�J�T���羞�����7�v=Y8ӟ>�q�o���@(G�6��9������!�����ѓ��x#9���D1x�^�*}�X��R��X}QG��{�	���׺��𣍕-�L��P8��X����f(W��Č$�{����yՓ{����뾋��	�i��c�6H,�I�K�8���QΧ@*��h�D /���O�;Q���#��P�7���ĳ��DP�Ge��H��8=L1x�\ll�E��>�ޭ����ó���a[�F�).h HB�:Ҳ��P����{��E��������Z��E}
?"ڻL��h��}��S=���q��8H��V�aQ͸��^���%��@��;�ꦗ��|����\�P֍"O��U�_J�y�Q��y^P�k$�Z�Q��,�-�̘�Ge>H0c�@�`�
�����z��WC�o٨C�IU�t^��I#'i���؟NCR�9�հf	Bn��}o���5�0���E�zE��w/����@����1�.4]�W�oD�׺f�#��K�� ���d}z���a۽�۳���s��^��B:�ץ�wKTU]?6Q_pSu��̈�t6VYO�G*��bL\�����;h���֓+$6����Yr���_ߨz���=����!��.!�}�F�X��
�&j�a����L�^�l� }3̽�Z��<oF��<��n����[l����^�������2^�ۗ�5���py�o����?��.��B(��a%�z�.���O[q�s�>"�7�$���`-�R�T͡��
V�c K�����)��1��������ZeX�N �ͨ�mȟ�v1�#3��˂A�fg�G��Q橠@�&�aZo�	�*c҅��8V8�����۰)����Cq���g%5�� �J9B��@U���+c[��2�����h
,�z�Jh\�z�&�u"����{cGOD!���Q�8��RAMP��Z�N}<��_v�]��n�JE�hP���'�����Mw���W�5U��8�y0����I�d��4��t���yD6�������U�Ϫ�?�LϤ�G�������f�؋� �M�ߒn���+��=���KFc�-SF�A�Qt���oV�*a���M����Gt�R$m��h�����;�1���!^{s���:Ŵ�Ϻ2����DU5��N�c	�C�Q�@����8:��H�m^�h̦����S�(�S��u�ߎޢ�8%��#�ȾQ�a��X7U�����v�6$k(�a���A�C��Jn����?k���j/-�K�+��u���i����cV��ak�hw ���Xk�V�m>�h��_��x ��/yj�	|�|�h����!�ֿ����fsU=�)���(!WO�F�ez�sW��1��>S�ӻ]���]=���%�*E���~K'�H6�����1Ɨ�=���x�-�GTI]Y���+��R�i��<��&�g'����7QV���S9����������1/JN��O�#�s&��1�'�x$�4��Z��v�bڛi?��g�I�Ә�&���ҫ��"iOCA׮��Vƨ�F�M��ҫ���m��۶t��f�0�����o~��vC��9�i���)�@4��8f8��W����>���09_��l����O5/]6Ց�����L��mH�Y�W�	�$�*���L�� 
;t�Jj�;^",bF��*����)�
���z-,HT���Ó�_�ŏ;�GG�i�E��'	�d\����O,X$9;��\�	������+pP��C_yj��P����jaI�I�4��@1���*nd{k�D4�pM�J�M�Xh'蚼(�Ge�j��9�j)#�K"�(�rU�TW���P	�� d�)�+y�� +]5a�.&�Vb�?�g���\�[�zc}U寠�g�����M"�YCIua�넆��'�7s{x�c�`Q
 %��;�`b �Q��' �?m���nʊ��F]��qw�Uꔀ�,�qu峼��?�7r�F��?��Ni:_�#C�J��)P�|B(��1�&	c�_K(R����P�ϹmW&����db@�N:W����Ӏ+}(*��Ĭ{���Wq��y�ά�	Mow���*ٜ]g��:��哾��
S�׌�Br�	Ϩ[��^�4��F�uFH��/k� �����J�����E�����j�U*�"{.&�V���|��!:v3� 6���B�Nq��/ސ�r�պ��B^���i��������|����^�w���.K�9�&���T��i�f���]���F2��C�hY���i��3;��1Ƅ@��VN��;�T���}�3�`	^����3q��b��~��p3'�K��m[�(ՙ���r�3���(n�s��!P)�韼�IH I�u&�X�2�-ϝ�~6��)²y�(B����KsI�b$i����Ep������%�lS�^�P���X�4���8BR&���������z�f|�`</��(����OT�/d�5  I�0�o	�se���tQ|�N��|��׭{!���W��7["�\UJ�<���	�f��Oa������
�$FL�g1��\�QbҎ�8K7�(R�c�����D���z.k�B�����Ny�c�p�i��<���v��]��������ɨZ�����D�B.z�y�q�lO೵��v'B�>Nv�h��j�]�g�9*V8(��Ԛ�>�f�J(P��� ��3�47��ѡ���ub'�%NA�֌聠r�	�(����bL��a�+!�o㪴ʶbq.J�q����_��E��K������HuH�u�+�"I�!��P��<�k�N��z�^`W7.�C�H���>�%Le"�f-�"9���2U+�$p`�c� �%r�V����k+Z ��޴w�@@o
��'o5Eˍ&-H���e|`gL�B���u����)h�^ut��}�d�ޗP-����_���?�یr��L��z�H��k�F']��\_��Op��󍞠D����*��.# �HFo%� P_f�⒛�������6J�kQ��^[���h	�H� Rk5��蟬hx�;���?��8SUe���OGw��u̳�cB�������m6�6І5��������"oؾ:N�K,f/�c�)����[��_1�^vu�jz���
E���)�N���K-�W��ʕ^�Şɣ�%�p�1�*��p�Vh�m�Z�z%�삒��S�+�s��
��7�g����W����e��c0��w�֯�s���y^���~�@ɫ=Ǩc�\<<�*_w�{��|�����hX��>XT���G�Q�J��7R|�xV�u˹����/!�X��ӡ-���
�z{M���U�Hp�aS��_8���2,ڌ���<���Tֳ��wp"���[L����	�����ׁ�_~8v3�u!��,�z%0����u�S�yhK
����V|����>�+K�>\6U܎{A��G��e7ݓ����l��#gѻ�#��|H����X�k^r6���O�~Nq�Y���j��E��:V��a�
��7ӆ5߅������A!�F��ue��~NQ*�\cGǿ����>��\� ���hv�%iVy!;Ծ�n������,��H�a���Gf���o.�?�J&{�U3n>��y�V_MnoȻi�PT?�hԠ���Z$����f�/J�b)�}�Ϳ���k�u p�����gi1����P%�ec�����%u9J�t���tu`��|�QѬ�⾾i~�ji��X{����x	��*_(���E�X�tU��7�c�|��T��n;���8��Ԭ�ʃ$a�5s�y?Sќ�=�@[��ƌ�l޼�/�{����|��k;���}�AC�q�<MU�o1SJ�c�슞lagѡ8�J��u��ڕ�Sْi��@@y���ԏߙ����v�L᠊Ȫ{ ����������C�&.�����Bc�����)�y�Y`~6���7s>FW@-��?�ǋ��s�શ!�D/y
Gjloi��̋�����~yu�v�%������)h
m�q3���	ڀ�����m�Va㟕0ӯ:ln�[��*j�ť�յ1�
M8�e�1LXy���A�{T9m]�����Q��n��J��8��v��&АN�r�B�B��DA�O{�2�O�H�9�/W/�$K�dDG�2OAR��u�<@z�$;��4P%QBC�y��?~�8�7�f2]�r����o�yhO��&]�G �
��d�͛���5�����72�jU�@s��n���fa��'~�`��_�ɣ
��pd�*T�{�2�Tl����[(��zVm�q1��z�]�%�5�%B;5����<9f/>��}f�+ s���2p�1v�����S3�a�Sky%��d���αN�����O�B �]&�6+D�����@KWaxT���j�ݶp��P�f٦m��;��sYj��(`����:��걧����#<�~oFW���᳚�>��w$�alQ_�jw��S�,�0��7����}$���q˿�1 �|�vl\��㵱r×U�еB��Gp?���{����E�	t��n8�ҿ~;_����Lsߡ�e��m��z�K	�I�m�4t��L�S�چz�QxE����R�>�Q���*9�@,�~�l��JWt�6
q���31^�����8���n�ڇ$��,��[t��[8�����9���u��x�"@��=1�.X���+A�å멪�����6�Z	�ڹ�҉�q`���Y	�s���_�QS@q%Ԉ۳g�MD��,{\2�d��%-q��~���մ�lF �^�g����cd_
w I�F0��W�Հ�����ѡO��~��v��~����"*(��w�]^�v��:�%�N�YY�<��+�+qI�<bt�W�,S�#��|T���a�`��>����oPR<�/������Gwp�@��!��2Xt ���[�J�\�����	��-a��y���`�:�eRmG+�Ji�+�,K��������#/a���w�����	[F����8�)(�~c�v�{Y� M�:+q��$s=D�p��=�Do~�Ve|@�Kd�yƮ��z*���)���"�1Pz^���,<i��q�Ŀ�^�[?�J48��E�p�e�f�Q#�
�kI!`颌���`14�D�f�IӼ���&��Ă��>^��H���==_)�\�	��?�z�2f3j�Kl�g���Wq�/j���/+�b�uYl��#r��O؀�D� )^�_�a[�p��$��#�y�����O����v�^�$�r��+�06����c"��4�Fs��a7w��@�� ׽�)��:��N�kǃ�f��c��H�~չ���Z��?^�Z�m+Z�T�g��n]�ό>���`@s�́q��Nqx�Y�qCO�}Z캍/<+~`+��:���{�	H�Z���+��){�Av�O%�q�o�
Q��㉢�����?�X/���<�-w���i����]�FH��:�'��ǰ�"��G��u
��<�Y EB�*���IW��l�ِS[�C�+>���k1���&�뻓\e�0}���as���֯�������֘�Aj�Lؐ-�:�S?��Vȸ+� ʒ�e��
��#���T9�G=��s�F(�*J�h���>5-f	\�'��cZ�z�dg�J[d
�.g��'�d ��{�΢�X�c_���ݾopN���6J#d�I8-����~�!�O�������P�:5k{%�6�,b�~=���U>	3qŔ69����f{P\����K��a	T��q�b�G�#ƞ�W�0-�v3��c癜��І�U��{o��X��:���|2*��%19�A��;�"٠ZF���Xq��7a�u�?|���$�lLZ��L@�Ӈ�G�C~G�5�����r�p�uN`�Z�f���g�`��]���k�D�^8�Kh��Q�����m_i��&�l�hU �,�G�_Y}�ijO���̉���]3�R��$�`]�?q�z��,n(��d�ޝ�4�x�K*0��v�t3�B��J	;�L0��T�a}���~�r(o�ա5r�"��>u��
?�,^0'.����	7�v��_s��o,���4f�A#�R �~?����/R�:��-rt�:e�:�l��dl�ig���p�-0Ej�lE��/����U?ם�\�n��Ǌ��ozRS/��Q�/e�S�Qdr�(ˬ��t��ĀC_��f���r�Ю�Y�J�B�9��ٿI^��B����_8����l���F0
9�����|t�pL�D)�&ᾖY:ˉ�Y���PQ�gT��U\Xl�])$��m�X�����;�N�&>}*K�i��܀��
�t��Pfc4=5K ��)0	<���g}ES�h�[tV��j�n��~��_e"����������gP�vǛ�Cs&6�G;�Bc���$ɿDɴ��L���%��y:?y��%S@����?�Q���	/x!�9���Pr�?d�W�Kɮ�~g��@�p�ގ��Wj��u��
����8=����U�cN���8�p��w|x��o�>3�LI��q8~}v?�$�/�x��Q��^[=mk�yyy�3{Ek��C�'.�I{Px&1��[t��y�5Є<uqÛp1���4���o`�}��3�F�6:�*�$���tbY�7�5$��,��I�x}T����؛2j����oyN�FI�`m���AFKw��(j�U1�%1I�%&�(��x�'�yR�KyR^Gg8÷���9���Ƭ5,��ޛ�7?�17����������0��t��Z:	W����^�Lt{��M$�^~��_&��>�wӊd��j��S���6ʠ�z[�����;����S�޺�]/c|���7����Sw��,���a��Z����A��a_4"{�W�RN�)��ʳ_T�{��<s{�B"@2ŝ+͢�-�&D�ї\rAu�&�9���C%V�+���C�~�G�,m,c	9��Y�5�2¼��)����a!��GR�Tmm�n�C�(������&��s�P��傞�(H
;�:�4�g5V��̌،�����U��]ifꕙ(v��>G|ܚ:ܹ����J\���3A�gp��
�n��h���H�OP��c0Bc��I��w�V� �g�`���}��[!<XB����+vh�������C��ě#�0O�{ug5�x���^�t��e�|��9�S^��]�;>��x��A#�����a�e����M���X��B͖�t7��8�=��I�m��;��4�&�4CT�jN�>A�baߜ��R�k�NU�?�[$��'F��p��hݱ��b�)|���)�Һ�����w��.�|���J����,�t-Ó�L��c=?�"cai�j!�=ox�P�l��ET�>��^��2-v[q��|�f��{���q�R�s�)�$
��
��+%�m��� ��[D>�xq�{M�C[��ds{�������^1݁�ǵ�ϼ����#��1���K��S�={p��sX�'�*��2�/�s�c>rqȂ���c��k3k�H����v� ���P��,���ϑ����B���-��._=��SR1��w��+��g�Cq�~��Z�J��m
��N=�0ϳ�o�u�}ҨbQΰ0F.�¨8Mb�n�2v��I�w/ H��n�٪9>�m	�s��<�����}�@�����g?�2��Haц  !�Tڣ����Vo��~��艤	)����c*��L��H���pgY�����^���(��f�?���F����w`ڎ;x�M����>(L��>r�#�berG��h5��i�`̔��6��#�xp��侟�f8?<w�é�++Zxz�&� z81���؏<��5�p��W ,�d���� ќތ���{�Y���Q+��M��f;8�9��-m���kMx&����-74��h���p�ѥ��ZlЃw�Ѥ ��u�v�!�2 ����l�V#N�#J����7�7_�Jl����9~|&y�c�XN�>�˒dF0�NS#���o�W-Q;:�M�p1�:��Ң�eh���0A'�;m��ʢduW���eu��O�C.B�� �!��4�6L5:���f`���"�� |S����8�����3b�u򯊮ر��a���D�q�K�cI�@����}�jC��/�B����U �zL㔹M{�>��p\	LK#���Y���{�d��c*�	�p��}������9���d���Y�J�w�B��<�"׫ߵ�[�3�Pos��G�#�n{��Ԅ�oU�`w���H��EûB׎e��W\���[�k��uw����c���N���	���<1�nY63E@�sǁqB�$���c!�I��7��C�(XA�v��X��7z-��`��g׸g-Pd�y"�̴���MD��*�JSEz��Z�����}E.!�IP�h�ֻ|�3����{��/W�a��R`U%��.�Ic���i�rI1��r�|�쓧=�>�:+��nz��C]�0]2�M��<=&Jo5^��oBƱ��`\��-�]�fȇ+ڜ��U#[� �����b�GaN�&-'�vx�T���?�o���a��M��~0�F�1���,v6��u3o�6�������J� XYh-1(����{�a��F�3�v����f��{!i��`��G���4�Gzx��f0#$"d?}��X��� H��?&����_1�#��$ D���X?�|�,Ǩ(LIZ�G>��T'/�/����8�Ľύ���!�Q��}>���S����xj}�oL�L]I~��\��a ���2���B��h:����oÆS��6ߋ�c�-⻤�\Cu�v�~�/5bH��|$T[˕O���Si� ��^���|��H�J�jV��_*���3���_��F��RTsj��n��7�����i�ܲ��6BN8D�cj-jB-S�}�5[�R	i1��_j�簜/�h�-��4�[v� ��l6Ϥ��h�NB�g�=����O�H�~<E���[�4�U��~"��ҙ�	МX�%��!�N�K$�v��#�[פʚ��e������O�2垃��'ɳi�J�rU:T�(�
˃>Y��7���\B7�ʠ��N�M̓�)�-�X����oqx��s�3DP^���AM�<�K�n��8����\E�,�<�;\��^A���~=n
��+��/����%�8�:�r6$,��T���Z�M��M�eo0>P��tLR��*O�����J, fru&�~Z��b�U1���)~�l:����pc!.gHʿ����?���G-VC������]ǃ	�lM�C1��=F��H}C�͒�A��/�U�%B�t�wf��.v� 2��HĻk;�����f���|e�C唲����7��@zJ�{�pfrܔo��}����fd�����H ��G����\���[�J�7��o�&�<���N�J�����'R7>b���0P�f�&�����l�N,�4�s�Odc�Ƒ6��%e�p�<|+��D��R#+�g�r�֤�q3�BK��&猓xlx�tr�!��7�i6'_)�P�b�T"�7��_����r��F�8�h8�� I@�����z�,�!=�M��P`8�)�K	Bl)it�� ���1����֦D����T�����8y��a�v'��gc�\Ј��ʝ�+�^����J�4�r�Q֒i�]ܣ��0w�Zo��{\<~��:�	'h<}�H��<����ɟ�uؖ��9�ϒ���+�k��J���@�ޫW�b�!�.Z�`ڝ�NR2�o��I> ���G�����փ}S����V�9���k[��i�6	\�H���W�CԬD�h9���Ku���[E�}��a�����ҴW������>%���<첟�HC!.����V����0�C۽	�	��D<���iHE\D���Y�okzY�o	��,YlH���i����g��`	����?����1�螷���%vo+k����s�}\c�1/�	5)ѩ���g�_c��c�U�c�83�S���T��[Q�����el��L���Ǔ1�~��|�9F&J��Q i	W�g8.B����ߜ��%�����ñ�>@�D�@MX�V���ҽ���:�6�%:<������z��	B��@�Y���U?ݲEe��U�Vx�_��D����3E.���)=j���{8- �;�1�)�(^��+�~�B�o\�bD�%�	 ´~�0�������n{��"�-��m����q7�� ��B�`<e��X�3�~I�AZ�Od�A��PNj�F��%��D��UNWE��y�u��7q���z�k�X����RM�Nu.��-�N6�RДǄ�(Y@�E�$!Ag��ϯ��:2m�?��4$�0[@Z_��Ae��N���R��:�2��;2��qˑ��^i1+0m»���-M����V�U%1g�d�%�b�E�%1$���|�Ϳ��g/d5K���3�ije��»��7�FvN���Z�a���������V��f�M�Yksr='uLɤ�����sމ��J�(m����ۍ��i����v?Ђ�C�7�jvM�b�k7�~]���05�TWW-Ѫ�H�>{B�>?K�O�Wv��TJ�����=���<?��:�����E�����������5�@1'L:����Zc�Fɻ�����|N9D�mv::Ģ��l����BH-D��ow����Oʟ�pu�b��EȲ�����kOa�gv<�P-{�*e.��gs,cH$Ǫ�"�"c�����A��aZ�XZ��w�:�HY���&}�!I����> ș>h;=~�:�p�V&j�cx����s��A����J��JWlWC��S��)�	�Ð���
e����!Z鏆�j�V#R]����r^s�a���9>���Χ�A
��P�����3��,���� p�+���=Ԫ���}f���N��-~���>��r�5�k̴^�ޭ��7�˔��vV��ׅ�(����}m�ߝ��-�'�;ߌ,s+-C��ǵ4��$�q��ӞAx�-�rȓ��<�����X�NS]��_�Vh�՚����B;1,�c��a�N��z�@3�����eJtLx���z_ޕ�M9[�J��A�*�ELl<��1%ҏ,�<F@`.��˳j���-�/N���?TY�8D����Ha�k57ç�Q���C������_��s�x!i��j�Zc����r�9�8�������z��s�-í|<�w�����;?��Y�|���NRe-��%ԥEs�'5�K�L���%�	֊z������ܬ����S��5�N�/����mɘ��1CC��l�l����ǅ�ב�3�-W�\l�҈.y�o�Dh��_���ţ���(�ڋ���,8��%��K��G�4-��]�%�άҹ��~��z�Ǎv�n�nS�Y^Zdw���;x��d��P���^�qT�d(���թ�*T:��l�4q������	
����D�o*�?$9+@\λ��褙�'��5oN3et�M���ȈK.K���{�'�N�&&G�w�D�o����+��ܔ�\H�lO��*t�B׿[����߶�x�,n����I�5ߌ�觅cN'�,7fߤ�xɱ��w"ZM��H��pmOX��g=��k��{��H(��ퟎn���i��U�z�������&(m�F�\A�V qu�*�|I��_<��O��mt`��7�H�1gڗQ��}�	A�)a�A��u��F�E�f�m/�V��l3T7>.�גԗ���:��s5=�_q ��\��,�g���"�P�b��7W �囏I0�`a���n��<��Fv�?d�uΪ�Y��cl/
T�Ya*�^7��qto�]���(\�%{b�J��
\Ώ�~�Ê�Cѹ�	�>D��o]�ivb݈�]���m�&4���<=�p�++�����,]YS[�q��#��IDιY�� 0v0�ś�^���㮇o��#�0��̡#�>�́vˁv�ދ����z+SO�T�-"��wX��X�V��|��X���ױ~H���nh�m7z���ܕβ�c�Z�A��s,�&�R>�	�0���K�灁�K��J�?9�uI��Y]��vO5�[b`.E�s���0W�MG�s�+0�h�YTW����\I`��{�z竸��@rF����YHƜ�C��l����nsc�_
}�YT�e?���84z;�⏔���V;�O��9�BC�r2iB2c�_��ApBN+.��z�#�b�1��_˱�d���Y�_��P_�L�O��&8xZ�J�>�Ķƛ����._�#Y<�|2��a��~	���,S7|:?���L��0�t0U�^K���������
���H�EJ��~��Y�����B���-�FZR�DHQ��3� ���[wt���)�]G�z�q��RVO�9�b��5�F~jB͗@\uޖ�c<�w!�L$�������(�u�7�ؾ��fgG���O�6�;��2C��{]N�;�̢n�����Qq>��yX�a0��0r�XH����t%�\n;k��C���J�M�q���=cD���t�1��O`�V"�QZ!k���@u[f.���]��z��c`��߼�\��s]Kv�ѭ�����*u���<[��8�U��q9������:�B�N*t4Fc��_�:���I��:[�lڢ�J6gF!?�9���	�ɛ6>��ԠU9����b#�����Բ���@�uܗ[���9
��N���3�Ƃ���E�z�j������b�Ywl�ۡ���	��/��~���.E^MD��m%Z�-��@"x�����/�⺯R�%{��g&�������sR��YM�j��X��.���0��U�)�R��x��T�a,�*��M=�s���/O%��ZWS�����4G��W}�������5�1�]�!�7'7E>hZs��� �@��kƸ� i��G��f|`6l��"�BG��[��:�Y��'�uĤ{MsN�ƿԻ���+�ף�U��������L�祡�
���v����kD6�����-=
'Ā�ҜD����U�4�PW&�p���H0o� -;Nߑ��������Ip�0�ϥ\Kǭ�:7ofH`�cwy��J����#�k�2W�mA�ƫ�x�W�I2u�ԐZ��)��JA���)�j�x�C��#��o�Me����Q��X]�Sc�������/�B��!|Ø�կ�fn(�C)�;��_m�Yd�r��*����Q���_C������;�C �p���r�]��Q�}�v��)��U�+�k�ݑ�����.�25p�zm�Z�N�:kf��^"����T��8sl������d.W��c��	�&a�6��_�g1���k���'���K�?޿��{�9Dථ$�A�fMy?�['6+�V�0��Unu�@"����]<�0qܗ���;��`R��6��t���\q�<�r�&{�5A��#?�����I�T��
��:�Ǩ����Y-�1{|F��Rk��M�"�rGy}��.�M;A�}Jt[�N�(~���?AJǺ�M�~d$�!��m�.���N^���y�S#ʛ`��LR�&���B?6������9O.�_A#���ل6�Ea��@i������;7�q��圪N�*��]���'>����.���b�}���IͶ*���x�I/<���-D���M>G� ����5#%��W���W�t�
�T1f���pZ֊5�%�Z�	��Vd����gc���y��Л�܅����Tڜ�����s�q��~�S}�������5߽��yM�Ǟ�k���L�{�j�B�6�g쁁l��)е�du���� ڵ��辂�We}�?�L���������s�x2<��};%M]OfCm��f)���旪e�@��}8N�)h�G��)c��(�d���h��Jz�N��d�~]d�É�c�j�2�I���
H��h��r�٥��uv� ���m��3K��iC�'�2v���E.�*7��B*=o�w�"Pz2�� ���FE�	2n�&ν��y<�H�8r����x��両�2��0���S��>R��]SHh�[o��G�=S�F �)�l�*M�)���p�V��͑1e�K"ט�%`u�}ktiddd��O�2{`cW��yǜ��ȘQ��l��������~����CM.�$)U��v@sڢ������9G��1^�[
(.��#�t�1_��n.kq����=�|��I��(���έ	�-��x��o85V��Pt�F#�ed�\���;�E�
�����:ܻi:�c����p� �I��`ѧ�V׬�A�����-a�_B(�s�]ʴ�H�c:ڈ���.ai������Ӿm�k�{�{�&��I�檘�j�WG+��#3�"¶l�w��>OW2�[	��O#�N�]>!���>��Q�EOĠkO�K�L'OnQ�;Uu��Ã@���"�T�Q��W����A��aU���kX�Yn��q9�Ly��=��E�h�?Y�{�ޮ��$!�vi���jݮ�x�mCSl�ſ��1�V��r�ӡ�N��8�k��w�N�\(�m��_YO})p������\�^P9�����e�	��k|�r�=���%��q�ڗDt��"�}��0���c���@B���Z8��V(�e�Z��e�z'FQ󑊞>�F9E����rp�p�N�{��M�O3<�4�^7�W��f�!K��'�h9�w�K/q��
N��_T_!��u Bp����q���}юR�9/T�9��;��"���H_�f\��Z�~E��/���tԮ�ON��夳2��ic�̜��4��T�?��A�Z�F( �Gg�İ�|�?�Y��ŵk��%\c��N��2�z�Sdx������M�� 7�	�3�����ILZ�_ⲥ\� &s����|Ya
�la�ͦ�kp��߬Sz�����9"b���ߊ`tlڻ&�a'0Z��1Jۼ�^YEQ~��o�Ty�^'��2����0�2Iplܽ	[���,dz�ϩ>� ��ܮ�I�+9S���S���8��f�.����(��X%�vaJ�6�Hݎ�2)�22����ϑ��2О�c��[����lu!Sһw�i�^R4��¬���J�����@�<C�pwk�Է��F����g�l.�/`��3r��"����Pa)'���� (֬���K4�v�,7l[��N��Hיּ�x����Ftn�6�Ԩ�������!�~�nYX���B���`���ݱg�<��7:�� ���L���.D"=��'8o��(�x,C`{�vT��;�^`!��-}��N��m�=�]��L4��'�/��?v����o�.���]�ڍB}�xOsd�	�r>�$	�����줊����)��|�Qx��˧P��{IO�F[���t�@0J؊LI���"U������G+�N�I�� R@��pQ��<�/�6{H�����~>꼇����5F7"�y=L"d��d��{�Pds�P;��o�d ��r�B~B��%}�9}Z>���:�U5��,�]Q���$3���҈���RI��ߖHhi%���Ĥ�IKiyQ|�α��܈�&�LhHS�st��F�
r��9y��ݽK�gaM`Ȗ�W�wߓ�7�CB��̻�J��G�W��#�>�:~ʵ���ʼ�c=��뚨��^y��'�����H5��RC�)o�����gU�}`vVv��%S�ۤV�I�֐��;r���{gY:m��832r�҂�!d	k��x� ���t�0�eʨ��z�4W�$���	�)��$V ����G?�k��<L�ο�>
��@w�I�3U6�x�V����\�#G����Fy���+ ��rm ��$L��Ɉ�Ak��DC nN!�C'a�Bb ǁ}�5�_�Ϡ�pt]F�ʰu����$4 �*2�=п�*�'��~�^���D�n�q��uI�kr�R���[�����jU��*օ���v�P���ؤ�`����7��'O��І�w#�̮����Pj�Ԩ-��c�����${�f��੩ε#qA
Cr�E8�SvN�� M2)�Ӣ㗍����s<$4��������🡴�l�}��	����FO0�l4��r�۞��Yt}��?
�͗��t�~u�psek��پ��^3Y�E>�1�����lT�{_	'�y�)e���?�����ے/�K"��x�؄`R�S���T���Ңx�"t�O�dP[ڍ����e�r�Ь|����=������_#�DĹXՈ���we}��DUlFiy���O<%�wl��{)Jd�f���� Ub�������wl���F�a���#�d��R�[����Zq�͵�B�u	�܁6=��6_,m�^<f�6�/�n��-�����6�[b`�*� ׺Ͷ�����o�9q����aS ��+�����$�)����� ��&�ɰ"��]0�@�`��p4l�m�ͩ��ߛ���G�V��B�aD7�>��v�����f�#\x���H�s�<X�0Y��j�%�S5�f�,��8��M�!��`�'� ��d:����#�&�yH'Ғ���I(}aU������u�H�z �j >d���pn |�YW /�Xܽk��8|@N�8${��V���իZ��ۅ�?��o��  Ϛ���y���J����;�_Yw��V����\�~S.^�@J�em��g������C��,.�˹�_�K��+��NN���}u�$k��|��ey��KR��%��hi@�4 �v��08��t�)I���v&-�x[˩��Y�sI�y>��Pj-� <<���x o��g� �W�f��	��%�W.}�I�hN�� ^�p�OԎ�������x[�}���y̅���3�u�76��l�&�Z5�4��FKx:�&c��o'��e�q��Hh�ܞ���L=�J(�Z���vb=�g�<��Q�HhV��5�*O�U����}�>��N��yfS�xr�3'��� �Vy��*�h���Ι3���6��e ��O�,��<���v�� �m}����&S�8\7��Ƅ�i�D2+�5�M�u�6I����gu���v+�1�wƋ�]J�/j]d��������W�>��n�l���7�d�`dL�!�����?����-�bkˎu�$��,��a��lCh~�4�-��	�Z�2Y)7���</?|���뎧�
����Z�'�Ӈ�j0��R__S �E�H�5h�NL��k�ɤ5�6�܏=��L��ȫ��J�����f�:��=ѱj;���xA>��9���25^D[��;��`?Z���*�l� ��W��{����c���;�;��� <$
#B�=�0ˈ�#ª��;x�������x oQA�~���/ x�f���4�;�N쯧�v��#G.nl��;���\�o��ʯߞ�1MC���u>�����GKb՚A�M��(0�0� �Pg2(!،�pw��6vraÒ�$b�����}&�n��6��a��[�=�S�n��8Q�;������ݣ%����%�� ��Ծ�0�u���P��̑��~�qu&|�P9���%�j�򙼤0z���7Hbuu�����4(�
�+�+ҩ�$GHk�&��D�Z}]%4���X<p`�<p��سSv�خ� ��VR�����o�W���mu\�Bu*	�&�3٬nF�Gaj]��W]��7L0Zs/��pu}Uڍ���d�����I�6�睷�)�~��-y��Y^Z�lf�Ti4�K���x�h��s ^Z�Mu۲2w����%2
����� 6�g5"u�lM� 8�^tZ����+O�:!��E�W/��?���q�#�
�j��lj0��45Xsx3�:>gs\�R�E��qB�ґnDL����~�/��Q�co �x]�[ �Z�� ���HzdBx |3FR���y	{�.�XK����7e��%���]"Yր"�~`�>-aȆ�*]���D+���gma�?@Ӫ�0&f�Bfv3;.Q����{^���%)0�t_�q�F��'j�wlSQ��{ i��{N��U�>ei��Bj�3V�����Q�g�{�� 8��N�g�� (C % �Ϙ��Y��Mց��Ïe/^mc6l��G�#�B�`��9���i�a�.�˦������V���Mb��R����M���~&��jc*k�� ��� 5�s��m']�qc풲�Ku}M��n��Ԅܿ_V�57�����m*��uc�HK�Rտwm���O>-�:*�\F�QRI��,��M<x�t�**�F�!~��������YGJ��Y�~ ����U2�n0Cz �T�b#uzY�7�"������ɷv
c��.���t~�M  ��h�[��ܹs��vΞ�r�䏼�!����8y����U-���;�7�VWV<�p6z;�!"�'��ah�Fm�YgOM)b|�=?j��ϭh��fh|6� ��38�6v�G	7.f�z�,Rw�G�,|{6vk���򎉄�C\��c0<�<����!��e�߃��n��?��j$��k���qgSId�Roť�H��bIz >��F���8F�Hh�]k�"YJ*�G�Oy��ҍSF�E��30%�2Nʵ5MH�|#;�7�zW.|xY�GSɬj���\�X��h�a4���H�.�� O�s\�'Ǌ�ξۑ\�#�vN�#���Iq��F�����*��⊜{��=�(��$hQki��V̅���t3i��+�	�_�5�<�4��W��p+:�;q$�q��4���k�Jӟ݃��
�_��7�ڕ� �%?'$�=k�W�W�����}t o6�NU���beyؚ͆�c�\H�0m�����Gm��x�F������i�Hh�
�ދ�|D�Z�N�#I�Z��ud�D^���%k��e��-I��Z�����/�;4;�����0�d	��$����rh�`� 
�5�3=��{?3����b���m��$GX�#�,�i���������}�'TS(6	�r�\Xt����ޒcǎiWV�,�9>M� �\�I�v�.cꭞ��O?�d�Us��(`<$��$}l8 �4�;�?cn�>�@H�x�s��y��B��&{�*��/B�~��n��Ǝm>���r]jݺFBx�PU���Ҫ��_]~��kOf�06!��ʘ��5ѪШ�kk��z��|&t\eToJ�>���˦��7��܍뢛�z]��4������е��?g���&�����?:+Y6ݦ$1-����� �'�� ����9D�:�6�[ᗍ��߭ ��$0~ m�8�6�'a�e�!�\9b/}x$��������כ�zRǜ�O�[��[�Hh�kDc�Qy��f�і/�ؿ����9rc����_�p�s���5?w}jeyY���mY��&Y��!���߼N�V;8�D�f�Y|�|�$V3�5�1���w6�����ծ'4�!P������ {�q�F�?j�mn<��n4Q�o�d�&��3�
�h�0򺕌4�ɹ¿��B#l!T�o�<M�
��ԙ'���;8o�J>��b6�o6/m�tQV�m�_)�W��=e��q:�%�Hk��jyM�+�k6��	�Z�=c�+�zY�٩�19r��ܵC�x�C&���w�������&�$�T��N%�O��5p�NcW�ڀ�=�C���&|�&:n�ӕ�Jj�#Ǐ���S�궤Q��z��e��]x_.~xUʥ����SR�4u�����!���������h7�t��Td"�հ�>�h���g���i#'M���H���J�ZE�����|��{�k2{��F��A����&ű��sDHb]Iw�r��>e૫�ȉ*4�O]I_�-��L6�Q@#�l-�߃ >���'�9v�p��I�͘�'cح߱�;�Xrv�≔~#�ak����&���dZ�F-�ׯ�̳���ٖ2�;S��ČvamĒIB������0g���t�}$+w�h���;2Q�riUskl��M+�W 	��N)U $�/�6��@��$�ʤ�9lS���f�(F�5<�|�_����?�Y#';��￯�R��$L9�3�ص���|�����_��JoH~EzC)]l��X�{{��/(+n�t|�&g&���_�Eme��>�/���x�ƅ����Gx�����Kbn����7�a���A�a�-����2����\�]7v3$��~�ya�>�v���r�≔j��ߕ_:+o�w^֫M��2Ҏ��ׇ�Ѹ5c�	���Xm]���\Vr�tn�Nӽz�!�c���'e|� ���\�xA7�1� �RN�ds�:��A�зb��)��'���N?*#��x*�(	���>�h�(�H~�m�6�4�=׆]����ϧ�p��"��~z�	�a����!V�n�Uu�^�s'�O\���B����ɺ�]w�j�����zi�Q+�l��/H,-������{Hm�|!�@��f��l������̾}sC'xqS �����^Z�� xxښG|XEa8����I��@�	��`LXh&��2x\�-�a��V�d����	τlN������3�������m6Bpnǎs�a���qL^ۢ>_ܝۘ���F���j��ie��y���j����{��s���k;�DVʭ��)W4� �N�!$��5�n}mU�Kw��lH�.��1 wJI���z���0��ѱ��Vg�&��hK�^�;w��y՚��Ȼ.0����j����"�8֝$Jg�=Pn�EO���m���r6,Hg�'�|Z����Z�woߑ���ȭw�VmJ*I#��v�S<I� ��ѢJh���h�7�4r��>�+p�M�� ^[�k���\� �Ih֗��K�u���HE|:���� |h76ۀG?gvG�j�U1 �Y9>h���:f�y�y^�Ԃ���Vhd�1��b}3 �N�7[���6�u�ۮc��G�ʯix�z=jU��ۨH�Ӑ�BZ옒ZiYJKwd4W�.�Tx��Ɗ}��g�n�H�!��&�9�o� 
5�ܿI�B@���{/�f���Hq��߸� �EO��Sa
�93h����c�y����ٟi������q�څ�����`{̸p�? ����/��2��F1$^�^�'��m�Z`��5Ϙ��cO21����
��1h`�^}Y������q�X5�2�!��s��� ���0�F<AE�@�W^{G��ZE;x75w��5@3@�*� cIJ�V�Ih
$�⛴ H���:��#Ey���Ŀ���%������D"��Q�� <�I׿sۤ|���ǟ=#�#���kR=1��a>��01�����:��hU��6�)|���}_Iq�l��}����
\�>_����K{�{ e��?:J��碘L���}&��_6 b��{̓��z��w�5ɷ�)߄�GTFc�U�$	�'�h��f���?���8p+������������۷nL�g�㒾|ٜ`w��|�1LQ>\�!+?���M���et���1:��㚁��s����@�V 8�~���o�v3 ?8��wΜ0g�yp�O�����9�����-cC0V�q$�_�}�)��`0�̡-��d}ŊL2��WݸT:1Y��寿�M9�t3EiI�Ee�K�K��p��Q*����ůRt���ڕ� �iiJ�h�ٌ�ڱ]�w�\��[wd���U`��V�����)ݥ	��HZȜ��:�1'I�d_^#�
��i�5H�^~��:H���hQ���-�cy-o	諷�r����pWj�5WJR�CHq:���CKb+�XITL��R]\�1���V:�� <W ܴ�\O�m�3O#'�f�%$����2�*�J�$�N��M;�y�׳��Q_�-�����?*HX�B+�h��1�.�d끹��\�����:�������,|�B�Q�nLHb��ڒȍ(/���ĺEx��\�=���� <HPN�Q��4d*���3��(�(_���d�NnG�U��x��>��d�b>�����>��%c���ƹ����9`G����ѹ�c6��������m���vΘI���	�,HF���EH4�������ɤ xzA ��[5�����������&cx3��Y?��?� ��\��sVn�6~�S:?���Z���7��1�}�Md��۰����A�'��Gэ����z�@n�~�_f��|�Ć��|�,�J���5y������daiM�Ͷ4 �p��Z���sj�S��Z.i�<�?�*ՆTjU�O�9-3Sr�ݷ��H��,�8Ѳ�GAp�֗Z&R��	Ԟ3��3g��3���h^#�l2q��ۏ��Q`X|1�9l��g�V����	�m��5*���w\d�T��x L��]r�y�ά�0ˀ}����Y�]��sS�9��Ԗ���<�pN�L{����*��+��+���n�ad��m��Ȳޟ�6��y�@�Ѫ��?:x�������K�U)�}�2��1ue��-�������lЙg����qM��tӵ���H�Jt'9l2F'gx�[����k�{pL�F�E�.�ނ�H������
���x�͂{V��	|Ϙ1�v[�ۍntm�3c�q,3�F�o ~��]zn�x��$�T;�ƥ��HM�Zkʗ���V��f�"����i鶚RZZ��꒤h O��ڒ����1��$�v��2}]�{�.zӓS=�&�j#ǮW�M��פVY�.aE�}4��G�M���	N�djV9#�ɩ)M¸ds��-Gʮ;>��L��    IDAT��g&d����e�T)��;�=�YB;��%�!�֒���ֵTo����RYBB�W	�V ^�v	5���_�Cg3�q���<2�e$K����_����#@H����E҂^�3 ��^zZG��!����F�9���V�����1a����w8A�SG�G��������=	d�
M�)#��&7>� 	�� x6ljC�2�%rLk6$o�D:&;'��Z/K��&�E�V-����������*;a����N3n H@�]�{��$$���U|B ���5��=��������e��0�a  o<xx��ϚL���D$׈�<�{�1e�����Y���dSC�(�k�grD�G��&�i6ܮ�^��}s= w�3��l$���!"�ԋc�l΅�pM����0�!��E���J����`�ues��5�[g.�\�8jT�C�3��7޺�����>��I暨tP�1�T�YX�ZeM�w��Z�� ��3Oʶ�)y��7��ŋ*�Z�	 ��� �k+��2==-��3��G:)����Z�2�sf׳� Y�-P�xŁ�{��0�fϐk�3�ƣ_�ޞG"՗�f�ƃ�n�����l_b�Ǒ����6\�� y��$�����E�~ܺ��>�~��I���dd/Y�v����(��U�H;�I�٪6Z�?:x��ٶmv~3ۮkh�|����U.�}��[3����2)M��+Ҋ�^P6�+���ǜ����暞/d;��f,��cGuo�������e��hG����g�b���Yl4n��� soG�o<<�V�'��sL�7�?�9�Q4p��o[���&Qj<��9�|0\O=}Zv�ܡ��N�B���)�g���d���H7��j��u��+u�o��d��b�%�ʺTKkҬU$G�2��V�!�dJ��s*�$' x����뛘��∔ʫN��If�.a�ݑF���T+�(&�h��ʬ�+U�*��g�V'��X9mkFr��l��!��cR]��Zi]j���sy�Ϗ��ɞ}��+M��{G��<�3+�;��.ڮ���]� �0R���Q�А�
�I�������SPo�&y3 ��Q[yk�]��ʬ}T �kYMP�'E�so#|'�9��?~☬ܹ� �����V�:�A �K� �˭�C?���:�����b�25�#����F�6u&����pa�y@?l�C4X�u�� ��K:/ٱ)�аn�<c�Y'VWAR�܀ޭ�&vǻuI�[�O�e4ёm�9�Ҭ��`uyIaQ2�����d߁��,cg(f �x��S;���fƗϙ��I^�Q@�/���Ȉ�>��6��Opϱ��,06}: 6��g�Qƚ��ءl���� ��D��X#'� ��܀7���.!{1�����:�VK��JGvN;.�d��׬�u����Xp��l+�������qW�z�>�<����5�&�M����Z�s��;�E;����3�޾gu��='gϽ�c�[��Jh����֪4tBբ�rwQ�Ւ�"��$�C�~j!�{ltDN�~B��'䝷���K���^:D#I{��p�a���fe���rdv��9��<��	��w |8��]]��!��w�<C�A����C�M*g��~��*�������~лXO�A/��(�d�� �"���� �N+�R�ׄr{�~.ܤ���<����q���"��ZNW����� ������J����ٓG������̶�s�� ���]��Ji�?_�;� o�x��w�ޒ6Ve!��x@�(,3B�g���_��I��lR�A���A'm�$��[x[86���̶:�Fǰk�j�l����1���C�����2�B o�a���`w�Ág{��G�GW�+{�O���8�+� X� /��ԩKɭՒ|��oɭ�Ty-��r�*����kuIt�!O���]gD(��ɦ��lJ�Y��B�a������q��Z���^P�19T@�Q�M #�I�]}�t2.���C�g%�L������Meh��H:���S;ed|LVW�diyUZm��^�醆v��JI�޽-UmPԖbqTr�V-��O�XU�r��V# �SV걖Jw��ݺ-��š �$�D:=��J���� >��Ҷvb����aY��.������+����O΃��'	,�*U;ע���$\��{}�� ��4~��r��U�
����p�l�~9��5���9��H�H����~!��SF OI:������F�IO4�lahW�#֩I�ӖB�#�XK&�)�T+��6��Xxg=Y��3kf���@ ې9��VN�{�����\�^�'��d{#��7�j6��
:��������ZB���"C�+�MMu���L���uٸ��O"�ub����6� �V��I� �O|�*�A~h���4�>���=��8{�:�bבQ��EO��='�O�͆�f��ml��諛�}YS8�~�d�lÍ��WH���'�ot=�u���DJ;�"�A���������@���v�D6�i4 ߨ��Ӎ�s5[]Mb���O���� ����R-)y�Lt����m��u��@�Lˑ���ӧ�GO��I�'wD#�!���D���; o��aXǍu���׭{ oe4{��3�ʒw:����ka}�ie�g��Ppk3ۓ��!�����c�H��;M���VwQ�+�>6/q�}��98.;�dH_� ���س���u��T��K���ߏ��U۟�ܮ�q=�*4��W�}�7�,�Z��f��>|��ݱ����� �����RZ�����m$�����J"E�1���:x���kȌ��@L�aa�y�|#a;R�,f��4<��`x���ǰ�نwo���6 kF+4=;~��{N5H������ͰMR���p1�8�aalKp��������X�1���[����E�����ʎ��%�v2	�r�eb�JI$�%	�u�ri����++զ�5�Ri���+�i4l&�1��p <�$〕xW|7�yi4k�j�]�lNk�îÐ�Ly=�L(XZB�^�h��|.%�����q��ۀ���*e�(��qZ{F6��\!��%���ZY��ݻdffJe	���v#,�nvdeyMr�M	��|}� �����Z�ƃC76��8p�=�S���1�&��'�
�:|Po]�W�=�=w]g�֊>�Ih��f ^���a��µ9����܏����}��S�^����R�Wq���`�8P��DdD��{;�1�T��<I����O#'*m��7^�`x ߿_z�U�fa#iQ ?UHK�Q�\Rdb�(��e�sm��CW��<�أ
�э��  ���];v���'�k���9W_��쓑D�X�7��kq��k�{6�x�{�m��*�h�5�k_�����1�M62��׆=A�XF;��$/�ms�50&.\�?��?�gkO�m��M�l�*����XTl��M�����ʯ���zx��������o�PD6@����G#�O3�e`w^.f�-��|�=��Q�٬;\�u+�H1�������J �	(�̩�=�G�r ZZ��Y��� ?��UhZ��"��x << �ʇ�����RI�+n@�V�U+��29>*ۦ�������3��ч�l*�D�i�K(�e�)I(�&��57f��sv�e����G���f��(����ʳ�H�I4?w�]
�c�QX>_�EȘw�LV�<�A��2y}��1���F�{�\%����duVV�U�Ɖ�kqh �Kص�p��9�������g��#v�[�g�Ϣ��5s94���g=���Q��Z����<x����s瑻���}� <%����N?1d�et�X�	7�Ü[`�S��C_���"��5����Aw,�����p89�P_��x*���ms��6z(��m3`�،y����.����%�v���O�G_�>�x�x���4#�9�7�s~fp����K���7��`����2�mZRɴJfr�V`7���SK���$U�ڜ�ݷ�#�-������MM6��!�VSlZ0�$�������R^-�2��{vj���%e1��4�m:C�7�`zrzJ�0׮\��Ҋ2)�4E�l*�s�8ր�du��h�OL՜����M���f ��gef�6Mꃍ�T�V#y��uy����դrMF��g�it�Z�x+ _�u[�K�^�Y��I'���m;DriJB�����P�s�͊�TF�z����z�>Hb�q xx�+����/< wo^�W^��ܽ5'M��= �P� ���^M�sz��������:�����m4;��2I|Xb������gP��q�<���&t=�8�jo|n�6�2Ge�b,Bz�=	M3N�)M��TB��F$4��t��Q���cm�Ȥ��h�t1'�nK򙤌r���(��z/y���	�>53�cD*����:��B[h �=ٛ�l{h7Co��>6�L��{֕�t�gϞU������>&����u[�2��6`_�G����,#[Ao�Z7�o�(>�T��ŋ�/}I�
Џ���Je7+?�}۽0>��Ձg|�?�8\��p��Q'[���لQ��yhޑ��&����fBI��>��5 �4�۞	�>tG&mT�
!�?!�+��koɛ����ں4aM�+�~'V߁Z��F[c�VW�U�Y̦����w���^�*���SgdzjL�}�M��!Uh���b�dw&U��S��ꮝ3r��a�ĳ����$�I��p�5R��QO�Mg����C���~�� ���H�m� ���w�9�2����b���:��p��]M8��k,E�RZ�4����M�jdz$�J�eT��vr/K��a6�܁��G�77V-����̍�P��.�n�\�G��%�1]?��w��yA\ �H�+�.�:��:z���������������me�q����� ���Y�ob�n ��h���v��`� 4P��C�0��+�v���l��4#�u[-ݐy�l<z�?�(�o���ez`H��T���	lt���E'���6Wf`m�X�0<����g䳶{�O�R@.K�s	Y�(�Î�AsN��N:1�ezrB�ټ�yɧ2��� 7��J"[��JC^x����ڛrg�$�vG�Նc���*Ih��f�Nx��q���5IfS�ؓ�O<&�B^�$�LHB���P6�P��o��ryM��w	_+R(ettD����E�vP/�"q����Vȏh���j��.��n�c#�2;;�L��?�ǘ�s��ju����������K�0*�TN��$W�4x	���fJ`�5��^�����Y^�b��d�X���L�H'����v\��&Q��Bg��19����E�FV�+�ȩ�|ҡ�����ڒ���Iǵ��]�e������?��;�5�Q'/�M��D�⮑�	�W#��[�4�.��K���Ӝ�%msl6`:f-dSԘv��u}Q����9�����X:�L�ڗ�ԯ>hZ-�e��c6�����E&'�u���B|橅�Ѽ����fKjm�D� ��i���и�prATjD8�{��gG�����4;\L�y��d�-�NS��2�KJ�Ӗ��iժr��5Y][v�8��� �S��o�1����?ԵǸ����v��s^��
�׬!6A����c�! �5#X�ӄqO4��c!@���~���9�ɘv�����.�W&��(`�#�!�i�mB�w�;@���EgV|d�� �Gy���]��P2kR��_~YEao���k�/�j~����#$p̧��C_�S>h4d$W8����^_��m������o�~��r��zU�v7�?��\�yK^}���%Y\��v��|�����O�0���2�VS}��2�]4�-Y�� �#r���$����Ņ�����u���b^ڭ��!f��V�{ ����ZN9(�\Z���.~���$g[�?�WY�Oͤ*c�7�#=m<��E�|�Ԏg�l� �񃯾��<���r��e�{��]�3�ΏRO^s�W1�'L�s�FK���{B��}0���ąF�k�:"��lN�+�-򬩿?2ZT��4r߯���S�/[ic@��3Mv�P���J�u!���U���������0P,��*�F����{�ݵk!���������~gmm�3�KK= ����%4\t�P�g�_ o������C�m��Nf�h�`3�(����K�a�pRFG)<oo7�ˌ�@B��w�^c�B���H�ABh�zĒ"�zh��s=�WP�(z��a�6�>cw���¿1�0~8w����ƨ���9 ލ�K�"َ�ò��-�e������~)����ؘ.��bA�4F��(E�YY\�H~rF�����|U޿|UV�u�����԰"F��0��m1�� �-If�r��Q9yꄖ\��!E�rZlyyIH�q㚂WB�VN����ڸ����9v���	L�/��e�2u�h^9�H~T�٬:�G��J'en�|��ߐ�w�dj�6�^�*�N*/�fW�@�(�η�p >9:"͔�#ټt�U)��K��&�8�\��LV���I��|W#�Ok���<� O�8� x]�A#�A��� �i����2����[�.�/�@�ޙ�{�T�ʖQ��i�T<�t��溴S#ͯ�)��I�3n�K�|�G[K�l���pi�]������ ���Xu۸���v �?�F/�/+6����ܹ���*R��kuI��l��=�|*џFK����Ƨ��)�FNie�\��a �_9�=P�L�"�amiɻt�#�NCv�e�HAR��Lr��������� ���(܉'d�����]W�Z� �1&"���TWO�3d�qI}6�D&$�B����xt����M#z^݁��t�2���6?�9Ip��g#�v�7�Ŝ2���\����uN�ٟ���ꕋd|L"�g?��3��o��6;�V�����?�k@�C[�5�/��k6v�l�c����ݻ�g}r�6�f�6_}�晁�pc0�υ�w,�=A�1M�DZnܾ+��;��{���4;1mX�z�^sX�M�/��C+���:c��s�69&�wNK��"�JI�F-������
p�-eޕ\�BM<!۷M��ٽ��g����{d���~U[��8�������*,!�}f9�����@3S����{4�b��ɦ��+���
I�S���,��WT�3����_��U+��,^?�C�Sq$Gɾ\7nD���k��u/��X�N��$%�ɨ���܃j���AI�]t ��Kk�Y9��$��PI���t�l]�_0�\�� ᙈfG�Z��ֻ��{��#�ۏ�??�ޕk����
��xW���:i��@uo�G�Q��H��-���Ʒ"6��!3$᱇��~#��wB�n����cj0�!#��f'4z!�cǱߡaw�5Xo������]��ǋ>�����x3�Lr�U~�]�n�C�I��¯� ��ڝ�ю��xo�����<��Iu^�LZ2����D�Y���9BB���c��{���_�z�%e�G��>�B�;��s9��Ձ�f��Ԙਜ>��v=m��K�Z����<��VZ��ξ!7o^�\>#�֮������������>�γ=��o��  ��x�0�0��ԧ�T�5u�8��'���<��\�q]�ߘ�l~D�]�%o�}N*ն�٬#g�A��o�4�@��	x�E�W�1���'�O�Y�c�9��X���%6�|6�|4 ��I*$E5���;7�(��s��t�M�8�t&9 ����,�kc�a�p�jU���27lPaz4���I�D�i�#���c1ϊq��b�p>�O����aV��ue����D�SY|�r�l��v���5I��*�*�5ۍ�2�$�)��I_m�5���<e$�c�
������?L���w�ӪI�ݒL�!�Oʡ�ۅ���\F��ܞ�Ӽ�F�տ��s��!ٿoV�{�"�o���j.0���D�#    IDATu���Vj9aZ.R3$�1b&�fo�f�w\D�uO���1����ɔ$V�o�[l��-P��": �?��?T  ����h]E�{ ������� �����l/Q��m�1���|���VB�)߁�g����]���zL6<c�+�!���5lR|#?|�|HT�dUh�s�!��3^�̱�,��G⣸��>�߃�Z��5��h����Wߖ��'K�t�l�)e�*��|����RUH��CL5Y��W�	��H.-�#y�$:r`��ݿW#cK�����(��]I`�A�I"s�$)3��
�?��9�o��)UJX�"�%fc�wlq��I�/Y�G�{�v����Y�6�M6K��W�]S�Ggi��XR}�a�0�jO�^��D�#	,r��V-����&�mu�t"�ֳ��k�46V>��*v�l-Q���a[3���6f�ɑP'��zP8�skYb淖��L	���!Hx� �u|�V_iJ��?p��ۻwi+4�	���sW�}nuu��/-,l__+i�&�>�4����d��|�d��m"� :���pj6w�v��&b+ ?���4�dƞ�0�fT��1Cz��Yxm�y�ކm��r���|��h+��^����q������k�.� ��e�[�>>�b��A�>&�J̇��|=^ǂ��2|�i�����º�`�)mr�����dz�.�ygQ��+_����$2y�5��$�5Ьad�i�x <���mB��#v��a����N�&�s7�ΝyvD�W���ݐ��m8C�����W���^z�'C#i  U@��ޞ���tK�u�{ێ=*�=��r��*�!n�8u\ل��U]���\�7�~O���eu�*c�S�L�V�!�O��*�GBC+ZB <�0 ��$75�c�	NBC$���1��F��:���)LU8g�QҀ�r��hϏ�c4����Cr��Y�uM�����uS7_iΓ��x�u�v\�S�V�219�rJk�x�w���%&�-�s�#����c�����-..+�w6DdzzJ���V�(�V𺰰��Д�������*~��Fdbb\��`.p�F���=lFom�;*}���,]S�nI�kU�� eJ���w���'��Ih���eI��w��n �y�*@1�i͊߿K=~Hu�l��-��q]�*�W���&{���u��!-W����k
�q�m8vC���$cc��%��5e�ͦE%���͎���ƃ����J��3e�Pz�fH8~d0���8��@��=�k���+����E�+��@�%>��k�i�'��Ҵ�֓�8���[�N:|��s�l&I�EO�(����X���i7����5O2B����_�X��"��u�3���F�J[�����c�wm����G|�}/�#����L��⪼����ƹ�VkI<��N�-%\Y��K�t��\�V�CC�<�fK�k@�T�#����'˩G4�{��6p_��.�9GO;7W�\��Ԅ9|@�};�I&�X����%�-�����}�ݛ�O�8��I�[�So���-�}�ޖVV���ڹ��5����e��HdP	���0�<'[���`�U�T�Q<��;y!�
2}����1�\\tC�k�Uγ��k���A���޹lB.iе:���mj�������1�5i�?���K�'\���j���R3�wGO���+a�޳������'�]����ʿXZ\�V^]S�&�Q�MBcF!�Q�����Q i������-��5��d����w8�	���]�0�oF�~o��.���� �鏢�t��خ;�?�I/I�>:�!����F�|}k o�O�P>De	��7>X�ò�9�254FҰ�[p�n �<%��t��Y�h��V[`����/�"��oIC@�"L2�M��
�$~'N��n�y��	��dt� ��Z����"�ZEA>����ܚWfe�̔?~TƘ�?�My��7��.p���6��A ��wjQ���S'�ӟ�I��,,���7ސ����XQ�_�ה�D_9==#�DF�.�ȍ����IH.?��}(z�a ��zvt��������zYrT.��Xc��j����P �O���Dh�qƽ ~p^�l���\k�QS �Љ#���Crw�����kR+�kn�6LI%$��8.����:�%��pjzB��$��I��R�֔�[74BBd�b�"��t�r�];��R���s����{�� �gqq�����`��0���*�7�s��^WL�إ�_l2@J�.��Շ�I�\�۷�:�>�V ��܈Jh��4%���I�
��Q�|�N2L����*����
�8�O�~��==*ӣ#�I�\�zE>����P�p�۷Gu�;w��w@���w�Ͷ��{Q�#0c<G�Ԥ=
�n���6��6(����X���H�п� [g�;�Ĝ`~���#sB�kcCbv�`%8��5d :���<36�� 6����C�H�.�+���3�WnBl��kl�8�φ��$��.�H��9����m`T��KRZ�Ebm|C���g� ��ڸ�߲g���o��Z��������l���Z��dZ�������Ⓖ��W�wߗ�:H䦄�o�cI�A�Re�q&*=n�dP���FS�keʥ����O>"O<��d�1�v�Vb��<wX�V�#�c#:�a\�ϟ:~D>���e����1������]�@%��z;0�8��G�,�'�������A�W[��*�F $�t��u��#Z--��ڨT\��2�Y�p��H�Ji�G$�:ߙ�ae;���|ẙsƞ���+i�r�^���d���q7wy�Z�����
�tz�$m�*qH���H���=�v��}�4��:���� ��6%<�xZ�9�f�n'��g�<�MMM�$�M~6e��_��ۥ�����4MF4Όp��V���c�p�e�%��a >
FÉNH���Cc��-��'��q�Ǥ���5�����]$�vM�����i�� >z��ۘ���i=͉�;v���;��yQ�W�0�����'fA��Z ?'��~R&''��໌'�w���߻����|��/�͹)�MH�L2j�F�>���	)�Ǎ�*����Rac١W�ݤ�c]�uI����M�c
��b����b>�@��?F��.���B�Q���^$º��T���*�<yJF�'��Ҫ\�zM�� (C�}��u�t� ����$�-jV�ԓC��>U�Kh � x�Є ���j�sy���I
�'UG�n�x�F|�<!D�,έA	M�#���:��'a���x$4�<� ���+7�_�f��%P=i��.��d�ސ�H����y�^]W�F�v��ɂ�����=� �gb�V j��JY9eYc�j*�����,--���`L �c���}g��Jk�w9'ue���ʊ�(�H���P,��8P�œ��jI�l��I4[Z�&�S �J�Fwc:'��UF�4��S����b;-�ڳ^R=�͞Ic�6*�lU��c���N��IrZr2Q,��7T;;w�>+6;v��9-�Sډ���� ��aS�xo߱�g{]�՚���\�����ls�W��Ι��}[瓎)7�h��20餟����MDK�+�b���q-\'�Q�P��C��JC+N!%�ix3%(3y��9�ɟ�I���ƀϲ� �G�2�d6T��XJ����_��>G4����O���Bʔ�&C�������U��簹�\����8G`�� ���o�������&�)	q��։�:1zm��l@����Ҳ|������o��Nk�;�]��Uu����L{i�5��25�WdfbTN>(�x��ݵ].~xN^���qM����CR��U;=�\��1��9>��S㣒��(&��v��P��# �{q�{%�!~���d�
:���*D
���8?��R*���#��h���E����V��蜯�n)Y�S7�u�X����<�2`�m����г�],Le��t��S�L�{W��R>�o����j؇k�=xX{�P��LA��v��V�s��L���>�333%��~o
�/\��[��+�]ZZ�Y/�� <���o�_AB�V'���p"c:l���Ә;��Ö4��h�h��ЀD�� ���DD}t�oL���IM��;�co�I��8#풣�a���:7����h8.�7�:G���Đh�������Ws$��=X�S'�ˣ�<�P��n�{�`�de�Z��o�+������m�vS��4Gȋ�;�D������k�fK�c��%��TC�|�Ɂ�`����N%�JiM=��w\��p!U눉
/|��T�+��q�G�+!���踆u�զ�'�ĵC�WMvRKM6�I�I��H�e���V} ���O��$V�[ۨ��|2��0 �J�t�lw%s�(�sJ��A�LN&��d���G�1�t5�T� ��|O|���P4ZN �� H9 �sPeT�kR
�FG]�AK�:��ڊ�2)��\�T�1��ҥ+�v�ޫ���������T�r���=��p@ #�Y���\�$�L\$Q�H���j�U�0 dk��7��60��Γ?Ak�ё:s��dn\5��dN|7�Q ��>�w�' �V8t8�������u�ֺ�%��:$O?��&���2V�jK��s����9'[�fe|lL�����m�����뎁g�q�p��c�-�e��d�3�h�=$_�6��3@�[�N�<_����vf��J��N=u6������y3�什}��Є	��3?�3=�I�4PG���/|A7���K��I��6)�t��\0]�]s���h�u���O=��֭G*�u�xY-�g�Ÿ���τ�������ưo�����������fJuԾ��E.�g�˞��"~� ��"��Jf

���+�΅e�Օ�V���0 o��Gu�TI;��3�-+�(�ɡ{則�O�ZyE�x�e����^)�%��q��e�)DYGF���]�#y��Q���?#�#�u��g���Q�0�?d5a��7��$���g�C_���͔(��cɬ��@r��T�sS�SUm]���ZXr  O��d���c��V�u!`�ښ�����7��!��RiU�f�f��R��:���L"/��4�z%��z�7~Ig�c�nΧ%�I�]�ݻ_N�<&���jwU{�;���A�hӾ���[������~d ����[\\���ˋ3嵒t�Y�K����~��!@×f(C �<��'�! �sD����=
�m�G�}?z��sQ���x���ޗ-������3�vMî%
���3|>V.-d�lB��0v(4�����T�vI�t�ٴ<�Ǔ�a�`:y��P��yM�,�W����o��y�swIr�Q��FGҩ�f���`Q��=C�Zm�,�:;�$'�LԔ;�nK�A��Q9)��hV�/�h������g�F�?q�l�Z��B��1w�ȤK�(�RkS1�5����Ah�I�9�pR�[�I�'ɠ�*��(H��+#ْ���ƕ�o�@PF�R���o$S�Q |T�s��^Џ ���|�I�� �$40� x$4��v;�=1�Τ�NB�kO��8c����P�X�*<8��zY�!�4��@��9�}�N<s7]�(�2s ��%��$/�#x ���eǨ�f���Q� �/-���h򩨃�����c�d������ҍ���͍�q������m�[�XJ��;1Ie� |'�S�$=�7eT�U��uh�gN�#��"c-dN]y��c�����HFF3�̦�`[*�%�Ь�P;����w�~{@R#qk @��vo�h����yF*��e:��0{c�7� �����`�aV���� ^�O^^b����� ��k���ی3��@ �!��ϱx/��Q����ɟ�����9y�����L����$1O�J�tDWE��1A.�K/�(��_�(���'��g�a�u��Ȃ�� 2l����[^��� 0��M�+��0��cN=yg`�χ��pf~�����`�=�7���߸�(���
�kݸ��l���k�/	�5G�Uy���M���V�ER";*g�xDfƊ��;g��J�Y�5ܪ�˔�絸���6�Ϻ�9"��?|���BN�Ӑ42���x� �#b�~}k ?���{��w �i��oR{�q�{y�I�n�ݒ������p��d}���r-���q��b����~����I͜ดmf�a�{�[Nj�qvl����:�h+��v����c�e��F��k53_G�$V4��Nw.�����=�g�;ַ�қ'�^������Ϯ,-O�`��4�	Ͱ�7�� r�gF2x���:�fC6������h��
DG�y��XQ�:���?l���4`���������akh(�xv��H�`>\�î!�B�g�����m��B7�f��/ǜ޾M�=,O<�t��#�&�����o}O�oߕL�oiwb���2)�}���TV�u��6 �'�t���;�t�ӨIL�������l�j&�E\N��AC^^_�D#����<ԉ���y����ǝ�F:��+�2�U~Ć��#qI{
�S�`6[��͎�a�ےˎH&G}l6.��l749����G\ |;�Q�Y*IeaQ%4�XB(�H)?�@��Haf�tH�� x:�R��$4�>��`���o��#���$V�`� �?,�?�Uh^��w���i�H��L&E��$��~�P3��l�Q�\kTU����$c�R,��c�)��_�|U��W�!�����"h)F�s.X5�`i����;
���?��T����B�y�|v�֭���3���/�d�=�|��5&l�̦���G@X�8�@we�,5*c��hv��H�>������bii���M�ɘ)��:�-�\��%��YgӺ:לR]��d�����e��GOV~�I�$��kwu#��� ˋKJ&��2�z����ߞӱS[�v�<�������.�:6[=}S�<�Jd��!J~h�M ,� ��r�,�OL���� ���7���r��0�<{����0�������QMiϞ{��������'_��W����ͮ���Z ��X�+��h���Oʎ��� �t!֑F�%��K�տ��ʓ��Cޅ�f���q��L*�E�O?��~xV���&���O�$��p�Ihx6!��'�Ο������@6����n�;- ��\�~S5��\�(k5g���U[	7Z����T��F7����e��gN�у�������߼���ؚN�+��ޑz����5�$�TI�����'{H>���_�lFZ��>� �C�o}N��pD�� v�,��C�>��Lԗٺg݅k����� ~����#��Y���I+��Zsj����j��k�y����@NM�z:thV��Y���f�� {�=����c��؃7���&��q�����]��"Q�b�U-/��G�I�+�k�@��V;�с��7���f�~���=_��v��e��l���t�7V��}yyy�Li`��>�H(�	'��m���������F�j��7�E4h�/�^�V 5��=<���~ޘ��D8��sD�Fǹ�O��gtA�����7��fKX�g�a���Y�n�b�k�+�Vi�<yJk��G��4���W^���='W�^�X"�ґD"��mt�q�aU1�k����m�M*-QN��� �I'Y�yIǻ��J8lq�&$� c�ڛh��3�ɱ�ZU$�,���4;���f��G�l�I#��Uo�S�$��<XƁ^��&$�lQ�Wפ\�I"�Q�D�B@8F�J]xj��S�#��J=M"$�rI�KҮ8 �[<�.,�& ޚ9} �s�W�ꯏA	MX�A?o��
y;tb����Q�/�[2w���#%Q�%��;
�~�v����欕WeiyA*�v)ur4�7o��
34O"^��T��#��MLL�f}�U��IL� �;��%?�r໨�G�"1ΙdsiM���ӚOi�n�=bRZ[��rY�Ъ*+�MZ?��    IDAT͎LHjd\j���ci�g��^��_��9u<hEb9`�zU~�I�u�nTd$����ӏ=(;�ǵ�S6��f5l��V������s���{�.��p�W.]�jP�*J������4�^�b��u��c\C&=7�=s��Ã��N;[�7�^m�G}��{������x���&��� '�����c�Y��i�D�G^�9 �׵nI�ܧ�Ɍ����ǦZ�=>o@�9	���o~��a��c쾲3����^��b���UqQ$����`���`�`� Y�uf�$ƌ3� 	����I��t<���n��V��VK�DQ�Hq���}y�|߹�[?�W%�$ �X��r����s��~�@%����,��s-�����L8�xb,�pY���X�Trl?}|ǰ�Oe�x�P@����Z��1+��T�HD��ټ'&���݇���}(��<�B-$��@� �:�<Y �d�JSbc�f]*�T�y����ǧJyk]�z�O$��"G���#���H��PvŬ}}���˯����~Ib�d1��ʌ�<�$�Qb��X������+�t���0��,`�mLX���������,#�ؗ����mjA�����\�������3�?�F�Τ\�"��4<�����⩪V���+T�����`��������<��ğ��`g������~�5�e��j�Ο{E��<5Vq���:��f�+�����_9qvߟ�B�K{���9���������6Tp�s�9u����b��ͼj�vC @8.����E5:��/zm>���{��D�O�{E�}Pt�������� �L_a��=ǥ�3��lڒLf̐O��A�ƌ�fK[��Fd����.�d"�qF�N�<)�N�$!���Ɩ|r�S������B�{�G52�4:L(��h<x� D�s��A �2����N9R��&EOZ�O�ɱ���ȩ��jDPDZ,l���"�`��[�&����:K2��>���s�[\|�oS�g�=_*�F�����ar�s�9����'Si)�ECJ<"�>�+w�< (���x�i��+0M�&��#�G��PL9� �5��ZxR���X\2�í<65���� ��
���������7z��p� �����qYx�X�����Hm�X����
`*4*#��!��"�eu�̋����T�I�����E�lFi0�p�F�M󠷷�@�D|efih��Qp�M��a �1ˈ��V ��T�!�1��-�=Y<;<���4`�F�ҁ2���n�ˎ������^V(פ�H*7 �ܠ��1)���gZ �	+�1���W[P��a�2֗Rhp���K�����>v��eb8p �"����*�P�)W���G��%��e��gO���ʲ]�@���	9�r4�r��44Bn��l��%��#�fKq���3q{?����_���\x< 
 �� \��ߦ����L�]��b.d#����!�5�%A���q\Z�1�%h1 ��׉�`.C�͛pL|uu��!z0V�A��p^������~s�p�P�o��e:��>�K��p��=��l;�49P�������,2����r� ���ȓ��*�1D�w�F�j4�F���VY�H�T�}�i���Y�:x@�֖�/��7e��A941N|��z#O  �u���*g��/_�(���*�I;C�l��N׸�6����Z'�Ύ�A\Ғ����� _����V�gPc���.Hw}������Sq�T���lV,�$�A��?�8�k����5�	Ń!R]@i=�����e����ݑ�7>��_�|��vN�g��}<7$�q<�@q|��3�ss<Th������ʤST�K%��c�*(�F�wd�Z������#�|���?�BZ�˫+��������w�������b>���@�S'���f�!w�A ��� �k�A���8PA�F��El���DSH{؎I�}81�ɽ�$��� ��t�����<���5��n� ߳�ǿ{>x�@�9Z�K�wlA��˞A�׭���/_N�
+X(��Tb�>q\��`��{�����nl0� �4��z�QE�^}��:È� �#�W��k�Oi�5F�(�$nTe�7+gN�s�O��Ƞ�,���Ҽl��Sn
�\ ��>�f���Ƶ�O�0w!��������Yam{^(0��p��������$A���I��lO�T�5���cC�B�*?}�*Ǧ�h`�h{<NGƽ\i�"���<B�fHjpB�OnPA��2���'�B��%��zr���[#�󧏓B3���?'�o��y�"�@�J��d$Aq�|����l��+x�Ơ�u��E�� 7 6 <�:^��Ș � �Po��h1(�2 ��FDݽΰX;�v�u]��,ī3��+UP��pPq��c��txd�X�Le�pD>��j�)�J] ����dߠ��	vbm��Ѐ-FPU=u��>Z�o�X F���a��0�Y��TLz�	�tU˨M �)3V�V�,�ш��Wϟ��G�Pف����l��	���Z���=�k��`�9�.d���k�7&ᳶ������|�i�#����	�ذ��O����ַ��sp�a#��T��yZ$� ��\+L��~@ �
}-)Qǳ:����,,�#f� ���۸��p$@���M�\��YbN�g�w|s�FO&��ڃf���|5Pܗ��/�.�a�5�jx�0A��|������,�~#���|� �÷�?�>�)�痥ԈHxݧ]B] ���I�3�Jf�U*��T�y镋gO���a�~|�=Y_���ތ��xs���[(�\]���e�dh�pbB������gY��V��:�k�<X�z�M�^��|�����v�ݎ�	���AªȄ���+����[\�|� �b�s�aO�5�c�3�ט[�?>�E�<j�7�? �==�K�/����w�������5�9���#R�0��5�����0%�6@Ĺ@�������ǒ����},x�͠�eL2�gd|l��>���
(���M|�+ջ�#��|���B!��]^��[�o�W������2 ���ֶ<�o�����M�n����O-O����Ғ��n����5`��͘�g�$��� ~T��ع��cn >x��?���2��y'��Z��Jp�������ft�{�;?李�o��qg�-4��:{�L<*[�m����y�,-��P 	2�D�N�Z��V��h�����0x͈�����z�a*/��Z�*�%�b�8vTN������6��^f$	 ���%���]YZZ�A�&���r��g��R��?>6��a��@��ȑ)�A2�`��Z&��ԙ��o��lP���lK4�o��O��OnK(c'd04�jM��^��,$�.��b� �$"5��Ec��w�B��U!�/'��7���x�#�>�h��� f�<{xW���H��JM��U��E�9�\�(B�A�N��¾
A�*���ɨ��U��VS3*�8 ¢*t
��-v,dj̖`L�����Sg �)�N�&�kU�@
(�*p�q�� %cZO�-�l�T�G��{"�JUѸd�F��a)6Ё5�6{x%zj#/�A&D�&imP����$
��zC�*�ĐA��`^/3[rhrB�t�59v��jD�ј�4`����Q�Q���1����NM�3o�L�
�۳$(rr�j�5�����=
�=^x����YED�?��S6M����y�Z�G��]��1��Cr�"��.�(��]Hۛ�c��D3)P ��±��2@����ۨ>��۾c�x+���q���3��h�Vd�`�4��9��?o;�}����mt�7�}�s�{S�� �t4@�Ge#_��oߗ��n�WCq�4@mք����b�\h���4�b~K�ۛ2ܛ��/_���I��-�~*ϟ��`Q�N�&�Q3]D�7�dii�*4����ȡC��MΝ>!�fE"��d�=�8'�੻!"mx�tṾ��u|F�y���3{QtmO��x���?Hu�A1 ���&%��Ve~qQ��
�0d��Һ+����_���U%�Ll#����/ȫ�s/�����ɍR*}���U��Td>8����I6�{x:�#}�am������y����d%�&!=���zᬌ��0 � >*���~<_��+��}#�~�̹+o�B!_�0��sW ��͛�X,�竫��P�����1l����o*�Y���� �X>�7ä��`l7 o1컍P���'f����@����~7��_+��ma�}� ��/8�(@�56 oEC~Dd���(�Ƞ��xF��c7��/@����DR��_�����&#�h�Dk
�x���!U�*��������D�e&f��^G� ϼ^g$�	��R^���K���S'%����ʼ�.j�k�8DB��O>�΍��}P�������Gr��nH���� ��P_�p�����_�����"�v�ޕ��%92uLN�9-�TR
%�"��L��vA���_�;�OY4(��MXAzJ��8 ���(�X)��� ���N
 <x5��@��G^�ʁ�#��� �@�m� m;���x���dPh �s���Ó���m����u�^f$=zҭ�0�f�T?���Ӗ�D ��33�a�,u�1��%�1$���:g��r����^�,�8m�2���FOx�
�Ty�Ŝ��6���J�"gޯS�QU���D�Y�'~�T�-H��3�\�s1����aTN?]��V��dR�*��Gk�&�\�e����?��TϠڀ�)�2�hU�<0&W.^�3=�o��xO?�����h������+W�	��A�.�����2�fS�(��Ss�| ��k,Pa s��dж��4	d�}�]�d _(� �#	�BP����*��p|�,� ��8���X@�*�.�Ng+���QŤ�i�3����m�Z�'���sx6�T��)������i+��1���1' ў��){��ql���k��ͷ!;�q��<���y�BCp� I8*[Ųܺ�H�y�:)4���R��~�Q��Eߑ9b0$d�
ے�ސ�\B.�vN�&�%������Y[�g���5��А�gv���w9���#��o|]N;J ���ye��ڠ]����N����t�������9j��8�}�{}8�}(����-,ʣgOeee]ʕ
��t�B��7{�h���e��cb�A�s��@u�3]__��r9�r�"�T�|r�cy��!�wH�b���-0��L���=2J T�����#��q�\}�Rkh�\�k��7� �\����ګ2:4Ȭ+��X̍�1la��r�z�d��9O ߙ_�=�]��On��J�򟭬�b����X�>ڡռ��nr�����G>ӛ�	��(�������E@m7��;�������;�`�����΄_��\�=4���X[v>��!��њ�iO~�x�NV�"��C��Ȉ@�q.D-���Z�(��H���Ҙ�5�GuJ.Z��vZ���0s 9��,�tt&E�(���F=�a����`肜:6-�DD�ܗ��9�����@Sj�\�.�v_��v@���I_), @��h��9hN :�p~�g��L9*+�Kr��UY�ؐc'N���~Y^]���UId���?D ����On�*' ���18��<8�5�ע(<uP-�6���p��? �`��n���?}pG~�֟��,"�(\,kaQ*&	'��Bhy.�ls^��ѷ@#���(�k@�
�Ug��t4\���������K�l�;��"c�9Ҏk����C\wb��ZM��ŵA2������P]b�� �_/7d�����.�|}Xc�r�΋mꌣ���ET�� �� ��.ڙ+�H����@�-��Gze��!93uH��t*!k�K���R��1�Nʾ�!��jo��
�	<�חs^�C�m�=�nv\���+8�g�{�-�����aa������?��� �3-u�q~�x�4�l4@��-2�v�S�� 0A#0 O��u�Ԯfri��:�B�S�"u�=?�a����3���;+���E��A �Λӂ��l�Qs����]�}V��uz��W�Vc^��"�pTJ5��?��>�X>��b]�� ��L_��EB5�Ͽ�h�P�i4Y�Z.nK*ޔ��ɩ�G�/���暬,����gԂ�����>�8xH�FGe|� �׮]�Ǐ>Cr��a��7�!ǎ$
i�Рi�@1��|f.m���N��������5���k�
 ��ܼ<x�XW���ͲH�r���
JXxN(P�Fx�6A�U�T)��h@)�����/]�3gN�għ7o�g�?���ԝ�={������L��5ӏ�&D��58�2�sd��Z�x��!�����K�op�N"x4�� <��K��G���~���K?
}��FW �ۿ��Cw����j��FN�H9paZ���wf�|#�@���^��7��v,��w�04�-�� okC�u��O!�d�wF���E���@~�q���t��� ���p�w5��aDm�-bh�q;�E�݃�!pE��<�e��;9�*�QT���&e4��hZ\[E5�_Ut;~""��W��	A�%I5l�X�h$�/I4�q���Y#G�)�zI��-����� �I��򒬭�p��(����r��%���OEG= l��4�,	�+�<ٳg���L�M�������;���c�&���+YZ^�P��ӁY][��A���#��iLW��R�I�a
���(���.�¶Ĝ?Ȩe4ʆO(b���	)p�!�F����Tw�I�P?o^A�!/uH8Ⱥ������Cr��	9w��<tO���ea�{����q6p¦�"
�ѱ���z��Q�.�'Wj�LYd`��}s�
BH��UMaG6
�Z��zD:�VB9�
�-8��&��;�4�;B�����H�,6���lE�8Vk��BǸ��M4)��aI�J��v#�亊C��E���O��T_ �:R#�C�nD� ��>[��
Δ~T.��l�|�&�dLR����	��eS�R^%�A�949�x�:��T�;4���R�QB}0�s ���_�
8vZQ�;����s��"�xv��] �fմֽ�E۫X��<��r�}�T[�����擿�Z�ܢ��L�Z�᭨:�e-h��Vk`ҕ�Jf������eo7"����ĳ����~Z��T� ���5�k\�"���cM��u���?��/��ĚAV7�8��O�2�ƎĹ�(ttm]s�j���3�cr��1�?�G5&�+���r���伟=NΜ� =�>���dckK���U�@7����|�r�Є��<x6t �v$Р�ƒ\����f��3��n5-�P���;�EHсޣ���ۅ�<������� ��E'@d�XJ#�t�K��[���J�F��^��<0�eW����y��W�ԩ����w�,���֣��� �YY]�]D�{��2�0/O��P� YpPj,�/�6W��I��Ѭ���+22���F��v
ܢ�!R,סb�����p����>�n\�}�w~�w�o߾���|�?][[@����>�6�܉ja�_H��vN}'����~r����ԍI7W���mF�65�:��6��ۻ^���{����}N���ﲘ:����N���� ���Ϗ��;�W�}�%!��ѩMظ�ǳ0�Vb'���6*,
�jA&�����vL���H���R`��Ri	E���/H�
����0 M��}��S�Y�x���B�"�D�������e�|��ֶ��%	�>�= 
��iR!�!�R��B����<k��T�P�����)��A)l)��<��8�{���5�~�f#��@���I�oW����T8�.�9.������Y ��=:�5���`\Q��3B�kRAZE��p$��������)��-i��e�;    IDATRV��Ғ�`�����*P4��\��:���l�˩Z�۽���/�>{����B ��)�2�p�D�h�(K.�����#2?�B���{27�pscEz3)��"�|2��.�4�e�M�0ZQ;�T��"ۆ�����z�#��}k��H�{
43�n���W�.m��dsLCMF��;fKIAlj�[A�#D�Z�\�F8&Œĳ�2v���^�I	�Ǡd���b�Vޖ�k�>�)�9WL���˨4.��u_o��٭�Q$���h��6䡦D)o,K**rp“:~L�GGث�^���А�<~T��z���1i[l�ш�N�g�f�-Xdo|�5�ND�v�u�lt �2�\�^�]��_�5���>g׋���gEs݊;qns�l��;V�
���V�b[`Ů߮����OD�D�s�6-������� ��SbM��ƞ����e?�c�8�G�o�����<�4g�H8}�zS>�䎼�����F^B��D	AԔ���<�;��G��`�h��z��|ce��fS���l�T�oK��%��ޖ�ϟ������dt����O>�D�WW\:s�|��_�CH�YeV�DQ�d�"���l���h>G;����c���ᯑ��S�cb�gI�P����[Xb7V���	�{8vt)������I�Z��e*m�T.�E�e�2;Ϡo\ΝyE���������-y���g~�~����>}&�G$w��g�=���b�Q��?x�����N2#v��AԦ�ڱ�$�/
�1�A���.�`mS�I3���#f��#��ʉ3�~����������u�֯��忷���o �.�qCn���L>����q��`�6{�F I@���p�O��T��-<���ư��4�g�:}f�	�	X������9�:_����i�7� Ŧ�~ٌ���;�$��h�Ӟ��LS�.�j-TK�b�#��;�Bnn'��+0;��I֔e,��l$
5���߰ X��&���5��T"h�z�J=tL'%��i�+��)8�� (:����W=x�qх��2�h[ݨcA
����Q��0��@u�r�H�(��� ^3 ^
������@4�Yz�q��dm�$�d��$��tX��,�}����\�	�Y����A�B���G����,��-�����ޔ�O�$�ׯ ��:
;uREBۉ�(��j;X������𜟠~0�А���΃P3�g�Qo�?�WNO��)�{1#�����H���b~S��L4"��H�� Gs��>������p��N�X��2{�u�;�{�(�g�3[�rX����L�k-�y��o�CR�R ����EcQVr�є�X�r3$[����'^�ŭ-Y�(H��l՞�HHe }�95�k�ny��!
��<xK-��m �h=��f�$�V�����"u���}r`xP�	4�P%���i*P _��3I*	�ߊ-�&��f�ll�n5��̀-��p�����9A{j�4ʋ�p,����-0l�7�l/�~d��@���6�E�>Ck���8�>���짍��'�n��t̶
���� ����6Z��ظ�y��ɱ=v��(��I)�r��]�ӷ�R��eiD�R%3��Q�Z�x�s�8E��Oj� �PVB��ެ�z��LO�I&��ڲ|��U�@�iv�G)I�P��	%��\��X_��db��4e�H�����)Hm ���b�lx;�ց����m����;�.1.�bYV��eyiUV66dc#/+��N<�����uG�Ѡ�1X����1�lF�/�z����Y�������'2ЯJI��~��]F�=~�{o��L:Ďϛ�[���3%���>Uk ���#))QJ��<0&_z��dR1��F�t5��*~A0%_(����į�:w��n���n�����������j�������Qe��Jq��-ƽ&���Z'������<�F/k�k�̢�Q��=��������p�z_�w����w˗�D��
���؋��͌�mA osŜ,64µ���Q(Jj��&��:q�#	��#��P8B _vx��ҫVk� �7�z���|d{z�wR]B��	�I~���w�l���sFdl�����Ph��f��TJR��]�Ia�ރq��`~�'�Ir�� 
?i��oS��q�(-��D���}(>Յoc��{����)�a�Y?��(윋1j��P���z8F �e[M�% FD[j��Ri��p���CQ;n�p�x��5����v��'(�pM��&uL���͢dlT����h� ߗ
 �5fC$�8������D
��2#6 y�3�_Q�rk�5�;ʻ�}� �?��A�v0�QR���/�-�s0 ��`�3b��g9�c]�r��i9~�<x�B�ϯH-ek,F�ɝ��R������A-h<#�4 ��s������CX/�I�$��v������@�i&���#�ݘ�`���} ����·=G�",�lQp�{p�����}Ƣ�8��R?�lj�>�
fɱO����-���w^����:��~���ߴ�`gh'Hog ���Äsa�Ĩ7������|���ym��zj���Ѳ�7s\�z5��F�2�5�7o3�Y�2SR��qAm L���6>pA�6U�՜�Q`�� G�\�t4,'������^�@������mfazz��9�V�7 ��)"�^9#_����I�V�(��.����. ������"�c{a� ��Y| O�KQ#�K�+- ����=j2�!c����3p�v/<��-m8
 �g��
�Mh�GI}���Twz��9�&�g礯7'?�s?���7>�����";�b/;t�:t������5�o?> <�4 ���*՚pr�"'��ʕ�QaB #h�{���Ǜ�b��c����\�;�u��o��o�{����7�K+++9�P3 �`v���43��i��(������t�}p4�������x#�4V������z������7������s���q��2�_r�z�Ɋ<�QYr#��2�QXV �V� o��D&G���U���H*h7 o�A7�6(A�A�d�r�}��dQ��:i3�L#:�7u�h�ԥV)J�V�pEI�tߒ�L��^��)�.�fK���������~!j�q"q
Ǘk�� �`�D�-P�>ӐK5��R}|8(h^��d�hT��7��0v���Uj#ʳ�q�a��أ�Tc�|S�����x0�y����H(��XON�n��śm�e�r�5u �'F��vxd5h�=���k�#"=�u�s�R�PX��G!^�D
͹S.?3+�_���Lo <Dsk�M	�
�$GGC�(�h��f64%_'?�������Cp��~�>v|��  oM�6��m>����5��SF�U/ԟ���I�֔���R2u�8��\Gw�EiPb4��d$���ԓN6�Y� �����c�Oู;+���s`���$�DBз��%I2a��p������}r����$��`s�����ap\�y���66��0��Z?��m���}?��SJ����~���Σ�6��q�z�~,(���i����_�z:x|`0�&<F���(4�}ˎ�y�h�}���s�-���p:�"�
saԑ��J����ܓ7��+Y�E���@c6��޼l�?�l������l�0�'�C�r`�O���T�E��y*�?�Bn�Sv�s ��jU�F��������פ/��z��n�B��5A-J)��'b��ΰ��?�ڬ��{{hm 5�K��ږ���YX���-�,���uF׎��=`�,]���8�8;Ik���vp��������ܜܼ񑬯�I*��
�Xo��T���@��dzz������3�'c184��=~�JQp����ZU������MҜ ����>#���7�Ii�\k��R���;}��~�ۮ �����q�!wyy9�Jx[4�V-B����нt���ʽ �- ������ �vL������q6��� 0�<��f�������u��vZ���N��{���i��x=�x�ϮeHCm �	�7�¶�~<��& <�@NM׺>W2�	@���$��g����K!`d�U#�}W�n:��{�����\_��ol��֦
�������F]�u�ax���׬JOO���jI�0�R�l��ڪR��/�5�^);z�c��8�i�ṃF�-�;��ل�����w -�Ǣ�E�(�I�RT���z$��apD�����\^Z��ͼ�Cqi�#Ҩ�$*�o�5�JD�9��C��t�r�4���CB�n�|$�#�l�4�1j�3�Z�N\Ѣ��m�Kg��Z��Ft@}�
%��;�g����]�"Q(�4���s'���cGdqfN>x�:%��4�ICF2T���dw�H�\*H�eP)vg]�UX?�۫ۺk�eW��^���`���$ sru����6� �����㔃"g5�
X��C�H4��p<������z�cF���i�dh8"�PL�op�S���N*����{���;�� ؓ^Vz%,jei��$�Sg9KOFF�rrxbBN�b���Ɉ$�(m��`����;=�����}ʛ�>M
����{���a�| j���Ì�bT\���]�Y@��l/��U����l���������G��q��팮��^l_�1��n��w;������R�D狿�sݺ��j���~j6 ��
eC��r������kR�v�M����%�w��9wQ��T���'�����A�?���ƪ�<}"s/ZE�6�po�G��&_�t��t/����H�lLiq���w�tu�a����۸v�����Xo(��Z�|�D����^ݔ"5ҵ�,��W� �ݮ�[^^����t���,�v<Pu�V^�p�*nh�<�чG��o�T%tB�:���?yJ��$�9����<�B ��)4 �.6��n�̂�k�K$�+ ��8W�8/$�'�o���o�N��������
��7s�޽;�]�Z���������" >���ͨ�z�����������m�����}L����wۘ옻m���^dl���+��N�g\\{]W�k���Ȅ�.��Ch|Ss�#�F���Q�3v��g4�,NI$��L�@�om�|�� �	��FQ�h<�5���蘤2iYZ\֎nu4l�P�	��O��Q�*���j�N&���I�:rP���K���y!��󎋧�66��tcc{��g�q	EQ��h[�C�M)��Ȳnǈ�c�t���*|�1:čOLH�� ;�${��v��S��,�n�9HRɜ��5�TkB�m(����Wo|�~����Kin�Q�#�I0 _�3 ����d�t~�ȰQ^vlvVt
v������m5B)4.�H�ՠY4j
��Q9zZNL�Źy���G�0��&,�rY��Iʦ$�<'��%���Y[��P������1R쮙)tr����YI�w8�s,}ӊ`5��VA]:-���i*�Z����HP�,%fN𓥠-Y�v�6R�p4��h{r() ����J��O��&�FLʉ���7��h8.�Gu*���a��v������cn�E�1��(S��FYW�}�v�R-lJ&�\:-�8�|\�z3rdr��m�F��!���A�J9� �6~��Γo�qƧ�A�^��v���{^��
�&�g�3�9���A�}�>�G�� ]�[�1�h��)�8��מ��|�N��J���:���8���)4/�w�ۺ��>�|u:�����w��?��~@��o�{ ?���2��%�:�)5q�kgF�օ��y��@��Reo��\V^9q���O�ާ�dei��hx��)bOſx,"�ٜ|��K���2h�W'��:KjZ�7�¹�ho���	:������={����R�*U^�B�����(��G���9��[[ۤ!ӌW,�5bx�{kOF/����Μ>I
�_�H�6������7~���~�m6B�}�88)LH	���lm�'�X9L}�۷>��O�j�HR�Ui��'U����Ċg�������x��j�Z������������v�`�]�w����۷o������ ~C77�Zw����D�}��ɛ�o�`a`lQZ�ª�qm>��O_�c�#�A໛W��N�Խ^{����k��^G�}k��T+�G�T�J���|C�:�+�4�h�Se���QĊh-"� ��c�ll��%Uh��$Qi/M���TD&�:�-� <"��+k�� �G*E�!u6�	I
� ����(b�H*��'����W��zrbL�=}H9)D ���!��{ s�p+k˚)
71�&�H�skr����|�T�N|:&��B�ӆǚ�G tzJ�''e������]]p�P��λ��{W?�p(%=���R���hz�I��O �"�Z��v���tED�񘄲9�dz$���32e��d$�g�VwE��-�o��~���TzZ@����6�o��(� /-�����Srrz��a�>�H��AJs$��#Fe{iVf&��2=u�ҠڶI瓪7P֫"�c����	`r����@�,+�S��C��$�L!���� �#�I���T��_�X��'�w�#�C��DHc#�;8<"�TN?�eӚ�r��+���evi]ꨧ��M�:ޭ�z�E��(���=X:�N>t�r ��v�1ie���.�"��d�q��xX$���@OJ&�����r���)��eπ�Tp�=��@?�#p�����"�����<l�?��쯽o�6�����(���d������{�����5 �;�ql:C�]U��1���+���������X�V�����n�מ�m~�������*}�'u���	YXY���"�]��>�p`��wQ�V1��ȉ6B���J��C5�n����?$��2���ܿ}[ʥm�e��>'�f�%m��W��&�/]��lB�����%�z��Kxۗw���5�����Nx�(���HefnA���!��32_�Mu�	τ�2��ux�lѬ���z\'�/8,���>u��f����7o����Z�x��7��3y��7�o`����EV7�Y4����񑩣2>>�4n�����ʶ������9}B1��B���M� 3 ���r���7��������{�->�n����?Z]]�����'��P���d�E�?h�۲h��E�ގ��~�7A��㞿 ���^ ��c�2B_ �)߈uZ��-2�Hw�\�Q�6O|�h*,0,L����Ѵ焟ܔ�j�u� ���E���2l��^fS=},b~y}�E����?�M��^X� (��e4BI.$�WV�	��iBC�"�&=T[A{���!�Ȁ(��!9~bJ.�?'��e��G�df�y���w���3�A&��7�qXY[�����:8��TNˋ��X���b3���d��19|������=CF5!��fd ӛ�B�(K�+���s_��c���-������V֦X0�p���$3s=���I#�TU%��q ���g�BF ��h6G _�frR���k\�D1uk�{Ԋ�<3 �`:)T��+��<���;��}��
�5ojx�p��o����Tx���z���"�M�{��I˥��K__/4%*I�w�ӑ��袡��� o�R����=ü`C2�;x\�w���P������Nr����g�4]'�[YYߐj�!C�Ƥ֌ʻ~$/We��A9s���w��ª4`s�������l��N���l��	�����L=����h��L�ByKz�	ɥS5%�H_6)FU���iJ��1W	�v�D�f'7?i;@�s�Z�f��y�p���,��~�ߞ�^޻��� ڷ�����i{����o����<��x�nXt�7�d���m;�������2׷�Iܿ���j����A'�h��:g�
L�rcA'p�0B�Du4    IDAT���O�/޾*7�>I���@H��y1G���]��B�o�S���W��ސ���L>� ����4�eI'��d��`>�2��H��ep�A�y���˦%���YE H����֗O�����N�S�3�z~�T;��?~�Fḇ� ����.���^�����Ɩlnm�|K*�V�f��W ��.�� wlA1�^'�jwu��H����Ξ���I���%w��ߦL$�#���D�z�-����c<���<��G@�Gt~bb�{�Cts�AuF鱘�*e�$:��T
:ybZb��T�%I��_����j�_M���G��z�N��N���wG߻�66iuu5G>�FU�@!���moYO�Er���O�H��qd4�tZWOO�ٮ'�ɴ�_�5H:���?��@����X����w[ߨwZ��3���i��E*�ɘ#f��v�:5�Qf�~`�6�&KiRh��B�a��DcqY\ݐՍ� �
�HD�;�d���m��AXB�z:%���hp�F#q8	�Q]��b9z�(d�=�p�$�l��(��~Y�zE���X�"Gt���	��p����'SSS299.��>�?{����SmD�t�Ma�c���T��*2�
 ��+�^�$��ַ��[Y_��]��:{��}�Z��.P��77��w>�kޔz9,�HJj���kD��m��\N�==RO"�ޔf�,1t`\Y�P���4��=��dF���FAջF�,�^��a� ����B-u�-�ތ]�R�#�р��7���AB�kU�IYr���;
͔,�/ɵ���m7��j�(�z2��W/���aY�y�n��NLK?d5�ȣ�v��4� y���r׊os|p��qOh
�:�ElQ�L����*��@b��a@N����c��;�2��'!��b�6������@w�RnH&7 �XJ���_��<wQ&����^�H�,����ad�(���}gO�9�\��K�,��#�ҽU�~��@"�N��wd�jҨ�%�IJ��K.��T��Μ<&�d�8l��η�I����~Z�����/x��}@�G��&�M7���h��v��6�iŞA@m���E��c�9$����`[�?�{��۵�Ί��vgV����ԕ�O`� �a
ؚn�t|�t��]G[kv���߶1�3u0s&�4��7%_(��ʺ��_�?��x�O�K��Z���q�}����r�: p��9_)k��Z��^ý=r���R��?���Z�	퓂� ��{�&���_���=sFz�((���m,g���*Ơ6�Q�Ɠ�cds̞����ݰ�?�>���a�	�^��*%2gfd~qI��7	෶�ќSZs�������5w&+����g�L8�_�XU�M�I����K�[�����"W�'�#��1����+G�N�ŋ��\[[S�h�&�=x(���2>9AG`kc�xt7��2���C� >�I��W/��C��#
 <�	����o�Z�{�ϝ����������v������mnl�=��`�� �ܥ��*�
о(����D
YL,�N��8�� ('9��Wг�#���xDݢ�"�����n��o\w�Sqv���ר��{�<�6 o������"U@<�w�b�rQ�4U
�x��4 ��Ub��T�=;�Vrɍ/�oQu.ɤ��\���xhE#JB�c�q^P����t�Z�h,$Ǧ����$�MH���J
4ɀ��L���<y�P��9��ݡ��������_<x@ �v˸.���<�qB����!��S�����!�t�|獿%&��ً�ɻ?��AZ/ۗc��68�H!�R��w��<~4#�F� �YU��VyJd*+�r9��d�G�tǬK��K+�,%���f����p&���PD����ţ�1��n���t<�-n��5�2�������رI�#�Ʌ�.�m����f�E�gOM���iY����|$��Ri��u��[_�$�'���*�ޒ��!6Ⲏ�np���K�#�B8�ж�[�Uמ 
�a���q�q=2pe �)H�� ��{m���<�8ߠ3Y'L;n��Q��)�)V%�;D ��?��_ْ�g�����;^��sK��@�k8��fOu���״Cf�{Rp��I��6�J���a�9 ?� |�Y�l*.�x�xO2J��ެL�$�&��Kb��A�g{�|��h�C��m8����mn�2pm�3��M��惁K�/|���T�8�*&9Y^���9�v->�x�������߆�s�G�w8s.k�G���8~�T��pޛ���� ���{�Y�6߶��*(&ciό�G�Vm�-,�����?�Og$��Q�v��#�x�� qu*t�+u�s�Kp���}�H?�G g�C�<l��P�� �SG&�_�2��l;�_��
��x�sN:i� v���_���=v��s�i�# �{C+4�_��2ʽ��"�����������Vڔ�tl00G�RC��l��aeu��ڃ<2�������,9��y��z�*�A6����t"0?��h<|���e�������<��6:���0�Zo��`�|��%�m�\�NEgH��B�_8 �U������3�xr��l`����]����_�X]������bQyF�@ɇb��f�Ht:�^�^�ߟ �D��ж�m�ۏn���o4�k�'���n���}/��1ZMov[0;��NwKs	�� �������^���N��3��������Î�U�H�1r˶���&3�hA$FI,쥵M�Ց�$�ZB�2�n��`Q�S��9�L�d`x����B��SA����Yh��; ӍuEt��\Z��r
#��q�QL��ږ͕5��#��E�V�O�=f���'�����@�>W}�l��5 sS|$���a9{�|��_�ѱ�|fV~������3�"2���!�JE;�F�����F�][c�)4�:��b]|�R����e%�IK >�`f"T,��ܜ��%I���װ&e���^I��R�b��4(�X|��0\��=x�wAP���8�"XNF�5�ݨE�po�W�`j��)S� �/�s������˵n0�<���	��W^�K��J-�.�ܔ��ؿ�NP7�)��9�����((ژȨ-~Q��o-n�CfŮ
*U�m@�|y� im����P���ܷ�������F�1? ���[bGށ��R�����e�P�cg����iy��G�baE�S����iwd�A�L����j�ޗ�"�p�[���cc�N�_D' ��4$��Q=**uɤ��M�d�'-GN�Y �#�A������hs��`ֿf�trĂ�Ə�����{@��S�m'@o`ٿw��MG!��]/�+�"�
��E�~!��m�G�1�Biem o ��vO��9<}�K��h<�3�vT��H�~�:�f@7I�Z�مe�7o�P���p2+%�9�%�B��~�@�q��9㸼N�q
a�rE���ȉ#��gd��Cy��3j�C� *i����>�N��у�|EΜ>N ���"cOb� �l`�]�
>��3�$8��@���9�A���|����Rn�M��.����,���F��K��4�iBx6�C(�%���y���8ƫX�3 <(2P��'�!�F��4�T��?}���`�x8�tE��x}k����|���M*�@����CtQiVk���|��eC��z�u
T�0���[��j���O�<�?�><���������/���gsO������hqi�z�� O�c�N�Vp�u;O'���i?/4r~Ԃ��K[���g/�����"��$��΅��P}�G�搪�uEu����idv4�jg7 oF��#�k7��?�/�[.R[�A���������!K��'d&�qAכ�� E��+��.�(`U ��(�W��K�_M��/����Ȩ�keY^]adF2@� ��/� 4�q�@��<DAꍲvZu��p�P�A��/���I���2:33#w�ަ���X�lO������!�PP��J"����q��:&=�}��/���d~a�� i�wD�D�h#	����&%�&P�R��@0s4.�����i��R>f�Q,�֋�RQ��$� ��h����@�E#�B*�H�;�x��t�+�c�P�"�F�h�X�G��v2c�&�`2$���G!*U�����'��v����u�[\b�8��ɿ������	�\��g�����D�!-�k�^9�	�xdnLm��7 o�� �_�j2��x�8 �|ްo|�¬�X1^��OՋ�1z�N�\0C�vt�	�ݣ�м�]�B�"}������@6
�:sNƏ	�s��9���^����N�Fŝ]`TP#��5� <7R���o���K*�d<ʦj�tLz�Q��&�D�	������X�@�$�2�>`5{tD�9ᧁF߱������?-�n�ߖ�r�[�ñ,��������G�n��`�������X����l^�ިΝj����#�v-�۪+ѽ$������w2����mcf��"\S�uҴ�T�u��YBJ��<���?��ɳ�i��R����L�yo݅] s+����� ���D�M�oQh#[���h��$x���d�t)���Tm�[����=sR��]�������:x�V��⋝��A,`��g8��~�9� ��A)Z���>���!��۲��&�[y���ՙ�r��s
��)J&��P��:�~�i� �_���4qd0�i�1#{])�H����"j�����{w�Z���e�мx�K�E���`BF8`ddP^���F�D ��0x�$��z�!�ǉs�����Ԣo+��������w�����qaa���b��GP j>/���":�w�4����mb�Qԅݖ13�e��>�)ߞX��n��M��q7��/�n@?�P��c�S�鸾A:B|ϋx�8�����k/�vQQ�i����9
���y��lS$�>iP ¬w��El����X4j"71B<Y �W6!#�Z���0M �o����!.^xߘ�X�i46jT�G�p�P�j�r���u^`L��[��)MȚ֫�>OØ Z�0� Y�B1υ�.m�>C����fh� �4M�wNЕ�#I��Ym4i���$�E�*�qD�2FG��4k��@	��<|$�.��N1�*yH]6�ٞ�%�Ϡ���N.4 |�o�� |D��Lluv07@)-��M�:�q�&#��G㠒�G�~�E��z��깓r��<�\޿��=C��.�ل���~CN> ���e��g2>:$c��1S��	CnV���ߑ�5�GJ1ҡ��d��Z�F��G�QB�[�<���F�� ��|PhW7Y"d?P�����D�7�c3	�0�z"��
�`�8Ţe��(�H�Iȟ��[���)GN�"c���;ސ��e�H��	֛h5�kfc��;Pf�v�u_��c֣�Y��RgHE�������KUR�0�N""�z� ����a�����8&����|r?jl�1��� ���G�;�xs|z�Q:���^�ϙC�SIl�����xXc����#i�s�{f�m^���3w��pE��hc��|uF�x��g�s�C����6&>���^\0Ͼ�}�z�q�
h�9|_iU��R����������,mH3�"�����v�S���eț��5�{	�WY�:ԟ��S��?����˓��I�\�l:ɽz� �R�1�I&���#�������r���fU��o����	/�Lt���ǝ��Acs�~Z�V�C����5��	�P� ��dss[6��4i��:h"-�YJ�ԋ�d�ف��w��:�j�PcA����Ǐ˅s����W*���A��6U��p�}�����jv�;�ame���:�����>�K__9��G��g�����8dy�����¹K�ѳ�����?]�����O̼�������l�P ���b�7���5{p��������f�T�A=� ��m�Y���{r' �7	����y���b��f�[Խ��5�a@݀<X���\Pa��q�MF�R�0��ކXP:ٍ�B<(4�[���r#�F; 8�n:�XHI���J���$���X�h� D\mRca'��ڨ�|LC���@(8 Iu�65� .b�R�b	m��=�d���9(������-��+��a��v7��h$-��
�|Cq2����[���������rH�(��,F4&�lVB�d��#aF���<<#Ρ�r��9��Q �N8�0���N�K+2��+W�ߊ��1Xg`����0�5��E�A���j2ؗ ��>:%/�>��޽N _cAjCFsi�ş���>r@�5�񀲄P���JQלN/T^�2���u�G�:�C,
Lb���nc��Y���o"� |M�x@�<�y��.,�bru@���$�HJ��"6Pa���F�(-_i���?�ŵm�����?z	��Q�]ӥ�B��� h8~�{�̌>����8���]���F�+�W%��H*��Z|2*җ�SB�S�I��\+9���4�ܯ|�b�O' �߯���������(x����7v�Q��k�:�&Y�� �7��U�x��f �ev|�>���G��9h�sv��}��������߿�}t.c��6�v_����|��k�O>������s �J�!��?���'2��)�h��
P�`�8�n���=�9f�+��B�  J1�r�; ���Ct<�<�G|�\ -k`ks��[���d�I*d�z�|��_��	군��!�0d_��L�5��h�|'l�S��nأ�k�Zv�e�1�Np�gf�duc��O���6iI3A�r�'���'3is�8�{�FK��h�cm��˦	�����xְ���F]�@��f6gT o]��,�t�{��$�9�, <t���s�F�1��]�jC������47>����}�������;�������������e��"' <[�;�}�`���_�ݢ����Ac����Y�����g��fm����D6�ǿkގ�3�cw�؝��A��[g
MpC���1���y�E�lS�G�/�F��A�ȇEKa�&�"u�<p��74k������di}[��H0�c�P��pQ>�o���T:K=�R� �rI�={&��M*����7��⡉�ʴ�v]9����[A���`<�\�1E�7���R-2mn\�	鬢:�8�SP2u{~�FB���x\;��cЙE4�� ����Z<zn�@����mQ �����;��XB�ٌԓq�G��A�6����f�K޷������8z��ѱ�x��m|^Z�s�a}�T��rʻxPh��v�4�̳��ğ_\�
6�F]������7���QI�j���BJyt�]c����I�ӵ�:BF�$��#�P�+h�N�n��ƴc/6�c5`�x	Z�i���ڛ,%�����;�'8pUz�j���k͈d�����ŵ-�����v� ~��Q����5t`�%�g��
W!�v^�������N}��騬j��O{�8�h� ��6�G�+ ��J�Y�2}�`���H�qJH�fuh��t�C��og�&@��z�ؾ�� `�%�ׂW6/� � ��g�����E���ߏ\�}�cP���_�����YB\�c�c揵ݻK��v������,�n��M�P/;��Q}
1T��[�ɟ��mY��K-�:)�*ɪv�cG4���lP<�	���>z0�JP��S��/������������r��[�xlN�G���#��vA�������)iT�Tf�g:p,�o� E�ALd����d���3|��0<f����g��c��P,����<y�� >�Y�5�&aJ �#�|џ�%�@�q�S�>����Z��/�HG2�|�֮����K���iA���p���Nb�`�U}F]�/1�#��\����K�Zd�1"�<�	EvF"(b]n�¿q����ꝘXl�L��     IDAT�����?��G��<�'k��?3??�)�5������6⌐�,#�,z��	��۾�7��z�� c��-d�h�Q��\��Z ; Z�c�����BϮC�5hy9�d�ߦ��)&���_ ���{Scg[�i?wr_�X�+�;5�n�}��V�c �	x<?�J�X\����$��6�L������X7OKO� ��<�]$��91�p��õ�+������Ҝ|�<���28�/�L���ಕ+�~9?�)�O4��V���8�ܐ����"#��t�S������ ) _��y��7�	��5d���Z�k8�h�g�L�$�V��>S�8ē)�4�=5;��b*%��rH�2���4#.���@� �#�DTjpN�G֍��|Q2	+bmH�UO/#�8�F��A"D��� �7�����+[Um��W�J`�w�D;���y��+���Y�FNK�R������?�;ߑ��$kHy{�]>װlo�h�=<��3���:g�#�� 	@w��,�5x�ؕ�ͺ4�+��6� ��p�@1<Y�d�R����hku�;6�$��zŀ��Ȋy�@K�$�K,��d�WW6����dy� �O�a��>����!P�B1Rhv�&��	��������i\[.�d -��PF���XH{��h;zH�����`S|+�
��t�&0�t��u}w���i�%h���>�E�0`�x�c���b|��>x�q��E�͡��|~���;>��wL�Qm��>G^��y��os��6&vOȘX4=�9��Tp|²���s�3�{���X�{�kPI�ʄ8��{���SY�.
�i-Ϭ��<6�J>�^ۀI*�nB��"�5!��C}rr����	y E@��t��<�{�� ۔�ޒ��MF�aG �у䵋��[�����:F~5D@E�c�:!Cpvg+g,Uh�kӟ�A,b��w�|��������40��y�����G�(Rեb�"�GGv��
Bϥ�E����躹����AgF����,82�����x2���#aI������a�p.�И,(>��f������\O�zs2q`�\�pVzs=R-n���΀�t[ ~����g��������� ����wzy}�YY^����\��ϳb���Ԛ��/�!/M/��k�-�{f�������4�h�eK��cB;y�Tf#�Fy(-悇m��L���\$�:Z���"�"�]����h(�k�W�
�l��b���ܜ� r'lo8Z��)�v#�H� �E�|��V_輀u<wv�k/Z�[��vn1�z�I������Eyts��"��@�f�v\E�XF:3&�#cR�d$9�%_�Уc���T]�d�4� �i7����)������X,��'�p���V�G���$��ۼ�u�G��h�����c!�Ӿo�L˜ˉd\�x@�,����v9.�TRi�%*���D�1)���c�?#v��c�Z�M�	����D��\�NհԪ���c�!GfA#��HB���I6qjP��))lf��ω�F*�i`h���Ij�� ���S0MЄG-��F�`U7�Hk�U�u����"V�U�C�.����Z<�M�7�y�d*=֫қIʫ����'danV�]�Ɔ!�:2( ��s�r��~Ʉ�C-D� ŭu��\��/ƻo���X<�b�ȹe�w�Ɏ���DbI'��N�v�ə7:�ECV����]1���R`C4�/uo�� ��	��M��#߳֔d&+�T�)z��I$�f����޿����:qZ�>*�|Ў���9����nK���V�l�ǑU{�F_m����<�3�:�6cN\de�@����$���`<n�Uy6������9x`T��0�� �N������Xx?.z�^������M���ր�z����G��s��mL�����������|��n�u|/Y���pl����s�5��h�1�Ü;��>s8�\����c}'��<~�������5 ��5�!�l���� ������l��ʮ��&_z����;$��2�H���|P��n�L���t�D����H%}�1�����QK]U�b�"	� A� 	�0�Df"�{��������w�%Eg+��\s�9�����k�Rj4壻��;\��RU������r.+���7��u�(��^�ޘ�U0�ac��po�ڿ�v��g���/����tv�9��g͕S��"�@_/����7d��TӢ�/�+"v�&��:5���f?Kb����[8��ieX#+��22���
��r� �3�k�I�e]�RM!Ռ߈�/.-h=R�F���(�S��	<�\�ќT�x�q�������b�>��k��m����o2�.��ɷ<0��L*��7ο.#�C�?����%�
E�ʯ6�2�bv"���o?��}}}�X���5�ǿ���{����Ϳ�9?�|,[ZY%��.�WL��|���� ���v ތ�3 鴂���q�y� 8�wmZ¸�h�J�?9��u~4�@F0���<��7��tm��#Pc�E���c69��9G*�ɦ��#�Ҡ1J-wǡ��>����~�*Q����m(��������~cQ�G������*	:��x��a���Ţy�)�0s�>)כ��7(�|A�דɍbԇ�����i����\���d��������iP�xF1ˁ�0�%2�]�:���E��1�9��Ƣn�у������/���FR.�ƍ���j��;rt0���e�\���Y���������F�R��X�z�vD����.���E�qj �]y��CW>١zd����3y�g��LӚIOiU����(4H֤��B�� <��|x�qNr�]���ʍ�2�����H�Y(��CW���������� ��d_D����MUx�fxwWAN>̖��������+[-�8�"��=��<'{6�J!Q���j%i6*,�ǼX�F�6��� O�f���rBU,,v�H�i43�����T��<8w>��YW��".�c�=� �%�6^�����v�Y+��T�<^"����e���eٲ�o�&�_�H�MM�iW�KMH4��.p`��h����D���ʀ:@@;�*<ڦ�FE��p�<סB���^&)ґ�KG&Ɉ���[e׶�,nEmv|�{�F���ܚ-���� ��*7����G��R,��x[����[=�#��p��5�a������{��v����lǵq��>�i�����F�c�{���8m����ֈ?�~��(� �)77@+cS � ����|t�y��UY,� r�a�#Aנ�y�7�1�f���y�cJ]�� ��JO>%�zW}��W��Ŕ5Y^�'=A�$� ����u�����[��%�0����X#�9 o��D4{:>������Th�,��NC`��8",h6t�*5�����K+(Z]��jIV�(]fV ���,/q_�\E�	K�~��Oq��7��̕�0R�N#�����e`��}G�Ưcɦ2��}fph��op��Bw��+2��G��}���� �\y>53��������������" �����37?�����ON<� ��뫗C�|���9cF?�7��qZ"ء��-D+��"Ct5_�iA�:�Y�>V�0�����Ȼ=��'R�c4	UW�C{�@z�_�àxx��f� �_�I�C�x Zx���y��QZ�@���vc��ce�7��WԌg�ȣ�\�k�����Fޢ���m~�������
t]#p^AO��b&/��>�vt��-;���)�/?�G���Ғ�y R���Yx�� �m�6����J>�y�@y��|� ��6F��pl�a����T��J�����ȨnD���`�ш�6?F_5͍s�0�謊�P5�G��h�E�f�4(Ѕ ���$��1J��.���&Px={��Ĩ�H��D$1A�v���2����Sq��,��Sp�W�#���x�H
�H"> �6���P��pM�T���P
��QQS�Lc���j�k�<�E8>p'�O��.s����8wu��cGd��]2��ܸz� �TEUE����w�<+{6�H>Y��OS1���07VKE21�M�Fd,�`@���9�>@���+S�8�":SF�1`�ش)8�B�Qh�Ds0BZ�]�E%۠L���kL������%�ӿ���E������޵��ljF��pF�1�T�i�	�{{�G�s�F�_?�m�p x�p� �Q�F��hd��6�qx ��4)��f#�}��K
��޻�6t�:.�6�N b����F�|"jR�`����v���T��T?�n�����ٵ���]�]�o�^-�o�g��d��n���Џ�����������]��ֲvڀyߡ���qGЌi��-)�l���d��R�ɇw>��/^&�G'D��}��'8+�Wä�h^�h�/��^�"��=r����&���;����WK��lo�.��eI&��L:.�R��{v�/}れ�K6#%6+�V�iX	�x>�����w���"T��x��,;0>�}��C,}:���,��/��^a�IMv��\/(���#Pk?x�.~ؕ�6޺9m�<(���vŌT���T|iG�e<�|��u�5��"�	�x�x��?}�<��2��Ҳ��hP���5
�J ~,���?:��_-�sv�������?�;=���f�O���O�W�J���og[.&����h�$�������߹LV�΢RR����X(� `C�b�74��X���E��	����0�Q$������S�Ɂ
�Q L-7�)b�BZ��s�	6F���t�ݸ2|m6�Э���?� ��=.�n 
��x��9M��T��`L#)t�-�'���,lQ�*���\�I�Ld��+�#�ԪFj��'����	YY)
f��49�?h8�׭�}���	�2p`�qK���MҸ�!c+{�.�8 ��Z���Ӂt4lF�C�v)�ղ6���.Za�{��g2:F0p�+�� �V��d�b)'�&�z�f5:Kc��TR�в�7�X�ѥRX�ii�4�;��ˈ���l�~1�'b�`V��M���,�O�I��"��PJ���4�Y�uuK
���GJ)b���x$�e�u�BCW���v�t��e#5`٩'��	�� ٘��O�
3xU�?y�#��cc�! <�ɨ��e��S~�«�}�_rR�<��F�; <U}��D��r�Iͣ���4���F�OVx:u:_I��ٽn�-�bN�H}�	��c�����y+�?�a����#��;��8�;��p����0Ѷb�drv^����L/Vd��c2�a��{��<���sg�9��u�b|H�[�Ϻ��~C��guu�2����̫�W�@��I2�|d�#��Ͳ�H��ȒT�#�TuN����v�έ���GweH�r~x������F�,�_o_ہ�}�@c4z<W��g�gd
B�������ǿ���_����u�Z�;
��zm������w����� d�!�yk��?�옌\�: <���:Z��^�V�@<��bHyDN)�R��wR��,��r��=x46+S������Ӗ!'^pYx�4 ��� |qeY�����ʉ��	��~|K��="��'�*}���tafV
�99r`�����2<8@�XuZX�.�"r�H�v; ��{�}�13Z�?�v�(���gHBpI����<;�^�v���x=_(H�RS���iLPT
ۚL�{���0
5q'�l��4p�ɍc�e����\�yd�X�А&p��e�H}0
�k���u���$ߙ���~� tvvȶ-�����2:<LǐrմofI8��K5Ph�t�����ultT�@~�Ϛ ���ϟ�|1�ݙ�) �$ �E�}��{-��5x�%���e�FhuajD�����(�Q�nxD\������]�iia�&�"X�G،��������塸�Gm�#-�c)~���S6g�c�W���&�c����������n���n����磯��u���i���gS��'��g�h� �G����h�=+6���FAi�Sz��Xm���y�b^*0��1��p.X�j�Tes��-[6	T�0�n�x��$��Zk@�f�PMcx��Q����I����BG�h �eQb�B�^;�ׁ�����g�eҷR��� C�#244��D0�:���TÂVD�;r��.-.�������,,�zC�	�������� �)շ��NuiQ���$V\��$�X�:���:�$�Q�d*#�DJ���	��j���8-} ���Qh��hwX���Pa䉉�K�0�@i�5�
MCR��֫���)'���� ��)�A`s6��wΟ�����i�I�A>�nzu��3��Ͱ���e���+~�$�M��y�0�ìw��G�/
��5����)����M�k���n��.;0�Sp~�a( S��k-����������jCv9.���;������4 ;
� J�z�H*�ȄOR4i &��;@���Ivͪ�����06���ف\�T�,�t�\aD��B3��E �m��  �
2[�Z������A���e���6 ��@����~���R���0��5?�����3���D|�� ��<����v,�G�rc���i^6��=
ޣğ�]@���:�R��QY�w�.D��W�r������T���B�( .$�:ʇ�kjD \h �F�$���;3q���1R� ��Dt�:ҙ�I�Z�g��H.���Ϟ��_���>xa�Аb��~�?f?�l	���VdbN���|D�9��`���G���/��=,��[��Lk_
���xt^AǬk�&N����
�a�L.>ױ���G��}��A��f�=<�ۀʇ�!`�����gX��
ɠ�L5���}��x�y��ddddD:@	bp���{�aP&]��x��ғ�s_�������m,�Q�[~�Ϛ �w���w��٩ߟ��>�b��K >���ܰA��_�q3"zN�����Si�Hn��F�jS
�3p�]G��h֊L"��Z ��{,dD8]����zXI�]������9�����}Wi�#l��o�����Z����b������ �; x�_%�6&���y2�m�X��h����x�"��3PII���=�)��̼����
���ݜtZ-2频X��G�1�{C��7��q��wW�5���B��Z.�g�)ٴa��߻Wz�{�Q\����e�勒:
�x��(�y��!���ʵk�uh�#�)���d��r��qٴi�>x�h��?4�̔�qj`�)6�`tuU>�H���ԩG�5�^��1�����Q����C �KҕJKӤ�	)B� �!�l��*e8
���0j�;���!r�>��ݲQ�������ۺ���xǁԎ� ����!'���{v���S�~�*��k�Ȗ��օ��e�G��UI5+����	��a�VSKB�ۧϰ�)
ܳ��]�m(�^�[�>��L�osT�x�����I���~�9}2
,�">�$�/���l�&{����,⛜�'�G��{P� U����\�q�o�73�8��\�y�w����U���h4<GU�:(vu8��;�|g&-=�I� ��O' MnPĊ�;�Q���=	v-j}L�'B����g�?�������HDmv�(�_��;��h��۱��߿��1}0n ���ڞh�u ^�3]���s��d�=zF��s�=7��wL�x�3a�ղ���Aj�e<M'��z�L����rQ���X޹xU�+��y_�%���k7t���]�E�AcDT�"� �Ǐ�B:��gO%��QG|~~Z������0������&���믝���nI�k_��+��!h�!��{�G���K;�����DBg���H�־��[����/�P
���vA3�Dja?�S�U$�"P���n�	�s}E�I��@�AUa �b6�D�t�?d�c�Ӽ�    IDAT�tB2���2�3���}�'��9���2S���ȃ��ͥI���Ca4��)P�ށ��AF$e��Z�����#���s��a,���_��� ~f��g�MM�'�j�ZI#���e�q�E�uנLyb4H��j���"��<�m,tK�@�lش^����@�<I7�ܦ��7�i�������x,=���<xyvŭ6�	N���Wo���X��MT')7+O��Z+�ޥ˽'����I�&�ۼ,Ui>�A�ϣƮ��?���<kB���Q0�>��[m��Jq�G=XT�'��p
*B
�Q0��H�&,�� ����eq�,��"e��8*�F'a`���q�����n��6[w���N6޷M��9���T���P�R������ؑ�r��iz� ͈4��Ra:X�Ep���a^�>��.�J"�ݿ/_=|D�	��;�:
b���%�����u23��u��������7�S]��s��V-�oݑ�R%d�0�� @�x�	��O�I�R��d��!gU	�c�4��l^����lL�;���+��CN�r���r��{{_��F��[*����u�	�F �f�w��O���KW��^���������dc_��˫���� g�]��k�Fn#``���?�n��Md�RW�� �?�\tn��ΏNښDL:�=Z�?���S��AL­�f���׬D�SR���_�� �kh����%�]^���|�j���рk�^�LЉ�6Y7���8�Q�Uc4�aO���D1kI#��C-�&�t�*4���$�#���^����f- o�÷{������}6]��h� ���d;���} j��y��������z�[�4�e�I0�"�QG��?�l���叧� ĺ}祉v�.�kc����v��}�Շ���8����z�:zx�X��`J�ټ�,���o˻���W�E�6A��5e�V��m���u�N��#U-b-�����c��߻s� ��}aa�4��μ���|� >o��WN˹WOS9��b�\#'+2��2�n�β|t�G1� W�Ws�������3����裏䭟����R�̀�^(��|)�ؒ
�!��L�5���1wY�W�8f�sן�����<�4���xF��6��4l�o�����@M̨�	�i�h��lj+2���Z�� !le��}+P���Ij�R�?J2i �������s?��b/�����4r�����L�L}*4/��Ǎ ��x��>x[�m�͗,ţ����)쪩�Љ���C �m�V엎\^�OU��a��a�Y������i`D]�E�����h"�N��Lëp@�Ӽ 3A������F[�H�K���Twk4�E@�q��J���7�vN�vF���w�B�����k�7�=�v �!���k���a��FBw�]O�27��Q%�����'��\�b��h�F�<�z��\Sr
�5CB3&�d�k�1��9K&Ie�`vm�-�I�p��UxhQ�<~BN�8&O?���RE����� !J����{�r8i�rQ�y6o�${��y�y�#���%'���E:-�#Ì��b~
]�Lg	�al���c�u�Vٹk�G�?�Kׯ�iu�U� 3����q�KG*! ��q���R �G����h�\Hv����0�) �����j�:��X$�FL�����ء>��M��Τi+h���d1��Wd~�PՔ����:vL���.���K�eb��������A���ʆ�e3���$�AF��va��>@�+Pe��@6.̴%= �yIG@m��г�*Tp0@n6�5L5"��!�a�I�3�~5 ��W���1 C����/��/�懲\�s����� �+%�1 �8�T��z��p-m
�@Jj��e0��4��+1�]2q_� K�IŤ���te�����)�7o�(4�dSt���5��=-�O�`��{&����3����~�:z>���}Q`�G����\���_�=�����*[V�>���=�`�3b׎��Ql�^���c}��SV�gM�7��Q�#��kŮ�1�����}Bn����{e��&d�L� �ʇ��{W��j5.5������\YB��q��C������0��#�"VPh���X&��95��,-γ�{����/>�/�JQN�8.�����K.��H��7���m�j�w���I�z]��\_KF�_K>�(�q�YD����OɁ_\^���XL���`�d�3������ ���.�� ���Y� ړ����FW쏢��Zf�d$�"��>p��p6%��sK+�F�bef��Qѩ�ű� 7٨k�HHf�xp )Y^)�������M��ؙ�~�Ŭ�at����f�w����MO��������c�եeN( x��w?6 -�kN��@ܭd��0���6h ���LF�褙N��� �IW@�ND�F8����
'�QA��аPG[A���Z�F���"f.�
��@����:&uHаU5�Ku�E��w�l���7��uD�N�V�h�
\�NXyC$�E.l�ٱ�Mړ۲��7Q�FGw=^�����C���E��y�f�bv��v�����:f|&���!O�q�1vܶF\��*���B�,���t|R&���Q���o���-��*�'u�^d�
�E�o�NyO_7�Àb�'cOY% �� �.?N�����B�y��+Eh�ڷ_6���׮�ŋ�3ڀ9�Mњ�`�b�#\�ըlB���@�Fc�������233'?��������xHN"	
~�1��H�P�`0���ѣG���7%��˵��W����-��9-8��'�2�� }Sz�y)/��³	��9e�j
f�s �7�"�&���@�n9��-��E��@�5P�qu"�FCu\�5T"�V��B�$�".�p�%�Kw!'G����̌\~�=>g�z��*{�o������>�6j�D�R&���AM��QA=֭(��J�~��6L��Yր�E�����������������:�2�崺5h 	�a'H��/?���ɻR��d�#RM���dzv���K��L�������~�7��AmsTC1.1�ޝ:� �g��bV4ͪJ
]��1)�3�ϥ���I6rڱu�lۼ���!#���^�b��-�e�G�sNw�}��fwy�W������f?��̾�{Vd��=��v=�<���z��v��Ι�{���Q�����c���9J�|��m�����H:��k���5�8X�ǵ�5o?����L�����  �1���Y���<��Kr���x�C�J� �KdU1��^�
�.
�����ݾ�p���եR^a+2EG�l2&>�'c��BE*��W���^���.��t*&�㒌7e��=���S�i���� ���|�F�e�F�(:�jX"�I/��l|�C�??�;:_�9�u��s����7�?���eo�jL��]g�u�3vP��1bE'P��&�/�9�(����;U3�ۧ ��x�|�-
���fo9��V���4�k�\�'�23�,+�ʽ�����ؙo�b����J��cM ��?���/�����ɳ�3S�<�geu%����oT�8W ���	�\d���"4���[ .o6�K:gB0ix<*��șEWVT��5�U.�n�@ (38Xt ��ȶ�Y�17 �I�Q��x̌�q�&�C���|)GB���� .���
|��u�D�Nk0��W��:(�s@�7~�Gj���}#��k~�a0Ȣf`�f:�d"�+:G T�AsiI�v-��:}W���28c�Xtƶ�d�C:���܈����,.�XD�p�A �<�����F:��	���K_O��8v����>��{��޾�ܿ�׾s�n} x� �>}J# ���ǎ!�0*
�$��t
��ݟqݠ:]�7���+o��d�)	p��'R��ƴ��Sg��k�ҩx�����'���w��Hw_/A����o���@/�/ʋ�Y\XІRM�cǎ���o��~㦼w銔�U�4�ROf�J���/;:��	����T�e��#�hw��/�ǭu�F�9�A���/-�d�7I��M-h����oK�E�!�`�ږ&B#��6Dh��O�e�έ��S�ّ��ߖ��~*�SS� ����gO���$)G�e ��Ҭ�fa���)�06�N��ٱ �Ev�`n:�^�8�
�rx>��dM�$�/�6X�DjD}��� RuD����/���r��'r��-�TN�6n�t��䔬BwM� B8�I�Mp��R�����a3:���5xX�ef������`@=Xo(��g��Ύ������+ <�0�w%�� �s$;��)ٳ0�b����3o����m�6�{e4�u �3pk{C�xv7�(=�e���o��/�@�agK�m�#�6�������.c���eAm�l����h�����}� <�k4"�\*�B���2��A)|1���7>�
����Z��2�� 8yJ+�F��SD��ߠ$�JQ6�"�G��g����_��U՗�1 �QQȊ��s3�I�e��]�ꙓ�a��$��o 4?C��%��x{�V�i�3:_�5��8 x�TRuF�5<�܌�3� �7Ԥ��Y�Ձr�3הI�b���Q֪��zv�ѱA����	�$���N�6>�ug�6 �dc�z ��_[� �T�302�[GO��v,�2D���� �����OL�O�����WV���-�Veea>X��e��ź�µ�n� �VR��5� ��E��y�'����:�����3��%lPJ�FS�~�[�4<v]�v�v��3CΓ:.T"S�����fT�2RWA�&�ɐA��R��i{#�Ĩ>x�p�,�� 2jģ��R��c܌\x��������i� _���$m#!����F�ю����u@�&����4�&���I����H��,,����@Q4P�*�'
�� ^�dO%etd��v���!����C��6o�B������ƍ��=~�jGP���O�S�Ko� ������bi�����ƵK���1��e��i����,/.��BW'��u�.�|űQ��s=z�D�ONpt��С@�h�Ŕ$3iٴm�lٲ������r��Mj�c� `A���o�]��!<��Tq�&�J�iB7>#�BA��<x%lٲ��LLI�T������4�!-��T�i��IMRz��-v�v�:޶��y�O6���Q�~�c�X4�2�52��%�O�����9�ӧ����;2��1M��.w��\F��q����]� s�<����mh��D�.��d�έC�5�$��Ŝ��xݸ��Q������v5��X
�<X$��̬|����O���̼4I绥Xk�*x�.C@@�gD�(��>�yo���Y�[i���� ��޷��b��͐��$$���f����>v.��\6.�ٚ~떍�ljYhL�D7�Љ��@��a޿+�����8�g}���a�Gk�����c�`�?��Y���g;�xӮ��D�k�m�F���5���>����>�|v�>u���qm���Ԟ���|ʾg�Y�ɾk�|�A'0�/��<�X�L�-���C�z"#B�ՄR��B�G��3���;��<d���P��$�JQ6����d>C �٧�(� N;2O�e �=�]���!s��tL��'g_9E�8 <��ډ����'z�}7�7i]��F�"��6�0L۾G��^�iԲ@ \�P�q�O�(�e�B�1�7�@��c� [����p�:U�`m3kf���v��(�=�*Z^�Q$�{����~�c�����S23�$+�ʭ�������3�lMۿ�&���?��3�sӿ�0=w�T\�j�,�K2�b*X�f���N� ����Y--)����#�=J���&� z�.�n��r�&R�*M�7SOa�nxF��!C�V65�]��Xy���O�ޛ�@���kX�V�,xLP�RUta��((3 k�+���C�������lhCߡ2�. �k����J|O3H�+�Ƙ����%p<z{{y> |�6�8P<���h
��q4�c[9P_�(��+� �Y)�TZ�T(������ 6lp���d�iY�nDΜ~E6o�$�c��{��#�~��q���K��Ё:}�4�EAG�իW�>�Xf$�MK.�f��@��<zTvn�"�.�\�߽+�ݻw��3==%�Ϟ��S��d�ƍ<Ɠgc��㸥b������,�#_��ò}�V�|��@EeǮ��g;
�����?~Kn߾MM[����G���/�� ��eD�k*W �#�LK�$Ց�FF#��\׊��21!�Ւ�`��1��
�/��3�C�S|������?S���M	���"�Ŵ�Mҍ���$��V(�V{"ސ�����e��-���|(�>�+>�� <3�ά�2��"jK#p��"���F5��:��D`N6�V���N�mE�&�91�\�5����bh�]J�:���qѨ�Nn�3*:`8�Y�3w3�.&��G����"K��IRj�4ƒlx�	dǟ>��[Q*8�-E���֨>��
��AQhp�@@�k��B,z'���q��g��3��G:��\J֏ʞ��e疭*;ɺ�;.�M$�� ��}����lbD�|��(EŦ�9
~6�����U������p?6�k�g��'a�}�>g������?k{��z���,-Ck��6&8������(�E�������3` �~�5F��� �s8`�< |*�!��K�F�kq��QĊ~#I��\{
�U������dI����{1����R+��u�T�����M���m�k2���+ԃ�{ 𝹴L���];t� #� �X�ǈ��l������ >jw�y�<�v��%����__���Q��K7h�"ߜ.�{��a�}�b�&�6׈#�z#�.��xV_,%�d4 l�sѹ�ɐ�hk�e�r{)�T�p2��� �S�i��2;�,���Ս�w��}��_i7��^[��/__�����م���
` ������kE.�Gt�b��m��꩹F&X,n�`<�U$�����cQ`��b�D!׈.��d	�M��Z��g�&7{�?k(dQ*M��0�T�3�F�u<�����`�J� rBkAk���\'���;O��$3��F�L#�e��u�Fd�V-{��4��}6�	�H�	�o��Ό��m��� D�)i�Ti�����gs+�
�c�*冪�Q}�+�P3!]���?,�xZ�V�ʙs*$��a��U�Oed���r��3�e�&{�H~�wK����I5ٿ?��W�]c��ĉ��������? xV'�F� (��߽CΜ:%�C���^�>y$��{E�l�,_}���;�ˋth��eGd���d�۰^VWK���S���s���ДM�S��ܰqT^�5Fዕ"��F7m�m�wIgO�<|�L��?��7o�Ԯ��Ç��k穵{�ڇr��U���f}\���PiIvvI�3/�tJ��#��rI��/IE�"���72I�������b�P��
�8O]c0�{/x�a�g�X�S8�&�X�� �)�քBCSF����e������+���O�ʋ�cĚU�V�*5�dJA<���
$ֽ����s
h7pL)O'3l ��*��
���9�)����!:r~�/�8ֆx��}@��+�Y)��憈�(�}�5̠��F�as�V+21��k����5ġ��a �w�.��P������k��7�c����w���;lA��&�1l)���U���O�ٔ����{v����9O�Y�rl����m��� ��O���u/���Q�Y0��$;�u�mu$ر};j`#
�9+]m����[msG��x-����m��~>��蚎�n���6�B�̏{�����m��-�d�8����#r�c�l(� ��|�L�-�p�&|tJ�(�w��% �ڵ�R��)�Hp>�CM	x����֍����[t<c��-*�    IDATk�5����Td>�$������μ�ݽ� A)�H0�hd�B��@��롢�gH�l���=J��t�9j� v� ީ��3&b�7�֋�s�����d@��]�)ǩS�@�GIT<����D���^�b`��5�]����Oz�C�E�"�!G�h� _�T�ٵ��?۶����� �O�����<�phn�<�,��f��7 n@���owQ ��)E{��8�V��� ���'��Q:)]�.�+Z)�X�P!���i?U�|���j�'٩U�3����NJ1a�>�B��ƴb�g�p m�K��,�c������'����) ��� 7Tņ1�9��b�i/�����tu�Q�Lj��1�,��u@��'�:�Y�Ӣ-�(�oP��pS��=6t�������8;<��ܹs'uP@�]��y�ok�D'O)$�8�l`T���SR0�|gϰ�"��E~�~h�u�w�}��?�Q���l�?E ���{ﲠtǎr��iٱ{����;���P���!�����o ���S尻H2%]�N9���>~D��H*ސ��w#_}�����y9rh�<|�P�gg��5��o3S3r��'��d`h�Q�g�'	�>�J.^�(gΜ�����kl����+�8ҋ����u7Kwߐ<���g���;AG�C��ʫ��cQ�����K�)ݥr��ťQ�KY��NIuuJ-�d�"�����f礶��L,2YMDB+����u���aD��U�xr�f�|�H�z�Tg +��o�A�FٚD��4 �:G˒L��g_YY��7l�-[���-;�t���\��X�7=>>���0���5���k>Ȃ��U>ڭ���Y�ǸB=d�6�~����ZP.��i۰�c�v-,����w&"�1 	���g�-���f���{�Yg�"�TZ)D�euA�!�x+�������[����w�V� (@׿ha�J�;�+�� @�qG��N�,�sp>��u��g�vٶu3;�*g��Y��H���=+
���`����m���m�Ou�=��C�	;�Z�d�5���mO0 ��a�7�n������^�~k�c�ѿ�(�q�z��Qw�����q�����˲h>��s�C��(���g=O:/��r��'r�ÛR�'౫�B���������R�jX�Y
�<� |�� <���Ɂ����Gׯ��O�!�[\]�\:-#�}Rȥ�Z\�S���)���W_;My�&��*!	%���ޑ�1a_�5c��z�|�l�??�=;����3��{���e+X}L�'+j=-\�S�;�H��9{�y5�-:�~��aL���X�k)��E�bG� x��i ��w]A�dA`!ڹ��z�R�����ֆ�{?o{�6/�́��������[��;49�t%D��������hJ��ED|h��Mc���� ���?;:%��^(��@C{By"�u�G�������#YX\&����}�z�<��۷�ޝ;��#+�H6�M���;(���`�*�D��" ����������G�UH{�+�.�7��͊4{�F:G�Zb�?�fn����;�˦��T�僆��D�Z
8�ZL�@ۢ*FW1�B�Y���s�Q�r!�MF�d8Ͱ�D�]��ǘo޼Y���K���1���J���f\@�سI��]�6��N����q�2@�<F��\�_Ju���"��V��L#���b3��3Z���\�ECr��)پy3�FP0��bWT���/�.�m���w�#������'?Q��Qg�ú�ٹ}�ܻ������9�������ț���7޼ ���R\Y���N��u���2�|��.��g�2�a�|��r��e�'��k���-?��H��_�'�e�&����*���륻P�O���}_�~z_J��$Si9x䨜}�e�]�!\�,hT�EI� �C�
�tw�TS	)C�;�<������,�RE՗Ri���b�W f�o '�\X��P׾�o�h7���H�QF^���u�'��*,	㫑_�Ouj�B�Z+J�VfFst�gPzzI��z0L�X�u�L�h��I���W�>Ha���vY��H�^��h�x[��O�kT>�>�r��"l&b�k�9~����4�6�%�s�C�tU?}&�jM�5�X�v���ֱ�|R��5O�G��[�F3utl4;j!�F]�;#W̎�O��a�7�tW!�^ ��gэ5���>ٵc�lވ"V�_�\z���3�+8���(��I�/{�ZC���$�m{��}��G���nG����P�����@Y��h��ua ���6�Ԯ���h6���?���XT��e�ܸ�Qy���㏧��Ҍ���vMV@�)dt�<N@�O��X�|tK*͔ ���>��J�ۈ���-�[R���"�}=rh�^��o^�O��e���ϟI�X���n��� g*4]y9|��@����f���P^����^]�,@~���N����R��ڙe�jT�!��	L�@[�mn7�M|��a��d�_�\[�/�*�j�t�(�=Pʲ�G�ak_sD��u�7�A�Bxͺ�A��+�[cV�e�D��& |�X�����G��u[�>j��_�ǚO����_����_fg^����+��,P�bvz��jE1J�P�Ư��>p�d��S^� @�eWWe*"F���$���������'�ȋ�����G���'��ݻ2;;O�.@x�l0TQU���n9q쐜<zDz;�T�Hƕg���1��A�HJ������/f�ڵ��ƭ;To�uvK�ѠbJ"�S�~W �)�6��y�P�)kt��F1i!��o�qA~��)t�	�K� bڨj��j%P�1^1'M�D��d�x�$�C�\&��g�(�)����3�++��1q<j�;��: p��	�oD-;;
�˩z�r]4 �_�~$���#���uy�x��E�k
�ߺ���E���<���L����@��}�t��j!U�s	��JY2����k���ÖKƤ��@��ё�R�"��|L����cٵk���:�t�2�5���X;rTN�<.�dB�=d���=;��H|��\8N�x�,����C����,M���R���|Vn~t[F7n oj88?2�������ax�M�+�\����!�j����e��ٗ����%���^c��������	�Q���������w��LH���1�E�X��Ғ��W'���� Liq7x���c�:��sѹeT̈́�O�1 ���TJ�� mJ�p��Ju��H�W�ڤi�%�B�n�屎꒎����	pD��.��]�����Fh�0�m��y�1�xR�6|�N�mƀu�x�KL��2������M_%�8�&=k�4��`��#<Y��@큝U�:���5� "�Z,Kww��˴c�;(��-��&�����9�!F����%l�5�a+��T�A��|:%���twvH:��l&AIɡ�ٱm3;#���K��R��wm��"�=��(�����=_k����2��`cۢ��}�jch���Z| o�� �J�*��-�2�X�Ό۸�#�_[@!m#�ic�,����qL�^���=;�'��}�6Є��4>�{Ǐ9��7��J�� >�@��X<%3r��;r�;R�b3A���S4Q�\�뾌5��P&��O�U���	��@�|v��|��g�Y�|6#����������ӓ���-�)��JqU��D��!x6PO���,N�����z o8� <m����3��u2����Ja�3r�|��Y��"Oˠ�ll�������S����y�D\�~j�l/�ě���f��ud��,��̠��hX#=�P{ir[S�� ��>��!c ��-,�K��_8~�7n���jK�>�f������==?�_�L��
�F(�/���(6AF�6���ZtǊ������y/x�P�*�Ά�pp����X#��Lh�v��Siɡ�c2-ݽ�� X�ك�����l�(���J�!�'&dii�W�����b�D62��-^;+��D�$�ʊd��V�9Hxǂ�*TP���,�*r�ڇ��e~a��	�:�/U�l�Å��*v ��J%Y]Y��GH^3��U�Rˉ���W��Mٽc+���	#-���+�0�	����pF�\4	�@��I��9F�A1@q*�y�������#��G֑�Я5uIe3_�hpQ�]�N3�Ð�r��4�ƛ��Lge�R�[���ū��Լԩ��m��JV?��?�����W��"��x�X��q�ut�Y�c`��	{|��yY?2"�DC&��ɺ�Q��钇��266&S����[ߒ��y��E��L#m��G�^Og^�^�@>�wO�nX'o^8'���-{�H~嗿�Ͻ���ƄFMEP��RoʕUy��sfk::;	����P�l�Ƶ4>>A#�놌���Rz��+��/dq�H�V�������I�����'�?�2��dd߁Cr��Y����߿(W���<��H&rW6����vH���&2?�� ���w�ѐ��@�T��U�xk�������ȁ� �Dޙ<�̈́�4�v�K������D�Xo�������ـ��|(N=gt��q��t ����I:F�i|E������]U�!����F����t��� tQ)C#�|NO ���J���#P�o��d�-��c" �mBP�`n�hn���:�9U�n�g@��H���3G�<�$��4c6l��M�yt�6���~=����� )m��QX � ��,Blj{��u_���uQ�CT�􁄽o�����H��"��9�A��lʢ��c�<o��{��Ʈ�>��H�-a�
f�X���y?zO�t(�#�k���ǿn?_n�Y _��֊���Q=��-�L�/��kɍ�w��LH	6#�.��\�~LX.��/�wG˃J]������߻W�o�TjqeQ����LOʝ�n�����!�N�n�M��S�NIOWA��*�>l�k�r�# �l�I-� J�R���lk ��yNX�Y �pZo�X%��3�����"�=&{���jv��]�_�i8In_j׻]_�xGpm�©5b���%&W���e^�yz�Cb׿��z���P!�C�L3H2;���Jf���ɣ�����_d;�u���l&�~�/���s/�����G����2�2&PT��M�6k��&YM���PoA��Fvt��Ԩ�a���.R���;'�z6
�-;Pn��V%�ir�=\��BA���%��I	 |�l^&^L���2	��:0�f�"�f]6�˹�'����oJG�A _YY �E�0��Yj�C9��՚�{W��ū7dvn��l�R�Hg<�2�'��K��&����%�$x��sZ��Ւ���Ϟ�3'�K&�
y��bGW-�Ө$�kH�6R�c��q���C����`�QP����KX0~��3��,p[\���e�l����$I��\_:���z�B�>�ԁ�L�Rk��JI��ɵ�����ϥ�j#&*�('��\��^2*��g�ФT�/�P�|�@<�C�nhP޸�l��O����'w*4��ܼuKnݼI�'O�d��? �Fat�9��I9}��L�?�����db�;�_���7坟�� ���W��3�����Դ,��K&�e�svvJ�|�������;}�tL�l�NSiuUf O���ɖM���ezv�kd`�z޸I�LN�O�~W>��s�4D2�9|츜=sN:::坷.��\�ڪ�#C��*��[e>/�t��&#d��ЯE��T\e��f�T��9��	w����3�m�"�3�q[ˠ���8��>]�(8ן�h����U ���#���ń��Z�iE�x^z>}�/b��0��Z��>!��V|�2�@�)bP�h'�Йe6_n�D��$ĵ���$ox�����>��?�7#�ȭ���|�5ӫҾ�.r�;
9ɤ��(sٔ�����ɖ�Q~�R�����?zK����q��H���L�>�7�O	a�׫M���"߁�A��(�6pu�5�SM,������ �T��Z��[.Y��5��|���_�
ft�E���9bߏ^S�yd��{�3Q�,
�m��9�I�Ş��=׈��>��{>2��]�!7�|� ^J2	d�\��9��9O�>��G� ��8�4Y��6|x@rY�W@ �*3�����;�0�B�Uv�F���#/�C�X8�� ���"h���U�}AC)d�\�6{�8�.^��l�O��&�0y������|�H48���t��-�w�Q�t}�*_ �*@Z�`Y��{/:_B��C�}��[[
�ǲ"Z�F�=�M����e�A���ֆO��s!�|��f�!���\�ߟ<x��uo�8���l}���|�f��W��ͧ/^��d"�eb�����H�Vg�;] �
�U�9�p(5Դx�ؽxq�[&6yi ���:�D5Z�%�c�4O�Ǥ�p �B����I�G�Ťq�C�š�� `E�h�J�R��fU�%�0�/��:!g��~��J+�%V+1UG
��V�TA�'��baE�~��ܺ��,-�jQ *��9ݘ�!��x"��j�(��ev`K���O ��V$V�Ȯ�[��_�c�(妴̸"���$�E�p�@-5�Z�*��Ŀ���r��l^�H5���T��(��a�L���P�FB�dV�x���K�4|���=�������JO����1y��ܼsW�~�@�_�H,�)�@�wp��0 O�~F���1˝G �E�� �	�����PI^�*��|���>�K������oʞ={X��֏"=�����<޿s���?�}�_�Q�x��?|Dn\�.������ gN��o��y�'/��z(��֛r��!:Cs3�2�tL���X��q�YYY��W/�ݻ�P�p�tf9�೤�'���7�n`���۶�ٌ?.�LF6m�.�[���÷ޖ���i�j=&G����g^�\�C�y��r��U>d��5���qn�F&)	�Ul�C�JB�Ot|��]�rqE���UK����+h�����&�χ�3����(]k��+d�D�{0��2 ��X�F�v�MP�f�� qn>���"S v�*A#9y���V OHd:��mؑy�����L��?/�_KQ�e:�i4��ǌ ,�l�({���'c���(�tkL.��x/N�K��Զ�ԏ�^S�䥿���g�i�ʧd��K6�ɦ�f8�EJ�s��X�r������TS����~���W�����]p�~���������9�f��6��שq{���DyB�����욣�)-5��v�>�c��uΞ��v�����E{����{����������5d��.jb�9d'Y͞H���iy��5���K�I(�A��8ԁ�𰦾�k <��7�;(��̗4*Y0^ag�ŹI�ju��
�|�o�W�?F �-���F�,Y��H��T)uZU{ݤv񺒊�s2blE#�6�Ƚ�Q;�>ֵ�E�q^��`d� 1�_o��y9p�S:N�{��N��^���f�-��߇?�}��)��"#z]��:'��s�X~�a�&�h�ؐť��L�;|��������O[ ����}��>��ҙ�f����KR]Y"�A�%$w�L)% ��NS��܅��;��ۂ�j]���^��o��`&PU���(�e;$�5,�ɓKUhj"Z}ptYej��l_��Sƴ	S\*�n�%o��}��[��*[F���8#�FEz�03E�Hg��v�)v�KR�?�����269GDp�A��"����IԤ�+"�rIJ����7@9�b{YY\d��#�ɛ���P7���p�}`�ZF< f� ��a�qt�t�dXn@���(�������kJ<a�`�2����q���E &o�Ҡ�COO�n�Lp/�ܮ���P+�%�`Hr��2�b�i�[�|*��3l��LX(�E6���-��nv��s�l����#<XW%8k�rԨQU���A��?�J|�>�s�<	͜@W���#���Q��Ghƃ;�{�^ٺq�|~��<�S��    IDATy���59w�|��w&��=|H>@~���q����23��Ų�v�$PG��[�dqyI�����¼E�?��es�~�(S��6�
�BMN>�l�C�o�B�����������Od$��ˑc'���I����r��U����c�3�X_��p��AaB!����G���Z���Q�B18�f@�4���P�s!_����eR}��T��1��Qh�=�3
�H.O��������/�U���3[�@`@����V� �MKs}-��s+O�̖���*���u$�G��@�qT!�|0�(}��.��Tl��Q �\?��8N�7�
��U��0��${۫�h��� ^=��Ш�R�T��*Q��H_�*:AV�����lR���qdP���	?�O`Y4�Ba]�Y�Km{Ѷ�,�r�5������9��>�H��u�~P&:���h΃9�~A�eS-��`;F���x�#���x�������}ٵ��8���;7���Nsb�I0�iM�`c-�n����1e4�R���@  ��Ĕ����r�. |�T�-�'�sN�@�%�,���斚[S��l�p\%\�^���kU��V���,I �Z����LJ���dx�W���-��lb�5�HY�Θ	�lk��z�0���&�!4����U�հ�H�aڮȎ��d�	��ٔ6ߤ?�T>�!��,��|��r=1��ozNqp�6�s5:o��z	�t/��n�q���Z^]��=������}!��(�6_a�� �\^Y�:����pttt���w!�ip���~�7>��U�-�dFb�:����Ab��Th��c�e�x����Z!��FA����sF��TL�h�� ʭB�I�'SR�tJ�R� �I꼣�A�F�:5��[��3�Mr���ˋ�ahHνr\��)�x]�29g�LB��2�6���TV&��ꭻ��;�\�3C��Š���(}H<i��4�8Eh	��5�R*0��)���RI�)��ȁ��m�6Hqy^*�IC����)Ɍ��,}e��`"����H�e �*�������QM������`5�Z�Z��C�ǫ�5h��"�,�Z��HS'��5���b�fW���/�x21)˕�� ^�y�3������B��Qڐ��F1��:Ϝ��Ɗ F�D��| *S���<8�z���h�b�ź ��l���M��"i�����+,�E�T�L*&��}E���y6r�q�2e�6m�H����(3��R.�d���xԀ@m�V��fI�������|���ӧ<6"4�X�n��Ks���t�$��)s++26>%��EI�PĜ��'N�����+r��ՠq�ld=I�5 n�3�b��� #�d��
k��-8�ŕe:��q3G�	&<°�uV�
�T�N�w�w`D�f-K�6��u+xj� ���#5>��@zkĴ�S��@F-Bmyis���x��>��)���l�-�f�� :خf�q_I��N:�
68����u���J/�F+�KE��n�~�/n�6:�O6 �m���&�RR@D��S�:s�K4e�� �׏���� ��3�M���Y���6u 9�GA���k�Ƶ[؏4G��~��G����5hTF�p,��b�Cv/6�������s�����o�~�
�Vs"�y�?o ��/�ۘ)MT�+ߙ��`�u�T�A�1V���D�,e7����2k��39i�3�tbF޿t� ^Ry)Av��M�P;;�GUC�Mx�WZ?Ȑ"Y�Z�a�N�\���Q�.ٸ��⼔�! � �X�b"��=�n�_^y�(k=@Y-����#�՛��)h��k6]�RP���VT��jm 2�u���*<n����r��}˄Z��e�PO�~|������!�ik�p�����^ƞ��@DL�K!� ��e�h���@��yx�~���`E��uq~b�L�R���J�AGw��x�����b�i��z���7���o��������Tilb�G¢�e�0�4���x���)0d�mj�:R�?Ms�USa#�9,X4���T$.+ ���GM��Hx��itr�ABJ��E��%Q�I!����G���}rp��F��������Gg��賉R@n��T�N-I-J������ZzЦK�J4��DM Fi\��ʢ��O�4h K�g��2��%���c��1-��z�H��v/���"]���8R�Â"�k�C[$ �L��H��#���/�d�-܃)� ħ�e����l����$�)*Ơ�E@�>,��<���b�)U(�4RK�Y7�"q��	 <��IB��d�@�$�� e��.cG�1��{���> ����V)Qu�-�q��z��p`�!�}����4��.q���5���|���~�|r�C�t�}y��!�;ʫ��dQ%B>97�f\VKeI��쬊�I/��r��6�r�<{���pp]�Ƴ�׭3��5G�\SP��1���#����C��]�rE._�A�TH�V�W�ј/T�a�4�A>K��Il��cc4�5�i�]hkB�L�=jϡ��z;lFU���I+ ��V���I�ЋWT��Q@G��>�{>�.�@Tp�>������'��ъ¨T��D�������y���ߜ�M�o!��U�Zח��H��c�s/�t3bÍV�!6lr�#�)Gi
���6vBK;P��d��C
�����=�7�HO��� @y-�T"�`���A����QN�#
.�[��c�q��u��6�Q��S�3E���$[)���9 v,�C�;њ?j]+�^s� ހp�d9 f���~�S-���q6U��8�4aT��b�|�Ǟ�9%�-��gl<}9�Օ%�Q���*����$29�����ܐ��>�z*'�
U�VyB�8X����,��q�x)~1cc�SW�B��.�S�p���� �,��%��E
�9�C����'e��]�h�s3����1 ����-Τqa�I%�Ź�8�ҭ#iB��}W��
���.�ʜ0� ;aM�j���;mE���~Fӟ?���7��]�F��N���x"��Rk�f�o/z`2ǨS�����8V1��ļ�-�����g�r�	(kvZc�@u���J �{�����=����/��Ϣ&���^�������g��f�Z�\�6�^��� >���y��Z�L�<]��
��!zi��4غ��8<�͟���E��� 9o|x������
)B�Scr���Fh\�0��e\GT5�2��T*�K�e�r��a*���Z'
h�'g�����g����$�,Xlt���i��¢=FWP�P��(`��A�S&�5�W��jԩ�sx�.9yd�lF�5hY�,�4��f3L?��[�LT�c�ql����DC� e�X��$�����ȫzC2)˨�o6I/��D�rn�����.���_��2��"_<z*�(O&�d	�2����B}"�׮vn|}���!ک6�0X���t��j���m��b1��2ښ��JE�#ʪ~T��}b�-jd�k��U�R�U$��Pn�Z^��e".���М8~Dgg��W����#�,�4�?^.��)�0v��L���GiquE������:�{�����<��^>����7HG.Cp�{�%�B���2�RM��d㦭����*������G��P��)�`C�v@=��Q�h@�4h����P8�m֪���>0����2�զXk�P������k񭠤5j=~��z�=E?����[��$�5@�k�y�����e]gS{�:ڦh)����t��|��5��M�.!R��͘ΘkF��s�"��j��2�Z���}�:�.�d�< ff^n��O�~M��ʬ�(t�pOAz�)�2�#;7��ўn��h��HA�qNh������e@�(8_���W�3��?�6"C{f�tߴ���w��G�������`�8v~ۯ�c�����[�sl ��Ӟ�]�eZ渋��g�vV�k��G�-���i�����>���'?ak�n��-�j�W*���x����ľ����iy�ڇ�����@��n��ހ�g*qt��� ԩ��QӜHk:<{mx����oeA*��R�����XK�쬽wU���ӷ�����n��̌3�q,��~_^"�-< ��A�<!񀄂(#��@B"�� )�@2���㙖���O��{�OU�����^u�9}۱[v�:�ֽ��:U�V������Z�9��G��������ݗ����LF��b=b��ȃ6�|1�� ��3�E�!�kV�1��[t��s0(/��g��6eJ��-@k>���m��M�am.fbq��}��ݶ��9��u�����&[=� d@�ahġ�<p_ǂDHֆ���!��U��9OG����N�44����ؠa����^=���Og������[��\�  �������7���&>�XE�-k��/�Bې��SϜ-'�
C.�.��
Cn(cQ�걈����>��RMѹ&Js%�PW�m�WT�@�X��s�4j����1��GvJ����=t��z�Qw��)��u�j��7�q�_��|]1�G;z$���l@B ���B��A; 0�[/����E�>,�17u�;�]�����ܙ݉{��E���wO^���g�n�LAꕺzg�SX.E����,l��<Z�ɉ��{{;|� �x���-5c@3A��Sl�� �3��*��uw���ǯ]s߿�����7Ǽ-'n�g��tGrs���w��M��#�I ?�}��!̦~��zV�Ar-i�	��!ݠ����=҃Ao���!��ŏ��)�թ�=��/>�>��U��Y�8�P��Z ın ��d���H2�sx�����7�r�0��Y�)Fw����g��d�J[��X�%����Sa����Mg��p�^{�M���|����/39ư��W�I-d5�A���bn
A�:UE �k�m���eMk'�5�Pu���_[��o������s��l�m��� ج~ӏI=�9#@c��m�7�I��pf7>-s�a dj��&����\r����<���M6�i}�Ƃm@_���1t��
�ؔ*Sah�`���H�>w��� ���n�����^��v�m�< �6.Y����r��C���|��=u鼻�8�-��s��/#��KD����s,p���)G��K�(����p؞$W�^۱��:k����o�
��g���C����W#e��XC�z��@�σ����q~F��͑D0�,��<��, kXX�s������&��5ֱ�����&�熏�jR�^������^��UWLv]:	 ��N��ɑ:}f����ǂ��+�:Ҡ�k�Αc�p]V;P~=��Ξu������?��{�G��*�B���YoYs�lzP�	�d,�C��@��J��a���AS<����\ �9�|��]�cÔND��>z��?�gh����Z������`;'{
�JH�lxh�H.���R�`TK�+��� G{Q����&�ob�ހ�g�F�9*�ɇ7M�OG{��x��_���*s��z���o��_z��k�z��˦s��u�
���c8 9�D�MV��LRH�����.�v�q��e��i'�)�]7 \�ᗅ�Ʌ��Y����'����g��w�Y	7�*�tR�-7Ɔ� �:��Z�GN��9x�� �#�tXv�7'c���kΆ)T5��Sz�l��U�t���JR=wE�r�w'��K��S�?�}�a��v�1A)���$־�h�ȫ|��RR�.Xyf��IH<C��Cg\����d��$Jxޙ/�۷�[���W_q7���Xyt���Q�dI�W�z˃�[R�_Fp�#�%�d�dʒ&�m�Ve�^S�dP�U"�z+�#�ylh"�/�����w��t{��;�7eU i�5����@�$�� �r�e��76�[wn�o��n޹�W߁&Ţ?}��{��w��üV������L%)�*�uPt<�6��뮿���s|H��+DҲ��+C=J>sp���U�{X'���G	=���C�Y�P�G�f�\��7��a�T(�K"GPoz���]�y�}����iU?Y� 	�k������3��IjƦgg����)�#�����qY�i��D�aάsF����I��5l��ڰD)C�^{��B�&\'�w{�9�4a }ή��F�+��?/��v�m�uΊ�.�Oݹݩ�|��>��Ew����|�&H�c>x����"z����}K��x��<&�u��;�k��۠����Z�ր�@^A��[�!��������z��{�^�$���)�T���]��=p��k�b;i$�;0�8�s��梍����{��U��G�MW�;{3W#q�`}�	b1e�����M����b5a�V=��F�z���K5P�� 5SU��gf+X���s1J��
�o���+���{�������s_�����i�d#��fr�L?CU����M��T=̖ʦ��C䊍��@5> �ܸϋ�rgTO�
+�}N�����Hyg��rP��
��@ޢ�^��s���Ca�l?O��s"7R����^?���d�J>��:7"��Ǯ:�ᬥ��n>�J}�Q�GAKM>,�^(���Ǟ����ހ�-�yҟ�����^z��?Z��gMt�E�ںcx�4r	�BKI��(�sLO�N��XyR�΍���+��6p�&ݼ���Ƥe��[ˤ�-��$���ɁF9�f��5xťG�����Be��ܝ��ԡb� x�� �V|�t���pb�Uh��u����n��s�Й�Lz X�FErUj]���K����]�p�]8}ڝ�;��g;�� �;͟�PFp�C���� r�A�/����z�ɥ3��ze��[����sw�h�n�s��9tw�Kw�p������F�^@�j²�؀{@�Q}��߿�P�ܤ�#�1�ߚDCfx��֓I��i�+�0�P�t���Zщ�ʍ�<�:�u��r"(7&&UJ��b�X�� �*$�82nOn!7���Ac@q@)���ل%�`�Vv��"�-�EE�z�0��0��Q��,���S���o�Yp�X�̮ϕ ��rT�Q��Iں��_�EՐ���2�a�Ƭ�"��+P��$��k�
�,�*��rY�2��'�U��|[�V4鲧9�n~'%uJ�g�ڊ������d�<Q�9�:N��5EF�>��7]���eT�Iz�N]��vi�؛�K��u�(;���C�;Ϟ�7���si}*u�7߳��7�M���[��?7b{��-0�ݰ�e���sWΟ������M�0 #�0���B=Q栬D䎟�1C�m�5T��6?�m���N�J������k� Q��,�d=���Y��b�[{7�����d�����ͽW������j�,�ݷ��uTM���۫�FUld��_/q\c�Nu�bD��g�r�/��m��W_g�G �.����a�X&�}�z�vi�D��1���sę�2��Z�,�\�ڕ����U��M���~�i��'�qJ#1x��ԫ��G�V)�-7���(���Ξ
�oa��E��J���ܟ'��@��e]#�袶>���:�Nψ�B�����#w�{�~E��=��ط�ޞs��i����c�w*oq0n:6=���݄�6J��ٮ�7�o������[\w�Q��6�m�Gm��l�tE5~9����ί�?��I����{0�������q�����#$�-����� �Bp!2�G��m���(PAn	��4�d� |OqЅ�]]a����k�6�
�pU�~o? 
�J4w~ń�w��wࠁ���;���ab��{��R�]*i�����X#�Ti<� �wH����(%���(WY{� ��O� ɴq�&�w���۟���l����ng:q�1<�#��H1#�}#I��� �YXƅ	�nvcP����1���>>$`�s|�V+�D���,�hB�;T~n�Z�xr9�,Sz1s���lgʍ��s5�E��z��"k���)�K�Xeч�rXS65��a)T�j@9��tx�X�e5�T3����#��铳r��` �    IDATpu�D;�g�f9�Q���U2EM�X��B��K}V
b�Gx.l�o{�M�f�k.4�"��k^ #
���>'^/?�l0T
��$Ei9�*.v	U���N����H���=�1�F���1 `q"H�[hB�%x����f�Ai��,��uҒ5�N~
�k�OCQ ���B�?G��G ���۪�u�^_��5�rP0jD��So^��p?h��^n٢�� RηN&&%[% �b�#wz\��ΝqO?���g�`9�Yȃ��@KT��xK#���(T�����w��3GV����u�[ �cR����I�G���x�N��Q�ci'��5
�9�l�Q�����=�V���q)��V�QJ��7��瑽wg����<��s��&�����gcFh�t�����o�?�/�_{åj�bQ�������G������B\r�֟*5���ۅf&@W/� �GcIx�O�Lܙ�=w�3nAi��y��y7I�>�t%�F`�s��������?�}nЪo�ɪ9�t�jC8��~�~@ْ�"#��=8�&�]�ZI��r#U��z�]9j��GҝM1IvX�<(��f�ڣ��~oժ�{�x��eN������	z�շ2��/.`���(a��s�#�mM�^�'���ϟ�%��M�@����������;�p�?9o��j	n x?ʉ��������iR�4�#)�y��7�.{��g6����l��S6A�,����iⶵ��ެ�; �6J+!E���3j��N� =�1������U��WK�,�c��U�qI"!Q���&h�&�![9�FltJ"�1���M=��W�pR�H��"`��\�/s�6q�:��C��� �	X�LT��  `�
D��y�"pG=qH���!'$�>>@%��#��\@%�<?�툋��םV��M�g4\��G� j�IԈ�[��[��A���0�h��A�Ftѣ�2�6�K��DF�s]���y�ǳ�����������N�D2����R���M�S��ڣ�F��B�]"��J�Uօ�hCn�� (M|h.]s�#�'UuN
��4P�c��e�T�@��y�7޽��Mn)x��M�%��h���C��ds-!�����W�����l��F��R��� �y�@ɺ�=����J�t=�MO
�N��)=xn�Eq�Z�d�>Q@��I�e�ξ�'��>��}?�o�l�H�v�����}[~"���}�R�V;�<e"���V䌒��X��ˌ���f�/gr�.��%�&��QA��ҍ#��
�}�?�t1����(�����̃��UpNA�{c=Jw��Z0W�,a���b�AЁ��@*����We� �O#�ii�ýؿ�윻��$������DK7\<�����"�'��Y0��B��!:Xy��}��U,c����E�H�x���s�!_X9>>��x�O��Ȉ�hv�eҚ�V��N�|�c]*�J-m�$��H�Vo�����~����� �?SP���>�(��Ȟj$Ot���ڋ�� ��M9��Z��w�"�{W�4����w��e�P���Q&���["Ͼ+'c*�4|�<�X+*AP���T^�����ҷy_[�����:�#�'��|���X���}п�Y��E��`�1Yz5�d�a�/ O�C�Y�\tr0]�#�t]�ַ���w`�bM0�)[64>k �ynE��)�B;�jqx��8=ᆺ^J��N�;]����ѩv߽��_+/��0T�S�X�')cn�\V����~g©UV�G,��Vy���۰{k�����*�lw�}~�� f�6̺���ř @,=̛;V�P��	�6�}|�Q#$���⛫�.�6hL�-
Mo=����i�7�^B�5��-IZ'4[bց�+Y����K*��i�wL�Ϸ*i��������<+R'ӰU�¤{
�k���x�@͝~jNҧ�������x�>��ɳY!������5X �úX�r�f��!��{c��%L �2����k���g9 �s��9uP����"�1��Y0�gG�Y��ܴ�<,��� �f��\�ۺp�G�d}�}��Q��"\�]�C��&�dEq�i���@
���rJ(Ɣc���T�٩����	���G�&�#Co>g��.QU������	�N�sIgV;q�����v�_R��@ZW��a��/|ܤ�l�f��.�o���M��er0��/Le]<hƞD���8��`wr��]�7�<��]�0� n]+z6���;W����#��]��'�	a}�~����ǵ?f�ZSC���җ7���^V�sS���R]z˛l��t�ʰ\�ڊn"�2(=�|��?mxgگy��I	m9!fM2ĕ�:��6')jT���U��(�{�Tx[~�(ȝ��<��(�L>�%){�� � !����Z?	��6J@�T�9/$V���ʝ���O��T����|Q�fG�\tY��0���QW��U��ŪI�dB�6��ML�Lؙ,\?�|֋�@_��e�'���V�g,5n1Yi^���G�.:ȇ<*�3�gw�-&�#�r�P�%���T qq&�>�v��`[���&z�f@� ~�� ���ɽo�v�=,Lx��}�p�n��%�jH	)-����A�~�A������%$z�a�]��r�4��l�������&R��$h����dIK��&=���y���|�����2�	7^1i��N��4V�t|q�j�ߞH(�)��9�
����f��ڪɣ`R|�J][��K\�_�K����XHޘY\�m��4j�a�"H�<��_V��W�¦g��>!��G�M�^Vƫ~�9~���w���sO3���������Ez���>K�sa�X��۞�����蝦�˻1��Q�1���YyR7 F��5�uK�6M|��|$�ɵ�.ç�8I���cJ��7|9����T�f�P� T�s�S��#���Q�3���ѫy7%����\9i��C��0*5Q���+&��a� ;�6�.�`���m�a�Z�˂�O0U� ��!U��)ט����W�0��$���gOip.9�B� �I�g�_7�z/�����lͣ��_�ZZ�&��Q����,��ɡ�5)v�ث�W1qE�W��V	����K�������f�����5�R��eǣ��W�Aη����V��;���m}�����n�!����?xv�a�K�s�a���k6w�����o��UXoyH��M��Ϟ%d����i�dbbM}^h�Q:՞���K$���g�w��_�m�����jRe�޻��ӫ{'��-[�~ o6�ֲTc��H�q1���Ǐ���v?]���2(�{���jT\8�j�&�[��	YƳ�Ka�룱%�3��ڄ9N����e=od"��u�8�;�ȲDS+���|uP0��l�T��c�%fnW�Lo/����J�V_�$2�r�U !Q3��K�@��TY��$�NO�M�i�C'^=����wm���W[�o�����i�r}H�]���}�f�mV�n"5��|¹/�x`Hl��t�}��A���2V��eP�<
$(��AM}�}� `�#���zY*��B�'Âk�/�wsLii��;�p�7w��{��=`�vz�^�~��aG�s�������+MqĔ���\�J�D�T9�k��(SU=�>`�䏑`)Y�#���쁆b���[%��>;lSf%�̟?��1��'�i��uO������>
��iF7jRhQi�=.���c7%V�b^5�A�>���m[�
O,���3�y�`��#碔����%�����1>��H�ș/+kuo8�w����5�?rp�<�ʼ�Sޏԅ��ZT?Ԅwp�
����NL	GQ|�IVal��7���$d�-.u��g�����|�{j�������VB޼r�Q{76#x{!f����8<��p�H�65}���~�/�����Ou�N dd�<�Z K�F�(kWq�����q%ֱ���~ +q���*=9�񫀮,@�Hy������8H�a�ہV�e�����	?y�T���<+M���TA�3G��P��_�k��[�rr$k�kR�x�"������<�@�xql}��D4�����1�B5BW.mq[�pŊ]�(���2�}	���Bf�G]�X�XlH�u��W�T�}�	��/��R��ۧk��i�}M~����J��5��ī����%�QOᰧr��(e��qN�%�	�9���Y����L�TK�<�W/��}uI����e�LfЃL!�ô�;��nN�j�f��sb���X�pY���5���)���J�h|~[�J^}%E�^�/�nΩ�;v9@ i٢��QZ�ÌC�"�1�=���'�X@��8௨}�<��~����6/GL̗"�Gx���X��g���-�Z�TF]��/���H�T��0����R�}��@��K�	�y\&ӟ���~[��~��tl���8N�F\ʙ�}h�9?�4����سRW��RT���&�I*�(NDBYۀ��Y��s�,���s!ʷ��sy�8(O��B*Ovm!]���,'������t�[a�4m*��U��ո��T�G���S�@ڨ�=$`��C���ٕ�gE"�9�y�`=9x��;یl��5P;�V���:s��v�s����)aFR-�m���;����eh�Y�p�*���j98Yx�eI{YY7l��
�����O�t?̺'���jQ�d78�S��'lb�Ӟ6��,E�zW�W%����eʧA�nYҙ�#��ӓ���B��d�Ѵ�*=�5"Ϡ�v��g3���$1و�잩��D��7W�p�틸�ʧ��Q
,O|�ef� <���ө�x��c{��3�U��8��9Q[^ӡ����������>G�����������$V��͈%Q�� uu���	����<�uV�3�����i&+�3"�� U�40u�/�0_�[�}��]������������jVp����ߍ�h��e�|hh�BE�� �V��*���E��{���0H�����@���e��.�n�@�)��\��A�o�g�!���3�SŮ�:�O"���_�b>@⸃w�,�(����싅���p��f�@���PѬ����y�8ۆ�Ra�D�q[}�IKt���NQ��q}UG��2�BG;�f�C��M�~��������͆2�u��� �#�\BC�F�\��"�2= kt�d#��ų�L��i� ��'�$�e���嫾�-���_��̾I���i*2ho�?y�.�u�4�KG3QcM��M�b�F-^�����伊U3�>	h�&n�DW�ݕpC�,\I�6.B��$=�n��\�S��N�܄��ף�>O��FVxfS��.��PCHa虃�)R��Η�f�J����kyy->�ꡒg�΋�U�g��V;�P'l���r��ض��쉥(q����E��C�|{yc�/�lOM�fc��4Q�� ��r��]�D��[�m�e��U�H�<[�-VzI�ZS?V��n[������y�b��u���
v��׋���������������軓:r� 	�k�D�J�ƛe�$��<�ޱ������=al��{����;��:@l
�Ƞ��d3/.���ē3K��A��|��ɤ%=�[�N�
����$9%�Z���(�iv�
eZm�+�ic�f��)��v��shA�b�9��O�d1ːQٍ�=������"�7��Hu,�� �Gsr��ik5��nU��i�����L�p��@��naΈ��hj�n�̊��j��&��?u����7��[E�F��%jh�=�ɍ8d�DY�=x/c�k�r�����P�:C��Ŭ���^J�8)`���k��e?O�,G�f�5�g��9y`��,��	�I%�C��s?��UJ����\a^ɛ�n���-�b����ܻ3ec[ڛ:���C�Z��\;:î\[�۳{0W9ү�ևU�M97].۷�'W;���~�W��wH_t�N��}�C�����iz֎��"��F���&��(��k&s�|ھ8��di�������/-@΄�������E��c��յ��)�k8��+��E��r+W�0��^}�G}hޮ6r���ޘW�F�N)o*�⣄�?�4�%���W�(ZS��L��G�s�׻�h�,�[es} ?��sk���sft�t
�����p���E&=�yO��w�^�k+�B'���u�44�g���p�����������Wܺ��ޛ�;[j��h���cOLN���)C?X��A����zQg��7%�^���
� �p_
���X�q���S�R�DH�O������������@�T�쎶���1��V�/��o'y�BHW.m��ր��,o���.�pE�H�D��T͡�W-�K���a�gFP���U�R*�WlOZ`��_jF^�����������Ƃma�)q|�\	�~� �����e��))"Zqn�F��w�1T�`��ᩓM�'�Bu�%����L�Ԏ4�cAhb}J��Qj�d]R�A��l7�� [�>�SA��IZ�]��Ƈ��ͥ�����=Az�����0IIɋ�쀭f���}�t~���2v��ҖO��k��1��v��_�*AK׻-�~ꞅ�����&K��Is}�-V}��c���^>����B�]���z��Ӻ ��ޔ�t@6��6��,AW�v�p�/��CǙ4�X� �}��Й��p���P�{�f�����S��*���6J��YB��z��z�D/~5ܝ��� �����+M�2l�Z�rg�]!��dD2��/gM�ڴ��O��F� 03����F��x�t�W��Q���G��y�w��×�__ߣ]ůj��o^�F3��4ok����}e1k�D���l�����V�;�����ӷ���h�}�ep��n���d`?�LWvuF�]�&t6�=,&w��U��`!U� v��u�s����lٿ��;�/X]��;��X����+rvܦ�(`�f9e.�;�t�'ٸ�k<,�& 3Z��}���ݗ�u�$>�
s�23s��/ۊ�$c�M�醎���d��			��_��7O�{S7�-�⏠����*�D�������� <{�ȩ�}p\V��%a
P!( ��"_ي��(W03�.[5]��q�&@.��QC�����/XNi����_7�X(6n����&V�C�=�8훷]������Sf�ZpR�
�ar̖��C�C�έ�=\��
���X�[�{D�)��ӱ�CP��՗�a�Kb�����e���w��6o^��7�,��hdPr��/�l�����	m��$�|��l�7�����_��=�~:�j0��X.��eH�߰,"[iZ��m:k\pq�3�V�DL/ �q��9Oy��L�N�6�}J@Bu�o�V��~j9ɘ#���+��j�6{\��G��F�1����K�J���ǩ\\iTk^r/9gl���ύg�9�]�!$���)~�{ד��d��,F`r-�y�J��K��B����:.�-D'�� Y�G��8,94R���Bw��b����G���j�2�����|٥P�=�z�a�z���`K��N����yx�9�)=Nb�x �K����A:t���0;�y!����t�7e_.�����6���B�b���R.\��=��(���MFX�
c�LMDT��F�ʢJ��>�o���HϿ���4J�GRY����k�@�s�5�����Y�?�U_W�m\N�6�鮓�ѳ)�ጢR�k�p���E-nD�)_�op�͌�t�z*;�$��EJ�'��H	�/�qs��`����U{}@�`�[ƃ'vп��`���>i����쪟�S~��E����=������pIňY�!�
7��ێcA�F�Oa;�|f�Og���>B��E`�@ڤGwD��V�����.b ��)�UL인��|��%J&�>`6h���Ud\R�`���Yc�[�Y.���0�ϔ�!W*�_r�t�`OZX��%
���S���Ӄ�?�it�
����6��!��>��ZS>�MG1�f�N�J�뉬}/L��(��Z�L;�dmb� L@"�6�����  ��\��܍;����Nz�0� ����|���G��%��>h��O�����]'Z���>g���a�����=�vX�$��V��?+���^�M$�]q���s��ڛA����o/����B�n��9���|ltm��O�+�x�jx`<�a1��H��r7薔\}�ˮp��ŝs�n�eK�Xz�����g�l��o�"��\��zR�=;����Ώ���9�ߜ(��%������'���0��ҙ�����W�
��
��fԖ�O�����v��)TSD�s ��W��*�J6�PK   Ŧ�X_��.
 �	 /   images/f557da7c-7f17-4077-a29c-07168c914697.png 4@˿�PNG

   IHDR  �  ^   sQ�   	pHYs  �  ��+  ��IDATx��	�d�uv�Z{�}�~��t��s�hH�R�DJ��HdX�"��$N�8��h'�b%NE��H��`D��(s�q.3=3=��{�~�������s��2e#i�E����n����?�w�ߗ7�7�7�7�7�7�7�����B/��ŋ�����o���)��d�����������2"�)��W�ċs�[��O�)S�s�Źν�Tǽ�V��{��b|�o����ܻg��w�+/������;��=��Zڽ��>�������]��}��1��W�d�c/�>��f��s�����IE�$v�B�I4�O^g��,O����{�����,s�<�u%��Hә䅓��Q�f�����ۻ�#gLw�����f;�4��Q�u��4ux��JPaG�H������;!������wj���	(.Kk��5ZA��;�������Z�pj�(:~�߉ާ�i��ӛ��Ⱥ�V~���c�8GI,�V(�,Qb�wfQ\HB�\7s�ɜ��
��@\��|/�@����"�}e<'t�s�(r��ƙ��L�i>�R���9��y�8�A�e���:�x�7Kr�����17a85��b,�[�|���V5���p�"���^�����p�t�YPk����+<�������IJ�H��	���ppX�8Ju������s�1%p� ��B�յ�2c��7/x�?g\,��_f��9΋���^��Y��}���t"<q�aڝ,���uC�S(����� �t�8~-t> ���3��$O�Z�����s=SZ
^%��H��n5�����/a�1�<w�8ﮮ�Wd1h��g��@�r�̜����p�s�	��7��A�N'g6M1�-|�Vo�3�Q�'(H��G��q�F�4C���C��NR'��4�w�%Ƭa\n��y�>��������a��
:��s���s������ ������`����u�@~�	�+O��s���LF�48�v�8<:
�Z����$i?�g���(��(��X�F�ǳ(��!x#ov:N���(�$������/�����?�����?,:�n��ð��9�!�P�(u$E�Y��yƏK^K�ÂF��K�.Ϋր�O���$�\�o����`4��������/����v����6'O'�Y����.ԟ���=Tւ�<���$@��!���{��̷'�� �"O1���_ĉyVk6�o���I ���>�܌���|<c�����`�o��O��M&�N��ΒXǆp��O_��y�7�����,J@&�S�W&Q{�U`qj�i8���gnel�Td���G�9y���A����>�����s�:i+hd�$-\Ld�]�_��?������5/T^��o>�΂���Z�z��~���?�������=r(����R����垜��K/��W���ʒVO��G3�]�b�s����F��q�u���ϳh�y\1,�����C��Y�a�Rh��(]�u��x�}�ђԈ8
�t��V<j��LDf���.&�Z�4+����A���G���(�3:����j��ˋI4�Q��n�i��q�,,�Į�`
���H��,���F�N�L&�����F�X��;�Ef���9�Z�M��D���/���\Ȁ����PNB1H!�N'x�M�V� ��@�� 2$���b<5 �+.^h_��5�y�L�%QQj4�� �1�cs
<�kzIa�뻼��.f����K�ە(��ݽ��tii��~`�X6,�>�K����Q��4�91֐k-� 5�Y~"���-�,#�9�r���:5���%w��l:�d�FB=��h<[X���fˋ�(#@�c�3���P-�f���~
�n�+�1�'�6�u��&H��B�Ҽ��U�q=]%������\R�
d��gT	E��vr�ρ �r�e�YNe��Y�%T�4 ��Y��Rh3*P�sf�@H XK}�S%B�F����� �!���>7��Ƹ�C��^�sN�LUFA�'J��.����JP��\�h�HNQ"�T���~� �a	!ˁ�Ʌ��e��B�����X���gY�����I��-��9�����[�t��j~���{�Ԧ���d6M��$j������������v+0@]�A�8݅���c���XXX̩&�{G>@{�D	�@�H����M�r�b.M{P��y�a�x޵z��S��I�5B�Ó!  3̒.'�8����J+.�9��"��h˨	�0���EqW�*aR�a�=��0��|�k��P��it;�D~u� �`8$�����o7�<������~��"]a�)�"p�,� ͆$�8�=��t����J��ci4F8���f�x5�ԜP\�Eg0�A�6��,��B] ����Z/�=���� j�� ��`D���R0�*�5�l�VL>�[_�w������[P}��B�����_}���/����i�o�GQ�I !�,Q�FhQjaC���\6��%��`��rb}%�aNv;MJ.��Q )h!�@�0GCwi�S�G#�.ᣌ�P\y�e��	a���r;�	�L�r��Ϋ����d4[�xaqY�h:����%�Э�~��kN�uQ�(��p֛���x��H��P5u��G��J���J���HjE%bS%0� Li�d���
���e���:i
�����'s;T9�TA�p��)���T8i��q:��)4.��$�(�����Ӽ]�>�A�@X�y�����3s��1%3�=D=�P�S���-��c>�q��Pz�z(���0&�v�72'����)Ȃz��^O��a� BО�Lr����<I�
���B`�G0��5A����P����(�Z������ۋ�k��xc6C�jfQa�2��Af��?�
���`�6��a�h$0f�V��9)S�[Bb�����3C� �+f-�RGA��d8�5$�Z-?&N�7���)��I�E�]U-p�O�KD3-��@��i ��-n�S�8����� ���F� �̼O�z����7ː���7�{5XU� �����:��vʅ��R��.wVA9cg� 4hj3U�������J.��x
���ST.�Ҁ��q_bdB5c@�x^�;`R��-����ΜZ{����I���t�^�ŋ�q1Gn��M�~A�n6�a8{)���aPX�J ��ѱ>�,I�ޘ��x�a=I/��U���GJ~U�E1��h�����L���0�d+έ�B�Vn��lR�f!�K�n��� 0!��2�wjE�r5q`d@�M��(�DF7=O=)|O�����Swiq) ����Jywq�9<9��=
�Ϣ�~�K��?�,g��~�J"	m!�bV6Ή��%�1�
FC��W���ũ�Y ?�h�H)m�� o�n�bʱ�YZL#�?�c���vS`:�~���àSo'��1�8�s0������g�ѝ������P��:�Ţ?��g�v���Ǔ�����A��ѩ���$���f�-�$���$��ޮ��x'O�ʓ�^hLGGd:�T2�T6W#]���n>��������O�w�?�O(� h����s�a��Ȍ$�K/~��T~�#�G{T�z����{�Z�(��Bw	߯A��dqy]�����ի���j/�z�T�f����N���1��@�P�O"	�M!�N��.M%Z�m7P3gjS��N�����i�9:��r
��c����<b~qe���N<갥�[��uX�X0c�1,4�R�������,=0X��0,"�t��iLW�3Qk,�z��p$ C�nueMT�r��0!�S�en`�8�|�ve�g�v�t������j����N�nh
�\?OאQ�KD�'A�~ =)t��CF��l2�������K����k�I��2�1r�uMp���'gΜ��h�5��{�a��󦳱ފW-�R����U���{����7��2�����
����a�W��x�R�O1W �@2�:�6���Ů�Z� ��T�4���=��1���hp���@ϫ�V�[T8x=L��#��%�_��X�5�zb�`����ʿ������%�|>3ʧ���9���Uo�������P���y=��.vkG���Y]ꀇ���PF�]���'��񁜃�988�ӧ����"Y[[��_>���e�'��k�����4G��d�ziB$�1:o�*��tbs�xM�K�X�+���)k���S�+�SO�l��1�2�s����=q�P��5:D$ŘS��wC�{�I#Ý6�NZ#ݧ>����K�=iB��#�
�I�)������L�YI��W��@(��+�A*�d�V?x*�Z�y���Q#�K�^̟����Ε��H�5�҃W V@��6f��O�0�����^k%�p��&�t��ww��kY�����'�^���q�s>�;�����L�erZBW���BGFN��=Yjvd���p$�I)���ăci�L޴�(�x����@��Z8J�T�|�`�������oޔw�㼜:uJ666UXo�8)����T�|�@�q�-f`����:sK2	��E0���"wH����0��D�`�m���̔��*XVR�`�H�X�Hs6��S\,M��p4������0�Al�z�<T���C�UAG���#ˡq?"�0�r��x�!}o��<RX-wۘ�t �J���`�!�=cë+#��EZ���b �[��Xvoߒ�Ŏ��T@޴x�S��P�y��&@��Mdt8�טV���Ǽ�BB�� �̘��Ŗ
�@���zC -0r���4AnB҅w���Rc�hh�pf!Uʘ����,.�`�d<ʩ�u�E�-o&��+�>��t8��L���
'^���Z��}`]�A�b�~<����O�C�t�R}�׷ytJ%�	,��)�1�z5�5����^Z��8+EV� � �u���^_?�p`�x�,Xw> u�ݖ)��ׅ�b��`ܗ��-���lt<�^��߫�5��{k�s0��~^��LaН�Ȓ~J\�J.tcn��EO�����R����;�'����$�!��2������}Q��_�{G�m�I�2�<�kक़�;پ�<�(��h�筬������Ғ���v:��zv��T��Y+ޯ�lm�BIֱ��7tqOi�z��S�S�tCoCa�'��9�2�Y��Fi�
Wi�w�Ь\�a�5ic�j^"A-��c�k@ᧉ^�kY�	דGѐ �J0v@M�"��`E0�ES�}��jK��aI�5<{�@��7��S_��F����gs�? !1�Ǉ2���,AcEˤ3��C	d_C�Wz��ɡݓ�G���wH��Z쐕�t��)<̩9�l:�;y�W~��3_��jQ|�M��y��N�{�V������cYA.uZ2�}M&��Ի�ȓo~P�;2��8qNKJ����ce���� � >�0�$��TaK�eO�!M'r�;�$���?���~�䪌���{�RLT���`����!�����{ 'W��3ix����`,u�k����J�C�D}�u�E9ؾ"^R&��M�8񀬮��7�h��W��̅�
��7v�dayh.��}9t�2�������� %q�ߧ������& �@�=H��[�����'~PNo�H���y&\`@�����˗��7d����A�4a^�����H����my����C�R��<y�,�*�)��0��aUX��p>TfQ���#�֠x�`j��D�}���o_����rt�&Q��En�37-�"S�%��[0Z��]97ADG�ǵy�;�)��[���kr	�s|���r��.G+�	�7K����VWW�گ>Eֱ��׮�3�Z-����{�^��3*y>6�<�͹If���稄�Z\��Ǻ�^��}��Hv�<�ߣ��,�յ� {�Q��*0L��pl�dq=�UE6C�����w���0�4�N�n�^,Oήm�>x�W�<*If��c/s)�k��7�|C��<�/*L@u��R&����%/sW������5�A-��+����<(��9�My_ (���FWNn.�3�}Q�Pj�t k�K2��8���d��!}) O
�Y�<�f�j�[�#y�Ժ>W��%�i^f ��?����_� Ҁi�k�l���͛�Rw5�`J�J��}�Y��mN�L��~��0D��.��6=6t׫r���Xg���`���Q�C�6��yF��a��:�Q_�5����m�/����wyqE��������O��t{tt����/^��7n(��Z�ܸ�|6��O|ʹs���]��׾�߭x�����o��$��<���0�$�fs2�gӕ+W$L�j/�gs�m��Jk[�vgA�!`��r��ډfI���|�������߿�/��+�����G��G^��}����A�.N������B�B��RX� ��:��,�:�P�,�i$�^~I�w��)��59���JT9��K�B �@O"E�5(���@b3������T��y��Med	�sͅMe�>�5'À� 06��L����'��\����*]��~O7�d��o�rQ��ڦ����o���\]�����=�z�ܸ~V�<���˧��3��uVN�?AS��K/�5�2��
�d�D?���B��an`�Aɮ����&�Jח[����&xϻa�v �D����!o��P���Uypk
��|��ɷ_|>�\q>��Tzrb�I_�L꙼��W%�f�@�5�i���M�$S��{�rcmE>���K/��!�K���xtP�i�lR����-z��ҏ���rɡ,Ξ8)�<�\�t��S(#�@_״��y�\=�����{�qQ�Roll��o}B^{�5�=S�������Z7<�{�7{:� ��9h�:֋J����q$X�˷^��Q�o�R��OS�P	��u�����{��N����Jo��)�H�����%��sU�T��}Y]Y��~O�t����Ĺc�� 0��W���M��I��2,��#=P/c	P����'�[�d�`40����D!Ja��|���={VN�<�s�;��J\N�5���\?*7&�Q��S��yR?�:����St��g�<� v8�2��^���0G#�7�q�٭�C)4��z���>�ߗ�7���rG�����.6d
:ܽ����ss�c��qj�X�$rԵ��z��'t�HG9�_[h鳾�·Tq%c�X��l$�L �MRy��<�r�
ρ!0�#UF��󉺣��
s��Z�z_�y���;sV>�����3gT��{x�����d:�z��#G�by7�'� qo>��|�_���%Jhf%J4������wn�h:�k�����W��ը/�m1*x��{]v�[���d��y�txSi`��ı�Gа�sA�����]��{�1��w!��s�q�Ϩ��,�@��H� ΅��2�OO�K/�h����8���V����x2~���/�G��_�'��K,��^��}����8uLN�K�d	mׂY숴�f��.���V�tzS���n�6aݖ���{�Tu�[�nG�e�0�D+��t���j ɪPL�h�nʘ,c�S���2~��P��5eC���נ ��1�m�+ׯ�&��@���� 7`���ч> ;�.����w�E<�!�x�|�S��o}�������?�C���!��7~K�PP	�%��\M)��"j��}0�!��P6 ���w��*�;-?����/��s[s���W���eL�e^�#�s,��b�a���-�◟U��wd���u�6k�p�����2<���	�?5e¸8ݦ !�t�n�* #�uy̵_L��WfS�b�Đu�ql�ž�VK0jS��]�1��x4W�\K��47��c=�i�Y��.J��� %T�m혞�� �ʧ�B`ԏdJ`�1�=���ЃbX���e� ޢ𠫑 ���8<Ig:ƹͺx�����X붜Xn����{Na���e)W^&=z�'���V�H��ٳ�C?,/����%�,ih Z�(��u}i�����u��߭-ɛNm��;�P�Zz2;��ڕ�I_��x6�B1wz形Ǭ���,�f�X���U��Y�#��͊;L�C3�P�!4rIR(�)l�u^Y]���F�2�c��@�罨@	ɿ��4��=�}�+�� )�˫r{gVYWN@Q,��h�B��`Eb�Ν9)K0+9�4�Y'��z�����N5�kI����E �Ul�>��	h��=Н�ӲV/�y�r���<X�nε���+~�g�¯��r-O��	�XW%0� P�����1��2����Z�1���L�)��'-aq}�EY m.u[��mK�*a����`ޘi��A�N�R2�'ׂ�e�p���N��3��W.OT�R��O���\"W�8�k4�ߛ�6�腦|��? _��3���*7omK�f<b�L�+��f'7O�s :���-����FCbK�����M��@�?`}Z�`�7�+���Z�#k�r��v�歽�V���������7n��vQ<w�q&ߋ���zB���@���%�P;��^�U>U�4%3�D�F�	a��z��K4b�(��-s��ɼ M��Z��D�o���0� �����K�� b˪6�UW`���q@u5A�@��+z�$s��I<f���r��)Y\Y���U���BPܝ�'+�<��{ǰ�nɻ��~��X�CX���`e&���8�,�i��&�Bb���:�y�������ໞ��FY�͊N(��IսX�����2���Y�|?����e�����}7��:P��H-g�-c��ο�,|����]((z^��+t�јA��L�V��qP�3,R0^�ysQŪ1PQ-ab�B�i��]�� �k�Z��+- ��/cΒX���}ta����x4]P�ZUo��V\�Z����)��Ռ^�?�����0��<\�-�9׋��s��zL�`O�Ź �o�N�̳ES�㾚/�0i�t��>U��0	�w�~-Ƣ�,�	c&�;�B���)�����<)Z��,�lm`c9�� ��W���͠�l���hG��Y�N�\�@55��a���N�.Nz�����L'��5K-TBŔ՛�r�bYl������3�qb�֤�YW����q��;�vv\�b� ��0��-G�7�^K�Xʘ����5t׺q����<s�D�S�w皚�V4e��I�a�����.,��,I��2ɵ	���ԩ�0�ϊWs^\��V���:T^Zm�߹�L.�K�4�c�:Yހ�jֿ.�UO�L�Zs^͈OUv������\R�Ur+( Q�@c��	@�����[FPA��[A;qn�<���[�7u��
dڭ�@3 	}\V��T�̱�2���h�������YfQ�����h�d���6�[�2lW#`�l�L����rx���*e9�n���(�>uⴼ�ꫠ�@���c ��͎!�,]���|\{�;���?-���ZkW����^���͵�7}�{���B�#���h��@��6� 91�\�$���%�A�:�֋*ҝ�9>:  hYK!U����!�"�v�Ք��ɾ�jkj񫐬b�d&FܘY�&��BhE�VK1���,���y�hŬ#U��D=�&�qrE�\�$;�=".\�8��kWe��o(���-���~�k��r�$�U|��G��}�sR�׈�M���s�tjw��<je�'�_����_>���d��rr+a���*ɠLHd�Z����Y�+�`��8+��.���g��Grvm���c�;~B����P5Y�Og�KJ�?J#�_�Y�Zn�Y�P��)a�ի�*��`���åۗ1c�5�C%�Ϯ�8�,��J��J���T��I�f��Ek�5�>Ž"Ƃ�n�)c}���@�"�ƯAy�N�f9� ��d��1���4J��|���D�q��ʵ!-rLR�4�-���b�vӔ$�-�!�bv�QA�|'�g��hޗ���e�+�*\��:&s���H�)�u�T�4d�e$��5)�qO�: �m��P׹�{��h�LT�	@3{�d�XX��5:�ߑ�co��N]��rkp�6P4�ܺ�z�R���3O]�L���f r�y2�:%�$\'���*�\��,�n}i�
%���%s/X���[�,Q���Ǚ �qLpm]�NK�Y�y�TM�*�s���k�қ����&}��F����`Iʾ/�ɯ���s�1ыV��t(�r�Yתi����ڴ,{GA_~�˛Ɣv�R/�T��q��~%]7|��z�XJ%�ǹ�Y�*�#?��e��#�Hf���<�� �94�d�4��T?�Ƿ�P~?;r��)9><³�C��,�Q�H�sp�4}�\�j�2Le4EO�%��8Y�j�h8��(\���[�����������=� �h9�#�CQ���錭���W�o�z�����^-���K��}��i{�qx@DD�t�Zd�\L�~g^��2��8	�uw[&����2>)�fQ�L\���s������Y��-~DB��y�D����؜���@��"u��R�|ӲE$�+KҰXo�ʑ*�e?�F@{CYXZ�AA]_�G�k/�	X�ׯ^�Ã�n(�?�O���9��]� �9K,&B}���*�,/�sApt�o�.����,7�Xn�_�?���wڗ,�D�@�6��Ia�T��F�d4k��.Z>�rŃ�x����˯�͗^�܃l8��2M��TMyi�T�Wh��V��0�UH-��)ˤ���s�U�eI�ֈ*�v� �Bfٯjm��A�74��D���F.3p���1�+]�E�B�(c�AS� ��X7>]���f��*�L��r5����z<r)�0�y�z��}o�[���!����Qn	МJ|�D�[Ě��Y�==��	�����:WeDړ�,#�:�T�w��IZa+2Xw�Z]�Ē>�d�9a̗VׄcȬdҮ���C��S��$��t��*���L��f]iy^fM5C$8��Ɔ���.e�t����j�j��uev�/]ΎV.`�`�֠����ο39ڿ�H�pW6a�y��g�
]�I�@���ge:8P��e�;�b��{�`eZB������ ޹KP�]�z岎�,=y�;ޢt�<U�@�9�Ω��Wc!Wo�S�e6��UVXWV-�c�g5�	|u��@��#̇4Ip��Q�V�� �r�]���HK��C/���Cnֱz$S �^-z�
����s-��$mz	��6�������њ%X�����yE�������7Z:�dWz��*�t��5��m5*�F]L����Ȩ�-v[��Z߅�fC�u�g�e����v󆜼����@@u�: Pm�����o}�X7�B�?��&�h�N�e5�H�����@���hx$�7��>qbS-�B�ΝmL�+b�I(*��Z��)��J=�m5��A��	�Y���جjQ@�Q�G��ebI2�@s�M\����J��+39&�i�V�B����+2��Ϟ;-���$�[�^�=[� �v��,}�z�5��ݑ�4�k�n�no"w��eeu]U���Z��œ��*�{B��K���\8с����V^2-}/P�2�����u�T���?��(y���"_��g�"@3I�xG�j�$�Y�B�����4�����#7&�a��.h߬�0V�C���>c��3��hR�P!P�xU�4���E�k�_��F�&N�,�M����@��Ks�2�Z�{��RD&��e��2����2�f.�t�^%x��K�E��@��nk���Y�w1>%�2�\r�\���^�י!���kuπ�v��4tS�,{��iv�cƲ_�}i8 ׮�Bu�3������*?Ԑ����|$%(�Qe![������ք���e�{ٷM�u�Y��fa���W����h��-=4l��͔�"?�J0f��M!Y�I�H�=wө*���/GG2<ܖ�3dp���U�Dg����]�Dk΁��T�r�\Km�ƙ[@ ��Y�ΠU;��n��e
|b�,}k(c��p�e�;h�s�9�)k���-Ti���&-y֫[R���
1>�H�Sw�)b�HJ��WIe��$:%�u��esZ�K)�<�
m��קȪ�p���ZU��h�n���LxR�	k�d�`ieXk�x2T�ǩӛ�g2/�������TXa ��]����f��=#�YZhk��?8���&S�`��阈�_���L������K�.>�V�֖%��5�k�Ӗ�þ���E@�� ����N������	!2aK4Sw8M�didY�X�i
k:ʫ�n�`�N,V����FwYˤ��%^YFS��Қ��pbXpU�����\�����.�*��ȭ&ݳ���	�^̘7��'�v���"��3
~�4`Q,�7�� ���m��:�u�8oo`�<��
4�4塇�G�|J���/>+�v�e��
;5�̹�ڭhM3�+dւ�28XVL��~@?oB��ϏG)t��+/-X��B$S�s���i��R�����!.��Y?�y�&��A��)�DѶYfj��L��$���V�]#i*���d����ךVeQ�NIݡ�"U�*]�Z����{�q_�o�
]-9��j`o� �,�rܓYZV�Q���_�1&G��
	�"W���%~��v�%Y�?��D��V^�^
�@��i0�۱��Gp1���@6��z����5,�3��� �Y�r5�`2���?R�$H����@L4"8u��w��lna��������~���А
A�,�J���D�*�?W�°FV����� �1�CN�K�R-J�*�	��Z����G~l�����,�����S����*:�[yUY��G@@����X��%`eBe^o+0|�W@��!�'Ù�R���7{
�ìJ^AD��c�U��S�ҕj�����^)�f�# ����k*��?-IO�[�'M[6�jw�6ֹ(ͽ����3#:���m���|T�KV�V�?z=�d�:�]m�l�[z���!W�k^1��)��"+�%tnJ&�fl�$�V�|*����`����P��0��"j� ]��0�GJ�μ�����;<�ކ�<M��׆���G\$����i(le}���)c�[�y�������[|ZR������C��p�w
�=���<q�%NO_ӯ��x�29e�gWcI��ړ��Y_[�,݀S3�&`�@��<�<�:f�2�Z������@�?򔛰�5ɧ��6��,�`�@��hL��l_��.-�H�����#�0�}��i�z��}<�����GU� 7���{�~Z�V7�?�ޕ�A,��EYJh�5dY�����r��,V|w�#��.ʇ�~R�6T���Veǭ�Sˑ)(�dÑ�\i��L'MbZ��:�Ii��5j�~��Á֚��br5	K3�33�D��nٲ"���e�[*s�+��=�����hZۈ⾡�Աi�E��2F�j8!.-O-wù��,��V��5w)��(-枱���ǠQS�����W+m��b�N������v��Q)��d�ٴ޼�"��T��o-=M�:L�k��hH�Ay�ҝ�D)ݶ$Wk�9|O�h�h�)"�G(�U�K
Q���%r�̪�A�Y�2�����i����xdeRa��|�jN�Q�ʃ�sU%�U��j_8����S%��}�z棺�5��ҍ�0�����B ���~*�t��K3�� ����e?+��Xⴶ��9M,[�֌ƚ#Ua�]U�����P����{�38wK�hz�U;z����)���M+�Rv�2w�,�f�!�sʆ6l��淴�)R�O��7H_�PO�S�I��K���)��RnYn�U*UY�=!#]Cŏ��>�1���x8���k׮���J�j)ݒ/�ǖl�j7>J3�v�Q�Fi$���0ƚ�F��[�	�vw%��v�*���;��,���a�'����hl囸�x8�vؖ��]i.�aL��,r���}��=� Vɨח�t('�O`h!XĚ�����zE�w��P�`��\ٓ,�p�tቼ���dԟ(:���M�wY�D���b ��V�(�ǲ��g�������%\��B{M��t����s����ey��m�0���+7�N*���:wN-���ұzـ��Z�l�ٓ A���)�j�g��;��!��}�����o�&[g�,qM��di��kșs$��e�7S���t5s��Y^,��`a��cu������׼�d�2u�D�b��e�6&z�5�X/*g
a^�uƷo�ֲZt,�����l�W���(\貥Q�Y�jW���]S�a�͔�L�~T���TImL�	j����MbY^Y���2�uӵ��$R
(
�.A`�7e	=�$��U��qQZL.���n\�6�f7lɚl6��İ�q��������@׬�,�����`!k+kX�H^{�5]�6�جP�њ&�m�F(L�bF�li�BܲU-�J7��a)�����֜��TW�X9%��cK�b�{�Xw:f�|5;MX(+��HbX�ݠm�	im�\2���W*�z4h7���=k翂�R��rEӭ�������&�>#�O��6�3����w�7��M��N���O��ER&�3sn��������5���L�̭	�l���?�4������]ߓ��&��5Yi/I�cx�V��@B=IjuZ��>;��g�ؐ�����Lϣ!�r�BKL�{���2|��d2���#C@ts���O�ܰ�\��f_*Mδ,�Zؚ??s[\�*3�9J�uS�̓�ʖ�x<+��Z�����F����ll�P�`G�b���C|�c<:<���*̫��l^H��:���Z�1��z�TZ/*NQz٬E4��|e]8icmm׮�\�<2��'H/|>?����x�(��ma�.;Z_�i`�Ho�:Ő'-r4J��ƳyrK�_)�R�Ga�]|�%	���^xI�V
c;#5�G:�hl��p�Y��M�g:�;���r��L���`ʃ-%�ngE����e�Ξ<z�Qy�⫲s��QZ��{$����R�#��SR#�����+ɚq��ha�+2�t2��+��߹)_��o�SO<"O>���ܑF��J�yj�.h�5X�_���e�M������(�}���y�]���ؑ��ѝ�xAç�]�I��Aw�/=����m�:���Row��˗�k-��"mvee��NX�A�ϓ�*'U�ncd�ۅ�pK�f�ş�zXk�)2X�Z/�R3q�X����js'�c�����}�=�t�bln>/ӡ¦v<��U�♛}hQQ�S-��Yݲ�]���5�-I�ޑZg�h�T�M�sPy4����l�j }�����6���k�T��i�s쎶��?>��	���ߤ�ft.�`��eB�ݒF�����ђ)h4y.��V��%���Za��pf����X%���ּG�{.d�LO�Kǲ�&�\=2\S*��2�Q�E+k�^�¼���m�Rz$�� �����{[�rݭ.��w����n�Vv�{������:�y�e�V��V�����D�5�\�fK[�~�#���wQ�m���,��Ge����@:������7�1~7�I��T���r�2�3P�4P:f�1��ύ�XSM�V��+@cI+����r�Z�j��^/����uSM���֠Eݿ��gu5�p�=��,E���v�l���t��W+�U��yК������ʡ�,d.Q���Z���<(A��kW%*M��{Z 73 �v?���E�%d�}(c��Vm��]��V�i�9��p%#*O Hs��h�գW�,��g-��c�p�לzj��
;
6.���&���E{T�ټ1ɿ�q�)�ܛ� @w�]�
��Ot]�?6���\�rM�����EpcxS�QOV���A��w���r�ʊD����Ť�^2��#_�r��,����O���d�^�(����H�4tQM���0z��IM���K�Pw$?��
����Kca�ڒ�C�NW?s�eL�2�XYY�ҝ���p�{M4�oymUn�9����AQ�~p�9�\�I�n/��M $@ۿ�[���dEYb���n��2���|LQ���9�3o��ܛ1Z�j	�W��q�v�ݗ��G{r�ԦZ�����bW��Y}��T���z����%%�Zs��EY^\V�FR�׭���)��H	T��ie���g�k=���ns��b!�b�]�NY�����Zh�Eg����H�[i���Mq��u�r�܀�㹽� �Д��e<7�̾�f�X<��T3������Vs�^�P�����U�T�`�yRMZ������
���$Vn��L5����;���t�6�TʗzGX���f�n�2�9_Y�^X���Lhr��7�b�N�3��L����]}�$�N(m�#�a�ܼD��;��#L>ci'���W�a�$�$Ɯ�6X�6��R�ֵ��(��w���P�s���1���?�MA;�r��k�f5N�U0���Mg��sL<��ʙ�N �m%J��:,�zݬ�ڈ��L=KLT��g
���,��uUc{��>���]�O[��p2/)����ng��b�m�0P�2c~K���F>��1''3חV1�ɵ�\u;��PT��L&@�d
|�a��Z����*PF�Yպ�?(O�^1-�4+C=�|��^
��u����<�����n��'��
�/��ȘÈ
V0f��e,�Qo�4���^ם��8��h���[�b'O��3Ot���<�FG;��~�8A�|Oʜ�}�Ё_�z���d9��4��<C�#]�ލ�HVA(;�r��	U�7��"gN��ߴ���dxl�p�Q���tπ!�:!�|�醮��}P��}�s���lo�tq�L&Ѯu���괴􂻛|�+_�O~�������ԃ�ً&���n�H�!JM3�������eʚl2�@��,� )�,�%i-�^ݒBQ�/K��,�� .3X)H�*���a�B�Ai�@�=�� ^"�Э���q*�%�u6����ۙ��>TlR��H='l� �Mi��+�XwK�;����vL�w�~�cK�q|Ua��Zkh}�Y�g��sg���ӰX͊c[O� �H���6��22��) �\s��猦c0�H#�5<�?+y(��b���,��sS`1����(?�����}��'?-�ݹEZ��iӽ�Rl9��h��lƢ�P�2g�k
\U��e�<�I����p�oפk;MLI��Wf�[F���Uz�1*�,����WetU����W=�uS��u^\��R&S���뢖ub^���3����WVK���������1�(�sVY��s2�s�+`}�yh_���_Hl�J����_����������W~�W�h9&�x��LS=hy7�i�!wU���������;*7�	d0�A�G������iI_��N]�P�.���bG����]}��E����X��Ҳ6
���s���� rv�0@�������Iys�:p�k�G��n꾵3�B'�ғE��h�c�z�c�\+_���<oB�~��p�9.۽����z�w[�/���-������A���^/�%ȚGJ������~��G��~�|��ض��zҒ櫍r�����?���c%x�-��{lEnt���&&�4Q�g:�;���s��\t�$�c�w\�o~��)��z%��Z��,�n��;��ܔh<��o}\.<x^n^�,�/��}����0K�$)��Bz�w������{
�a(�7�Aʎ���2�?�'O���m�0���^���'�����O������������s��$$�B��*���I$��� |�d<�x��2A��^^�>�0pVrC��qny�;���<U̴*-�(SK���[��A�'�l��eN��ey�Z����:/�cY�U�quO*CZ�k����ٗ̾�yBN�-c˚�\�b��%�t)�sn��+�\V�a%=�<޵ybk�lUsYXY֬ov$3���
*ԓ��A��A�2yP����-�e�dxZRt�_�yC�P�T"Þ�:���T��w�
�[@�����z����L!<xAK�h�j�y
l���pgހ�V;��h�3t0���P�:�+s�j-ԙ/�%D��������n� ��y�ñ΃��	�J˸�p��&��s�Me��+����sH���Myi�!���YIi�7� ۱��A���}����"Ҍwz0B(��7���i��c1P)w<����,ف�@',w�cb]���C	so��M���t�[/��BP_���ٟ���W�^���[����rp��K;�z��$ ���E.�y6��Nx�8����׮^�fD�q�9!EYwHK�JAK��7K ������T�cX��fG.�ti�,[^;�������ۅթ�
f���iХ��������W�Rg�AZ��S9Em�0ِ�'c�]�\6,:�ۗ#(4W[�Fꦣl^��Ӟ�Q4�UR#��>=] ��'"=T?�Y�
銍t�{�&D����M�E��ח��O�^MA�h�C0!T�A�K�~s���J^��K{�8��C���L~��g������]b���]���rcZ��m��~?q��I��w
��ǣ"-�����C^�I#�RkCڰj����Ң�`���r%Hcb4��֩9>�me#���j�1�L�a��ʋߑ�<�fiw�rp�i�0� rh�{��a��#�F0��U2��՛7�ч�+�<"��ߕ_��o��Eƺ}�
�u����S͒�49O�<��h֬��%�J����.�#�=._|Y�,�u�W�n��T�E�X����IK���S�N��Զ4���|��%9��&	��J�oYl[�rc.�ײ�]Gw��J��������%9E�Ԛq!]�ui#P��_�5o9iI_���.�����ɆT����v) ��<XZR�S10����Y��/K'�|�r��-9�L+��4 �VWt(�g�^E�w�n鞞a���!M���v�fw���o�X��#�ϳwx ���g����5+|yyE�5�.@�Tض��Z��>�|���0mS$�z%�TǍDZ8o0�^�d݅����"�^�s  I �mؒ�;���QX,�k�RS�Z�2C��Z�fIy��% 98>�Y���G�O`J�H ��{����~�
�)���h�"�ttl;���5k����3�/�Z���t��>L����5�&I�z]�Lx$�i@�W.��м����/�+�-P��9G��ǚ�׀2�u���=���[Oo� ��ᑼ��d����Ž�e�����-���y�[�K�&n��PQ���Y.{ֲW]�[@�� ]Riq}O�>����dZ͑�ʜ%qE�e0U����pO,�����s��]�j�sⲛ�H�����]�� ]�qV�8j��@��oܸ���{�����P���ޫ1h�&h>+�j��q�^��SC�וi���7�``=pO�MϥV�Py{�^�ߙNw�u ���Ӓ�����V�Ah-��)U�k��p��́Xz{{G�d&���z����`�{U�RyD<1>[X\�u#��e8�J
����̹a��4s������;��Y���&~+56DHE��� nҗ���)���="��J��D:0л��ץ�_ ��Yjk�KB��LD�i�S*�\;�=x���oߒd2����P��2)�� ��صr;K�5GӉD`�-�vo^�'��/���޺.)���['6��934�g���ca&�P��R( u�Afé|���/�?�9��/=#��˿,�n�&K�'���78�qק�� f٬B�W�xH���C~�ԕ!�s_|V�Mrv�)x2�X�!��d7s4��2���u��*�2S�CE�A��My�ŋ2����S���e��1�Ė�� a}4Ks�2��kV:�/?-�K���zpÉ�ݤ�C�՟T3���*;5A(����j��P0�����m)��tY�9�V�n%)[a]��_�i���}\�����*�K�^�g�yF�
�D�  �M��nm�Qe�y�Z�#����ߴέ1Y��d�w��������b����{��&�� ��f�rUr�I�M&�EA[l:��g�[�%:T�,I�6��B�C��{}{��� ��cD"p]��XϬ�K��@5	��,����h	X���u�,ҿ*�e�祥JE@����y�l9�TF�������r�x�5����@�7���1�25E�P��N ������6��>yt��,�v�3�NE8�?���j�x�e:�T{7�����#�؟7��i٣�5����8�]`���p�8֐*ɬ��X�I�E�ߍ��rgo_A���S��@�j[]=��hd
�t��'�k�ӴNIﺦf���/j�Zh��C��|�Y���Z�gz�>��K�@=h� h�L(3f�[���Ώ�S�)��u�=Nn���F�}�Ħ�wyЬ�e�Hǆ5�W� �@����L���X;!6�N������;�44�^X�L�X㳅u V��Qo ܒ���,��R*h��),i�)��cn
֬���'��kus��������|��o��S��ec�w&��d��APw�@�@�1�����5k�������]�q�Z��mY^j�}X����v�҅LD�f�6� �cW�)~g�8Nf~C`QЕE+�^5�(���?����7Hl�ehs�0���5��<���}X�~��D��Ɗ�Z41�n&1_���RYY�����ީ˻��<݄R����g>�ek�6-`OK�X��������)��k�V�ƺ�������7�uQn��ds�������\�n��*��qRa}�lD�aq�֥k���� 06e��Tn�_�x*#��г�U_r6�����-������Z,S��͎[ז�����־�����|wOkŷ��UJ@t��W�1n
 �-�,T�h
�nmZ�Z��u$H�B^ZY�hz;(������'��O��ё�������\P�������(@��TQ�뵘	�Z����~��SW��t��9�B��ţ1��������h���y�$��x-f������uo"�F��Q��=���	^�2�hU	�Y���Z+Y�6�$hBg���e�XT՚��<�cb+ز*�}i����>�Z>x����`[�#���j���J
�����bKN[�%��:��%��cW�ݹҒ�,Ϊ1q���c�t�����+ �܊sme���t��sg�%�M�Ro�V{<��ey��5NG��i�b����sA����&lW����v[,�r"ܻ�tD���qc��8�;�]}զJ��E5��Wfֳl�e{Z̆&Rm<��\���f&{;hwZ&�L�bM� _�1�(����״�[Go��3�k��vaa	���v4�) Ҍ��r�r#�2���9}��U�B?�H����A�Nٓ��̩ ����4�8�i���j���>=
P�{���?t3&���l�1,r���gu~��Zu������74tH�$�dX���\�S�=�u���t&?���^\��m������q�)to_j�;��i�ueT�m=�ɧc9<�!��Wey�F}���3�j�-/w�o>YT�O���Eg��1r�Ȟ:�%_��/�ç6�Y�K�em�S���-�Ig��ȴֆ�z�i���Wd����\�|E���ք�7�@tɔ���K����_Ӥ^���յ�-R��/�������Ɯ;y������2�%l-�v�*(;K*䋲	KQ6��c�i��<ֈ߸~Y[Rۻ���O���ݿ�_�,j����Xo*։k+β���e��ي����H��͗����tRN>(��{����lk�Q��n�Il<���M)�:t�[+V��K�@H���`4�ض<�ج�o�@{�S@Gq��!|��@]WFS*(wސ���4fIK�.睽]�\�P�¤
�/�K^���_~��PY�e����
�������>
w��Q�--PZ.���y�Z���ĎzCuՏ�}M�Z]^Ҥ=����x�Ca>��Ӳ�-�z���|&�Ъgrύ7Ԃ�~г�=�m�R&�Вfܒn�%С�C0f�y�=������{
h��UX�d�{Qf�[��<����O�MQ��&O���~?I-w���*t�Jё�5n��~����}w)\��R�����Jw��Pȏe�PZr��t���mN��0�N��C����x����:jS(LƧ�:s�*��3�5�����Q�Zt�l��jw�N{����h7�}��e��*;�""�դK�� �sP+�C1�I��iR�� (���,KԸrh��Z݀���͢o�[�ˀ�eb���������Tx��S�Q�{̰��΢�F��\�(�ֽ�NT�p\�u�:sc*�(@�p��A��Og�{*=�9=�4��dr2�
���`8P�{��ZU_�֫.�������yLfLR�T��&�x�:�{#�����{<��f)4"N��|����zq_��'��q�)�2�p
�l`csMF��J0uX�$P��?T���T�.5m4���\�9.۶�B�u Q�V��V���YI�c�:��x��1m�tg���s���v��":���t��-e��Z�NU�b��l���7^u�BK�;1ﳟ��&�,��}���jl�j�!@)29��S������t��%����학�k�!�M����r}W~���������Ӌ���s+=�Px���Xv,�?�F2���`�׶w�ӟ{F.�<�0�-i&jo/�����=��SM(��8�Y�a.Rv<3W��s^&�ini��b(}[��M٫���9�g}���j�l��[���.X�k�<W8A���r��Ui�,;��ge^��Vf��x>��Ϩfv����_�lp*����S�p�:uN�oc�TY�\Ӥ*�S��ɧ?�)-�j-,kw�P�k��;�!�g�}mXA�����QI�/�
~��w�����X�6�䘥[f��剷ʃ.�����gl?++&��y.3��1Oa��hVR�m�%�����+?��z�(���F��.�naZT�Nն�?��e���;ıXs�{�G�=ex�6�����T��p�Q�	y;�=�v��{�m���3�{�o��W�����'�$ӲDN���K%x����:#O���a���f��^��3���{�fWY��?���5����@ �HW@�)`=(b=z*�sQ�
��D��	��T�I���}��ٳ�^���w��w}��/.�W���{�w��S��װ�[��{Қ� 3C8���J]C-+Au� {¾D�%t�������c�`�:���u����VK�qf��LO���k �黗��*5�:�L��G?3VUc�>CxSt�*���gE�%�I^6ny]�s޹"����A�bz|B�ܠʙBU�\�Ϣr�uA�{��^_���^�U;����j^%�4��B�l��"aI���X� �?�g�/�.���ܕs�|��,'?,�S�d'�\�V�p|�l�ca�\���ww핃����T�7�Cw4P�E�y��`.\8_�r�I�wkf�"1>y���9IW �R�S��2���yjuш �z�ٷ�W鱹��0�9ZS2��>3o��X�-���5Z�c���em�-��FCZF���k�<��-�M��h/��-dz������<��Z�C�,{V���M�	ʊ��佀T�#Iy)y��F�[d!NX<5�2>6�����Vt�;w��~u�|�}�#�X( �ʔ�P&�tcej�1���z�����M�e����揳g&(�f�Ѫzb0��쒙��S��!f�f���e/	jh̥\!�08��}b9z�p������8tF00pd�+ �j`xD��fAP��РY�$���L������{�Ѕ��3�8Cּ�V�����tǌzh�Ϛƫ�΀� ߫ϔ�4~�E����{YVh����.u�5f�@���z�լ�mŌ�3��_/��!��l�I8��K�C=�N	�� ��/�H�����W�������n��c�Y��P��W�\�����| pA��G��������qN?�� _;찊J�������
����p��0���%ϙ9.�3���� x�Yz�AԸ��Kw/T��0�L.x3����u�M�Q&�ݣ�1��bH�|���,W<D��A��g�� �%[A��{�s����Ȱt�@��bMC���S���&�>�|Y�d��A&���+ \Q��rF�־ >��(Pu`�X<!g�}��^���HJd]�u��x��m�vY�n�t���"���t�"�f7���/�--�k��9��G�`�1HGF妛o�}{�K�@���N��#����+�$6g ������H�����J�5F�5�Qb�{g���f1e��nVΪ�>s3h��<7X���x��`&�K���W���?�p�K��L#�m��c�|��5\����C`1��c��EĲ���������Ћ���6�3�[	�*%3�A}�@��2T��j�'$��,�p����43P�,���0�11�V�LjҔ+ߟ����X��Y��Z����푚�N�[ �̙m�Q �bƎ)�!�6b
[����J�ne�_F*�N'�܄����'���"1p h��kz�r	543��$����%�7�,oY�BN�I�dA��e��J,I�}J�hrJ^ݸY���5 ހ/� ��c"�$�e�f��䄭 ��'(���rPU͌��OC�[p�ְ���M�UQk ��7�MIss+�+ԣ��Q�a?/��^Ѭw�!�HOo7�i�H8j�{R�NN�,}iD���K�N�������$�Y�j 8y� x��m+~ϧ����	��۸I�.�&�9pz�4�>ރ���sUu�fd*dX�L~s������;��wY�rv�F��u���uc �e���o�N}���?��@el	�᳙��M��st|0ⵂ>����({5�c��������錤�#�A�L*�Ȃ�m��Dd~�/ ��w�\y�}D�N� 9��V���dT^#
�-3����z��
���*_��~`M��|L<w�ӣ�PV�~v����m����53e�.|Ş��Y	k:�:���r۝w�Y#q@0�V����6��'u���J��`�+B[��˯����;.�l���?8��>�H=�a���ѤlذE��;�����el�d �Q�w��t9�]�u�_e���'���n�a��!pv��x�I�a�qY�0>�i��D3���N���f��НG���ƼeC���C���\|��"0Գe�A�����W�14��Y��T�%I]�X�
?�)�0"�!��P��}�l�I^����С$[�Ԍq�[52l���8D���i�ޡ��ե���B��Q�h�B�j|ri��Q�]�u�(EST�\d�9>>*��ɪ�E9WIuU��~-��c��2K3�Be�J=>�w�@�����Á"U"c�Hv��L�,�E�e�idw��F�^R���P�u+{L�7q�]�Eʐ�P64 9� �[%��>�W���>h�HQ�X�+Ã=���O��tтi��Iscy�GF������z�HR�S�X�Cp�qJ�BF���F��&�T��0��z`�E[�8�E0 ��?�p�ާ� �y �N%{'SU@3��8�l�F��{X>��N��D�Vg3�:�X4N'��\��9��x�k!�����^$MM�>�R���}N�Pf�φ�KN�i�L9Y�rS>7  ��1o
��L�D�(�����%f�Q֣��d,u̌9��Ѫj����3Ih���QIOg�� �W;�O ?�m�ݱIcL�f)͢��T��x��?�}�Q~sӗf����x��
~��d����g�=�|�Q��'ؼ<�����R�8�k��%�q��8�n�˥YuA�xUO|Y�f�Ƕ�Ď!��t� Y⿩��6�;H�#F9���Ǡ�Q�F��s��e�l��c����T���<�����C�F�|��-
��r��@4j�r�6�ЕC�CΪI(L���wJy�f���0���ҙpJ!��7Y�ҭ�[ Q͆׼��� �b��gp*��"��\�s�w�S�'�`�Bڲg�_+]{�b1>�,�EJF�hw���@[2�Nx� P1>��c �w,s�eMI�<{�k�T*0�B�B)\� X��S�#b�D���X)y���l�EZ��Tq�����b¥P6�To+�-�xJ��;��|��z)h'z�13��Q�S;�a�xC<�H��h�8��s��͚m6A�<�ʈP%м��� 1me�L/�O��eE+R���wZp�y;�a�DXnˁP��[F�Fe�qo��s܂
��G�ec�%���5�_D�8�%�Y""Md�9�b����8����ׂ�#&j�S�#��	J�ۃᡰGWl�� ��$��!� c�gX,\ �z��t-�$@f_��cB3��:�foz�C�j�b���N�Y�M%�L�	" �Q�r��A�m[��e3��:�
�`��a_�k�m����X�hgf�]�<J���y<��O?��č��ȭ�����v�,��y�GF0� � dJ�3�(N�}pC�Z.HOw�lڸE�>z��_(�*�M�T�����쿖@�1 �,�)�Q�	�d�g��:K����{+O����S$h�Ufz���3��,��MNJ]u8K��y�ZC�C�{��)�Ƥk5*�p�XC\'� E�I=|���f�'���Jp����»^���0*�nא�4�`�=�1��T,(�C�hU�Bc��E�a?F���|��άZ��yF��%�1ѝᢧ�Q��W�b�:�������}m��0�,C�Sjq��(R�d��
�)��!^���W)���1[�3����`���9��,��xMP���牟���������5e�A�v�..M�ul	 Xt,oy(��C/)�q�s)x}����
���H-��� ��@ ��pq&Ѣ�N��~>���u��/��hXyN���
�c�����Y`*� �_9lFyQAd����^k��= =4' �T���Ӣ�?�3�ϻ����02%>�8����mU7H��ܖ*��!�@��o����2!�ɑ���¦|����B9�������4�	0&�����L'5���j�s���%�-��,�7�B���X��%`�% @���W�6K��Qcر�f�v�~1�/�N���:�I��ե_�t̝�2��M����p��Y�y([�0�
�f��J%	^�Y�-� d������+zi(e�(���y@��MQ�gT�����<�á%:lS��[2��0G�*QG�U0���	��C�M�����:��tun7���IT7	�A�UD
��f�U-@/ ���(u�����,���,
�k�q;ʒHD���Rd� Ζ�YJ��� >!h1E��:�A��K�cO��_�$<x�:�՚Q7�c�>!ms��#ZG�\��m���~���+���Ǿ�a�WG�K_���v�i,o?���|fcc�,�NL$Yy�F)F�鵧��<pRÐ7h ��(�UFx����Q�'�g��0��[(�W�H,ZE�����|�]$.;Ԥ��Mg���eӬ����r���UŐ���f�Ӓ7q*W!"��A���U�s4�=K�B-ҋZ9���>�1������� Ɛ�����H�� ��̃eֿw��{��i`��k->��Tz��.���K��q��l8�����]��t��)R��Y ��}�k"���1��� EA���:R�
�"�B�NϠ�TSWO����yϒ�� ���y>7��O��%�����2��H�a�ےb޲��-��?෾�4��-�\5pzP	�g���:��k��E�P�����C;��+�VZw�^�1-3�@��f�f&�cp�#�-�#�T�!�8��>;/��r]���6Ԍ�I �����GȘ��}�9R��W�r�w�&� )i�e�\Y�kj�	�	@T�����Ρ�O�x�L��~*��Z�wx��}�fG�%��1����f���)˪��D#T^��k�.4�T��t�5�蓪�_|�2��٩���%��j�B�R����,��^�Hk3N�Yx�f�}ã�=2,'�q4{�������3��EnD�m\��;#������z�c:"
O�rP4D#t��0<�=0��@L3��4���FfQ�v��#[��SF��=�B�gb?pH#951*}��t�����ԩ�y�CÒ��VG��d�z�U���+h�s�)�I�dl
�Of77����s�Oٮ ��I��2�y.����,�,��}�b�e;����\Fv��8�tzB~�˟K����'���{噧�S8!�t=�=k�n��Z�p!9�����RW�`8��S�� �v)T=����qn�h]�u��V�&R�L# =�xTzP�G�՝��f�"�Z�f�n�B`�͚�L�-�ӌ��pHG|q������s\'Z-���g��0ͨ@���{H�Q���@gT�K�-�oC
�,T��w1vt¶l}U^��m��!�5�Q\f��xF0	������qAI����wN/�L� H����X�/��yj��n������ɋ<T6�9����جߨ�y���!N�X6EruC��1��<���z~������S�ř`��JӢ2���c���X�����Af��X��"�Rٱ�a�!�֢��:H
j�5D����0�~ qKA��㧾G��"��H��t5��Z�Q�=F���(��5H��E6��������>�7���Ǥ�� x�y,b1�FnզhG��=e��=Vx�P�ϔ���p�4��<8aDih+�(s3�v�,}���k�./G�b����
W��*Sά�:�FQ~��NYت�װ\�a0�:4� ��z�9t��q�|�&P큱�C����}��,!��4�fR�+�j=�׮\�HYt�F�)�%@iK��� ��X%����m,q��w��`��ԁF�k�0K�"#of�9#6����E�:�d(���^zQ�>����P��ڦz	'�1LO�9��J��k��'����VsV����}=����~D� 3MY�D�a�h$ �����'^�������Y���$G\�qc]��kTgB�+u�S����"*v��nii��s���ޝҹq���C2=1)y��,a�FHf|L<�)�� �NM��wɺ�at����&��NI��:=��=z��^�)u�9�%�$jN��ɴ͠�y!C-2�Ʀf�Τ��Pň�e�.�yy�/�����.�����~�۵K@�
��������Mh���XOR������_�x��޲��6��5SG�Q[�h21�yp����ߖ9m���s��H��t��w����wj�Uk��2��3E��_�yʦo�ָA,��*�00E� ��b��w�F��/l�p]� �2� 3��C!��m� `���D�q��=q�g\��b�o2Sf{�������Ir�J�)�G�tԑH�:�Es�P3L�xٟ�ؑC�R��G�����+j�lvg�c������3��O��)���L� `�A�d��W�Ǽ�Y��I��� ���b-�̯Y}ysnq�1�Y�#x �b���ʄ��L�%�5��/ ��B�$s�9�1�� [��	� ��xM�k�L�^���ې߀�ж��L�JE�{���p���}v|�� ���A�M8�Ǆ�an:/U�& @	{Y��b���QM<�f�6����d2�}��cJ���F�À��m���������$��І�� |���(ׇ�n@)�č*��qJ�N�㏎i�-.N�8e;�`��P����{��n.=�<��{{��6f��C������p����y��>���(�� M�Sb9�
���4+,���`7Q>T��ƣ��M:w�z\�Y}U�b<�f�c᩷m�?�$?�?(Y*]{vɣ�=/'��YMw�ni��mz�荡p���n�щ!�;�+k7m��'ǽ�T�T#fF��L3������֨p`�M6�ɕԱvʜ��ŋ1 O��H�*dj:U��n"���`���s��O�����z��\+�5(�M�F�\�H�F�(��ԩ��r�4��Ѐ�]6n|�Ս�X����-��_G�����������-s��`�?Wc]3�Ny������:�@LIks�&�Q:��XP<	�b�-x��sE*5)�hL��fYe��[Y���:md��xD��}�oPJ-���j��k�^f���3o��f9�mo'�"���l� 9�HY��# ��eG��&��f�8��f�`��$���f�?��/䥗^�k���A����"m�s�?.�,�����=�>w.���D�U
�c��Xr4���<�L[3��.�
45��#Fґ�j��Sj<��OO� Rp�~��_�	����#�o3ʎxq��&h!� ��NT�����7`< { �x�i\]j�CP���,�1�g0����U�S�� �]v0��_�դ c��R|V56k�s��� ӥ��&%#/�OR�}r��F9N�A����+|�y?���٬۰�Y5=L'�mFg�x<��햐�s��,&	��j�������\DK&�7��'ا~#���E��  ��?���(x�����{�H2�"��4+B.I�2U�Afu)����bn��̦,�A{Q���� ���Wѯ/�qP��4�:	��Z8�j��Xu���c����O�N螨�ϱd@�T�<K��pY��L�,pұ�IE�,U�b�J���ת����n��r�;&0 7��2XiX��n���ep,z<g�"����dJ^�w6�=�C(E��V��μ8m]�V�������"R��"�}�z 0{^�<��y�����tR�us.<�0ܿW�}�U�hj�%sȤ�`��\�0P@;�����@�WF&'��o�w�y����ь?�Yh�)%Z���[:tn����n9
�,��L5�����U̖h��mg5�Oy��e�VШ���I�5������SD��F륩�Z7j�m��xӎ�-D�á�y��k%��y}��ֵ]Zԙϟ�!��~�V,S'1A���5�IBؖ�V���8@����1�4�0�Z�t�ɨjO��UF�s����yS����[dv	ֲ֦��(G��=�Sԁ��,u;wn7����+4�Æq �_1G���s�
�;J�.�㫯�*g�u#�m�����?]�	���?��>�/ o��C}�B�;�p~�c�=&��2o�|*T8�s��.Y�x��Èt��/�`8#`�|��׃�
��UEtx�l2@d3��2d�ܣł-#۬�&V�N�\�[+t0V��R��8I�A|��l�\�ك�c�!�`e���i#y���.�|���q���3�c�K�h��@�Se��eey���Ԥ	����خ�,��޺����B�l2[(����XA�D��
����D�ϼO��lC�rN�G�S�j�I������h�Z�ͬ�׊�`���X}��5�n��,C�#�IN��Ѳ1(o �B�PAO�,`vC1=5�f�e�l&��ud �a��o�(QÁ��.��=�7X�|�+h0�@��ɑc�#q���S|_�7�GSDy)8湃�-��{�������@2`�G��Ũ2�OTq�#��.�L��e��O�����X'��=Ҡ��!�*.��8Ro�I��	�M� �X`" ��@��Z �yMۇ|��py<�y�Y����L1 x�(��l`+4T7���m���: �b�� �����T���A�n=H�`������^|zz��1��*&�#Ժv|e�=n�p�e� �A�xR3�̀��Z-#M��G��7�����R�khlT��iiTc�r��d�
��6��"�&Ub0�c)5���'#&?���ǈ�q~�\�`6�q��#j�TI�O���de|����M��!�	��"(�=+A����!���%O?�4�·5A�)����sȏ�gg'y�Wq�tn~Mҹi蓋>�!9�S��5�˼�v��k^��aF3˖�V����/Rz,���3��,���ԂΙ2z("�3�(���^p�5ǓAxr��'��Ed߾=�_�\v��A������4����S�C~ء��fX�k�d�2�cٜ`P���
 N}��E�/��vtt��с;Ne����'��6�ܐ郌Ƌ�4���h�G�661n�KE��(^ĳ�S&�#9PԖɊ��ٷ�h@G�˔0��&�'���B~����I C@��`��O�(Y��y<3�qz��(T��bplȀόh�'tok�<�8V�� �'�I,�=�hƀŴ�<�,��	U�@�ᐔ�QN8����/#�b���ދQ�$P�M	U�Q9	���rO��`Fa�������\���w<;W\	����C;*e�N��@2 *��R��Q��k���sL��ˌ��-���pHP�C�'b�S�W���l����^`E�bM
P"����rh�� �C���f=�Ӛ8��}�-�ƀ���KT���(z��2 t�s�]�w�m=�w ���ho`���dtlXb��\��ɑai��&��<�m�hg�Z�˴�F����VC�k�:��#,�ψ;�,���R�f�\@`���}Ҧ�n�M��`��R캤c�o)�m�2�ʻ���R��z�9t�Yͺ=j�g��Y' ~ݤsϑ�-���D��Fh,G���! �V_##��^EN��@�VS���C'�J0��KJm�F�y�-�ɔ���+S�Sf�7�G����FPo�+���V7��\�L�z�q���Q����x7J�K"�	u�,���Kb�D�Tck�̝?_|��Y�qk� ��ꁍ�o��᤼�n��M��2�/J=����m�e��.��N9���D,���X2-?��lX��fm����x�w�N]�:7P���x��e[��z؆�qhww�Q[[���Z��CY$g��t9�����x�I���S�/���ɽ.V�Dײ*ed��QG�E�aJ�4;�ƒ�����bQ�NO���a���~�Zv, �:�n��yi Ɠ���z�*Y�a�<���lܴ����ٳȳNv9��F���.^�b�1�n�ҥ���F���p#C�%���eւ���|F�,zQ�?!����ό� �G�c.aʛ��ZZ[��r|R��������o�۱�j����a�{5\e��h�e`�L�7�.�����#��3�m	|�lc<G�P���iР���X`�B
���L3��Q�>�,�ů(K|T��%�� Z�� �i��뮫��J�eF�ݠܥR&G�5F�h��"�>sؿ#CCl� ����7���Ag>s���'��xn߾��Q���V��%�)�d��"�z��SB��q�S�3H�S� ����:��ǀ� 9��)����iK���L9lYX�m l��՚�&��[�����4@�?uc]=m�	&�
��[�PK;e0/F���M�(^P���L��$`�B�Vp�/���e������1�U�m��lm���^9�mo����i��^�����N��3�~ �:��C�yfo���aY�&�<�G�'�1 eQ-�ހ-jh��~'�qٴ�����x����#1e��>�v���R���z]t�����s�d�!P������2���!��<W�_�"���t�&yHZj�қ���2��r�*����s�c7�1=t�")Q���B9q�Ӡ ���m��n�������/�NbRwT3�,4����w�Z5��P�hʏ>����Ñ1��� ��!��=�Iҙ���j�C&�Z<����.�75x��W��i�h\d�^W�%��=x�I�y�ʱ�M��G,�@'*C#��xg��1��9��Qk��W��`�>u �D��t�L����C�p�:y�͑���b��Q��Y9P��jթ�4���H�/�/"!�emK �w3Ռò#S*����"t������hF� YS[E����H۝����}��[Zi'���c����A�72�����y���A� ���D�I���Ӑ7j�:M%B|��_\)ɕM��7�N�瞗�:v����dx(;z,'9j�� ,ت��?z"mj��I��0�e.r�I���?ʓ(���Iq�z��hmk�{g�O��ֲ�y+�f�"�1n��7`���㰼(�dG���0�����S R��������ՈիW�\a]!���E��=Ҫ�i�R��-z��<�Y�ԛ	L`��ܰɩ��uuI��y�9�
��[�2�?�^�ͤ��7�[��9���������	o'X��c1�ۙ�5��?�������wɢE�䥗^�'5@�({�_*�x��7�
�>����һ�(/�����-^,��[�mN���6��_լ6,5&_�N�k�����G��{�4γu}c��$5#޶��#��e_9��� ؅@�1}��&h�77��~x�|�S����T��ȁ���zvA�}���]~}<'|M����h4L����-�/��+�9蓏�����O:Y�bq��뮻�����z?Y,w�qG�m�>�d@���d�ø��%�"{����ADz٥�6(zzY�JN��u�1��|FZ[�e��3�]G����/>��C�}�{B ��v_��� �応���z�~ܰJ��Fxޒn�Y2�U�eD�j�jB2�;(�RT�j4}P��,����ҵ�-�,�Q������dVbԋ���f�@�2��l���@��)�qe���<�J�&)r�$ U7=L�-������g{H �v"ƅ<�و�����,;@ ٮ�d�΢t�m�֦�,�h�ͯo��;%^� �c�dhxJ�-Z&s�-�J���HMm�n:i�h��Pǜ��'�@�^h:ݭٮF��d׃Ý���_U#1$s�g˳�>#{����WJ8�QI29���9J�~н���t8d�e&����s�%l(ȍs.}J�ғ�<]�62r�K�8���׎>�����ǲ|�r�����-���g���Y����!X�g*mʖ��Ȋ#����!���V����
\Dg�i75�p�P��3a���,?�;�����0Cx�;W^)��匌�w1w�g��&h;1���K�I[�a�נa:3%�g3ڰ~%�ϱ�'��^[/O<�� �R�2d��Yuv���Zr�"����/� ^pp�w�lQg��˯�\�R-N�� ���L���J��{�gQ
��$'{��*��Mk0QW[ǵZ���_�琱����t�[5S	�?��:�nI�����S,���T/'�|�|�}�`eĢ��5C��o�M����B0d�M��W_v��!S�i���_s-n��&:�o|�r�9gɶm���ՠ(D��(n�Z\g��1��㘵O�D���{ｗ������_��đP�'��
����"�A�=��9�#�V,�˾�9�˥�^J�X��2�_�Sʼ�5�\c4�>�3�o�E��g�{Zf�w��d����d�Kk�-GEb�+u�s� �vD�-qc�ߩ��X�CR�imu����3��w�a^~y�lԵOi�̬��,�QCp�e�IjPp�i��ӟ%t]���~�ߧ��*�A`���?S��G��=��c��_�"�?��_����pO���Pپs���!G�ͳ� ���wH���&�w�L�?�����Y�|j��s�&T�B�NK���`�|�;ߑ��[6n\/{՞a���j�J�ʗ/�K�>�=}��˰���m���*���t�8'�5��}j���]&\:_�P�]dVV-[*�-m����h���9MR2Ƽ��h���475ʋ/� ���w4��t��e��BP0�e}rd�X������������ذ��FT�_���@@�4�=�����:R8�;�h5AQ�e\[�Ze��%���N9Y�unֈԑ��{�~�f�u��Ï�$1�r�wD��̙�$��UR7=/��B�m�8<�Ǉe�������P�B[Z�t��40�(k_y�3�E�xC�}�Q#�m}i�ٵs���T��v�~����~�cP�-���n��`�Z)*�13�jqQ�~���塇b|޼yҥ���@�JT#k���P2�U� zTj�aܰa�l�����30���H�,��"W�eVF��c�Lf�F�MT�rU�ܙX\;��u�ֵ���: `^C��H�1���h�[7P� ����挔��M�=g�B���Oo�A.X,��C�P@��у{��'���<��_�>���[o�_��K��?>����ߧ�*id5�LO����;w����?�m�71{���~�������IN��<�5׾��4�nrex� ׏�
��oK����>�ӦJ��=�ϹxL\T��yAR�'?�V־�F~��1(C�+_2�k7����_���g�Rz낾���K��}��v�mr��,��|�袋�����,U���}O.�����t����A���M�|I������gk0�����+RԵzL���?�Ij�,�cϺ�]5�������pV]}=��{���_.��B}�4��?��s�d��-ë���z7Է��.��|�s�'��]�M����}�5@�կ~%����ѩ�$*��ό�cv��m�|�����_�y�;�� /��G�ьp"�{?��|�#���`[�
]��Q�L����>Dн,`X�R$'zFP���C���X��e˖�W��Uͪ�����_��׽�L����ˬ��k��]�ws�As<�)�v2z��� B���a&�����O|�����@��Na�#ீ�<Ka0~�� v��}�Z�(��V�O�d�Ο�}@�S��O���3��#�w���Ϻ��[$Qe��`��ݡg
"H��Ge��C4�X �>���Ҹ��a#�bH�K�cpYof����\��Ԕ��޻g�̭���-���Tʅi�QJF�Q��A�9G	����������i��4�R���P�Pf�U�|��Fs�0� �@V51��*����ѫB6���5�(/8��B�4V1����f����r�����1[������E����lwL?b�F�5*��Y�!�g$���>p�:Č�I�-���+/����ʦW�1;��ye��O<Y�;+�Z��������h�Pm�*5U��`L���dLdfm>s��.Ģafژu5�X%f�6�&�5��/�҈�V�wM`�����@f53��0���N�r��2�2�%~͘�y=41��X�w�~׀�
9�� �Mi�����0:�F�UW]������[����Js��f}8h8_M�$���9���e����=��E��ׅ9V����*P�d��#�=ʯW_}�<�����7�,�xT�uŷ��w�Et�-�_/us�13��f"�q�n��/_|��5s<���5c���j�%����DD�}��`�mָc�X�Bn��w�g��܎v^+�lQ�mj���;��>9�ثh4����1g?5���]�A�ClD��#C��}�N��_x@�$)��7#�(IDP�����ɬ��c�=!�~�y�/����&Y}�ѲJ�;Z8�ࠈ}?N4 �mhd�]W�H�u6l50�:�v�j`���4g�0��=�k���3c��o���@�'���`��=�K��o��o�}�=_�u�Y���7�ɶ�dr_�~� �M�6����k������?�C`���:����_�n�Y��x\m���/Ӟ�-��SO��7Ƞ>������9�m��)�V�p��Ls��[z(�������o]!'�x�|�S���.2��~��u�=l����u��cK�"��'~��Z�
��S�.���Xi��k��G�'��_�t�f��0KG<졋a��E6�� W\�=����o���7(����=��s|nhI����`��	�r�t�a��>� �؛����d��ax\���N�GǓ���h��6 6I}��r�s����4���HW�@�i*/�	
Nj��������|�?}�a����<6�N@�WPN� 4xv$I�5HT2�Ǎ��`��p�J�Q��jQ�4a� �\:A��<d��,Za�$��P�C�'�~L�D�&r4�3�4rvV�\N��p�R�ΏūF�����S@��M$%�0�ƶ�6^ٻ��5�YP���',����=ʡ����>��%�Ռ�J!ʴS�$b�}ON���|�C����ww����VЊU+�\q��;2��)�ca�q_]#��P#�����(g;��7��-=��{����A�˃ %a�T����@���Հ��� �cf���� �*�2���=����k�q��\8@H�B��}��L�RB����ҬN|���LA2�?�q�4/>�����,�\+J�p�pX�}�r�f7�`�ա�٭����	�� �k��Ș�wp�1^y���Q_}��.�uBv�'a2�Vc�%����	8��=�F��Z��E��Z@CvQб��s�� ���T.cK��r�;ϒ�n��̛�Č-M�`�3���M �@���L������o��죲D������a��k�54:"�K���f����z**wP�ۼe�|���t}��ϓ�%�SN=Mv�ک~!dHH�E�L+�q
tT��II����b㨾5��vG1#�`�|�^��ڗ_�3O&'�T�P����3��}B�Մ�}�"��on�h��SO=�^0�Vd���P��GǆyޑXxt���	VD�L�@S�ԟ���%�v�I�X/d�U���gm�F���z��^.������̡$��נf�HB���8%�xl%�ـ6AF��^����[�n��r�O��g������O��M�=����߶}�<��c��A��=1�Y�e������Cs�d^g0e�B5R9*R ���k1k
.b	��� U?:��C6�R�z栄XY���W\q�چ�Sv�*w��z�>���g?��M>�p�o�AZq�[����7����+O��&}M����޷H���en��N	g���Ş48"�F�$ЇڢY�@i@7X��l ������ ��#%���-�~����0��n���p��N�I5"詸R�@?���X��l��+�4��"A^/gs=�e���imk�Q����i�T������&�-H,�W� :�Ň�����-t���AW#�}w��hPP$o6������@�F�+�Եx����d��ץuv+�y��
a42�N�����-�돲^p�9���^�#6t��J
���T�5(H^l�1y ��8uj�i���J�=!J�0*��+�;��=�t\����0��>�N�ȹ�F:1��A�j��򶷽� ���r�f{��ի���^�١��/�Q�cP� a�q/ ݐ�W3�}��T�q<��5�������Ge�dH�*�7�IF4 
{_�f�p����;���xk5�>���%ґ������'�|ZV|�R��G>"k׮Uc_'��9��������4��W&g�l0�	�Q��@={X�=�=�%�0jh5�� ���~ �J�f=�"��0s��{�a��'?)G�Z��#�"��D�Z�>�X�6_����"�(�X(kyI���˚�{�[嚟�����3�b���O��Fj��<�W��c(h��`	Z��\��կ�ͷ�� �C���|�I򽫮���sz���; 2!��P��� ��\���6ȱgX,� ��O��E���� Y?� �@�޵�Kz�C�2&G��# �*e꾁~����V'x���p]v�ed!�B��6>�����9K�_��d��]s�5�Z׽Z����6y�'�]�{��u�9r�]w�g������í�>��Q!����׽&��r�\���j��ΊF@��0��㣲��`B�����ZD�S^�����X�:�:���;��}���}�@ �l^���Q���~��r���~��h!����w���]�M��6�-������:.	�<��]�S��9��Hm8*g��-#P�[�y`4p]v=\��>�q��,|�C���e2=�g�O���oI���~�#�㟗h��-C#cR��,)��=9;go�t���3_�:8���4z���lcZ4	�?��nl�pՐ�߳���l<Q-�7��2)j�8�r� ��������<�SC8cY�`�#�"�Ñp����r���P�A�q\�U"��ل^C�Ω�p��@�l����R�l��)�ã�+D���7"��Tth�1��['*�_�)���½#jO����%��:�!���Y�h1f�e���/��{vHc{�E=t�G}�<��qS2��*嘱��`��+�{�ctK�.��l���,��U_���ո|줜�<�n�Θ��k*M��〚ga�`��(Rv�d�p�x_hR#0�ԧ?��3Ͻ O>��f�r�g�u��(.��G��s�gy��3ϖ���;����3p��{�0����c%��UG��O�4ȗ~��w��{-���ԟ�c�:�`�۫5�6�0p�.;�;�-5 [�����%���	�kh����c�������'��w�w�+���ƴQ3��d�^�O~�9��K"��]�(�y.Wd��4����q�8�Tt�UuR�$4�A���ñ`��	Y��wܡ�|��}��}��[[SO��m[��&�L;5��a.��N�@`���� g�~��VU�-��=���R�L���#�YF)�JfG3O�[D���R���ģ?��|���uM���[@�/=�S�`��^C������͙83�J�x����>� �K���^fn轖��0�YE�>�hXKh����47�ľg�>����ʑˏ��_~ٌ�����c�>)�Ījm�E�ԅ& *Bp�2������:[�lbK
�Gu�Ƹw����o1@���n@u��(sj��)�����`֨��]���?�*����$�nū�h��<���_4!�nج�{J��̓*����M�~	ɕW}G����^߯�i�<��"� �«c�B�S{�q���h'�N\�cO<ì;Q�� �d� ��$P甮�C�}@2z�12H�X��%���aD0 �g:�L6��AΖ�g��W��X�g#px��qM~f�n���)yE�h^�[г?���B�R�X�n��|��u��$��9t@Q$7�FiްPg�?V��H�LdEz�S�}�~���j��)��vgFѣ۷���c�[I&;)Sz�XJ�?(�#����lbU��+�G��BQ�/у�HQ8�Z�񢿅�w`�Y:�:Ȃѻ��C�	�8� H
z4H@�/�}C���.�<�X9��p,L͞L�F�Wc�e��CUR�8[��=j�։'Ҭ���K�|��S�]�C�%�����ݿ���j�5�a�5��&���q�0c���rk�,��� $-8�j0w���N�b�������I Y��Q�_� ��9\"�Mf�
w�ed9���S/�����L�g�{p���$c�ɐ(�������K����O~���I�s�.
+��w@��,�cs�x���):`�aTq[;_���z�|����ڳ��풯��н:�L�14����/����z�PP���A�R�J���NP�)���h�e��n׮.�x��Y�3d2�*���]3��o�Ev-����=]�я�T���- P��
|*h��h||�k��?>�1�_�Z�A��c�&]n�U-(��a 8"��(��~�5O|]s��tO��s�3�y~�GѪ�uI��W��֛oe�<�A�-��4s���,1o�B�Ώ���r�C��������oZ�Tz�e����D��#\?�T�����d�s�2��9�+����A� ��+��Ї1{/b&�&���Z��18�	=�~�R�982.���[Z�e`p���EK%Z@&됴X�2Tނ!b��۲�s;�X���=o��-��3�ɟ���Ĩn��>Ӥ50T�^S��8-�̴0����i�:-]H�b=jKӚ	g��Y��.p���ڽGvl�����XM�K�C�<�����ZE��I*�J�;��h����߀Y{z��k�����:V�h��NW�̫����9p��h ��7�hz�LV��N�LL�R�r> ��XF� ��Й��r(H �����2���%�Q�"c�æ0��g��I�d*��lD�*h�K�/��]�����g�
 �A��1����VIM�"���=�2:��YMU���M��C�ʂ�6�n�-�?��BM���,�^_߹����{�8.�#��K �a��(�>歲s�nyi�$+q�Q�ʓ�F��^�)�a�,$f���!+Cu =��FrCãv��?{���1.�r�̝�PB�2�l���$��-�-_)K��W�8&�}Z�����W��%Gɍ7�!!��;ϑ'�l�Lx��H�F�ý�6,1	�5<>���=@C'}�C2��M����� �CF�.�]3��p*.���c.�n� ?��sv����]�Q��V��������a0����̟���\zTD�$h��R@v���-��>��/��l��Y88r�Y/��Rin�c�}f*��=w^̂�`�(Q?������*"z m�N�#j��d�~���D�ׇ �\��^Ȥ���a��Lv;5ܤV���a��GaZ�4�m�;G�43�>+��9�ʊ��a.���Ѡw�}�5G3�Y��㏗�� ��G�ȣOH�� 3�\� ���h`�F�����$�AI��7��)�,�u�ev����z����@����Mj���/}Q�z�ye��A�Kb3v����f8af�S���~���1_�Niv�LD=F��I=�-1�B�Q*DOy=��(����\��E�PQpw��[d�� 1}(���^{�EG��ɶ�3�jвo�.9����+W�ş�D�����Բ�1�j�NBʔ��U�p�H.Z�̕��i�7P�x��G�e�l�i�7W6o}�<
�i�>)��Ñ]��� j�"�m�t�@zi`(��9u`~��#��2'?A�IN��y��t�鳬����7�3�c�C5`�H�9ZA�d�p�8�H��[��O�'9��� G�~�	�M@���ր��F���)iҲ� ��_t�<���b�<���}v�b��Ǽ:^>�?�L�GG�W8���{߻B��I��5ײ�9�R �BU�aX��O���C�-���K��}��cX�zk0��	't#��24�'����l_4WZk�r�.�: FFF����Q����8^���q��v�<�ee]��s4@#�`M[/k���H^�!��Y����I�A̶��"F@@u�h?���'L����-��<0](��u6�Ȝ���D��c>Q�૿�NHy�Ȋ凓m��y웭}�u��/���VJj� S������S��:S,�ȼ��:61l����w��ꈾϸt��=�-�����;��ӟŜ%���Y���>�}Z�\��XH���X#g*j�|	�u" �@��1����x�4��Cw,��_	H�7�m*Y�{��9{��`�`� �2���GЅg����+V�)�/{���q�O�{��0���'�̱P9����k��7��������B0�����o����N9����sϥN�]����+���X���u��$�	�D����T��� �ͼ9�[j<�؇Ϩs��]6�f�� '���캭���c�R=�-����J2t�Qi&<o�r�������6��� �'OF���P̴Ur����Z�`�4��C~�yr�;ޡ��"���sɻ����~Vv��Kp_����& D٧Z� �N�{�6J˾Gܫ��q��8�J`@A�Y]r�2�ajz��\7 �^�~o
(fu�'�Kg�X�'��Gf*t��f:X��A��ey�.�e��̳BP���4*�w�H�@���Ի�j(�g����Mr�}�˿}�By�;ϖg�����G~*M]
йs��\�R�Qdj"�2(��ԧd��L(���:�J�а����W�.Ct~K �s�5@�ǥ��躡�)��d��Ӡ>��=bE��TL�*C04v�����~I:;�˃���$4��)ź�4hEU2͉�V.���=D�C)[�Q�mD���&���̦hZv�Rh�w��Ǥ�[f�~�W�*g�u����Z=��|A���������<&��؟\� ����cwM?��Ҩ�qQVyP�O#�t��#�S4m4�����8�@9��C��/���0p�����a�L%'�^���#���@Ü�*�P1:����yQ7C����q�~B�5���2Ң�xZz4Kh���'(��B���9;��L3SG���o@����O���3��`�B��hs�T���@��yFd0�6��_vl�#�씑�YP2K�Au��%�⾇#{��Q�վ@z�%l�$�-���ʒe�k�Q�DuT�j���P4D�ôF���xO�d2���`#�7��G�����a���0��D�%J���ۀ�Ȍ��/8\�N���9��0077l2m��%."޼w�)VF���p3ms���4Jn����X{�;�:��h-<��\�9��a��ߣk<��[,��:��	p �g��b[ˎ]��G?��s� +br`F�a<�~�s?����7��?l�r�ʻ����[����w��Z6n�J.��!��������[��V��������İ�]��o��fٶu��5��̼��Qڬ�6�����[��)���C�"�u�������Ih�IP�:F���{z͋k��w�/�.Y,�_�	%"�s�3�:�4K�uG���k��P$�);���@�l�I���F�� ޜ��eÖm2�z'�z����jCcKԵ�@&5�(���u�����ydbD�K�`}���5��e���:F��<���z��(*j���'Sz���c�PA����5h8�dO.{��{���g���G ���f�	�z�p���(�9�{�b��� ����Y�CFخKj����.���!�K�In*#����5����ߞ���1_.p��W]C�MX���Fpz�����ЬVI�Gߩ` eꌋ(wQ��qh����dP(� �+�{_4Q��A�N=ni�o�Sj���x�y���k^0��{���#�Ŵ��sy3��&�c2�IpPH��յ5���Ya]�b3��%���?���
?K/�m�]r�ѫ��o~M���ˬ�P�<��H��8�裒&H�H���ԵN'u��'����K�K8�5�+{X+���7K���U��=A��� R�=ZH�y#26�&�b�C,����L0k�����-��f��Y�Y���-}���I��Dm���v9|�rY|�!r͏~,�P�|��_���[��#�S���T���h�bgLk���#��;N};�U�H��_��׺	3r���Q�p �/!"����d8R#�Cc��*�}Z3̎y(��F��8��9~�hE�xFR�]"�7D$�N��e���PE�ǦL&vđ�Ɂ��eˆ��ŋ?-+��53��f&F��PNkTif�á��p�2���:�pл⼭��YO4� 5��sT`48�v�qMYyN
1P2��uLZ���>6Թ�h�G#���'֔s��sp�)�F����l_�B�p��pO��Cj�{0��YD�f�; q��)��<��Zin��׭��ǭ��F3�(��I�\:�	����2�� ���K�K}K�L4;m��������-ݽ}��o��:$Ḓ�YO>���rڳ�s�#��o���� x�#A������ݺ�S"���~p�~v��X� x��LN��x�����S)����b�a���׾�"��܀e �P�����430#8ҥ��2"z���_���A������=P���C(���w�iPUӵ��_)?��'���X�g8���P�Ek
�5�M�ՙ<I���ߑ�a|TV�Z�j�G>�Y
"5�5p��@��PӁS�S���j@^�o@��Ɓ0������cU���ƒcIc �m�J]v\vX���@АH�[/韍��)_�UU��1D `����u ��
Ջ4��u-ܟ��ɪ6���zQ,��E� D�	/�\+8b�i�tgk0~�y�ʷ��#J�&���kT+�����Zl% h	�\���z�z��L���� ��^uYw�ߤ`5�x�%'ALfk`�s��EPC ��ł�7r���愃*[3iac'V��@�69��Q�4A ��Y����X< ��v�~�\Y�n�465�Рy���GW���Oq|�1^���$�U�Y}��_��-��?�Nbz�M	M,���?(�{�|�S����Kٱw�}QL�Ʊ�9a�{+r�@ ������p/�k8<@d	j(Z�{�� �B�%5�L٨�ԱD5�-������O��6�BS⨱n[p�'����%K�-=x>�4U�j��:�40<!O?���O�P���'��~�LFFǙ���p����&Fsш:B�����"h���R4Z%ɉIl�c�Sup8ʕ-xDm)a�R_Ck�A{�0�a�BL��zI�\ٱ{�Lp�D!��uj�2a.Ԓ/��Y��Zb���^�����+%z�����vI���ׂ>�}qP��k��oE���i�G@�l�0��ZєK֔�L�+F	�1��3@�\�Ku� ��ei8]�w���i�.�����ia�,�T0�����nnn�1��%����M��g���er�1G˪�G�+��'�$+��U@D�NX��	�գe��` �^]�Ǚ��t�igA���G�
��G���	![����]%~�C$������i��a)��	�x��CG%;2��K���~��'q.v@�]�C2enu���k�1G*\�(OC�j߁n�J"����!EE�S�REI�m� p(���~��mۤ����v��9��������J%���s�;zݸ��[�r��ҡ�n�����l�/KΜ�Q!�(�+�Z)
y+��`�e}3h[%��1Y?�˰�n*�֩3#9�h�N~��e��x���^��h��ƂSC�j���v�|�c���}\�m�4���$@�T��5��y �"p@EN����;�zP�8�ly��5<C� �����Q�Bok�8^^�܂1���Uv���k����l�|��op����<�y&+�Y���x�͙u*�P��rL�ZU��5x����ݺ�Z��k���g�u��Ĥ��߾L��_ɆM���Ε�&_���4����{`�V�\�}�jS�>6:� �������o}Ku��5�X�A<�#Uu�c��Ǘa��s����z�9�b�s�^�!��,�N�FӼTr�����NF��f�e�0&�x���F���q =,�K0��LZ�#�ҠQq���_~��]�=�}$5;? �h�t���$
��r��}�">0��`���^~����%1u20��bV�d�:�Z��碟��V,�Umz�$n�H����^f4҈VM~��` �x�ٻ�K3�i��m��n�dP|e�u�@�SB4Ѝ���Ɨ��UEÂ�H�:�|��7><8d2p,&�'i(\`]��0��2Ǵ�OG�_˨:�10�Y 
����3z�p��=W����΀A�Z�=S<�'<ZT;�rpW����k����@���ij��4�~�2w�|Y�d�<������~F���>��p�ҩ���u��u��5�w�yr�m�Șf�>x&S#���_���<p�_e"9����=66��?�u��n���q��q��e����r蜻'���$qDP	�
"�+⺺�U(�����k`]VTDP�40L�9uա��½��<�U�=�������ҡS�����9�G��[���c R"z W9��\��cG1y�de�z�$moO���,�3C4�<��g�o��˿>�P�͊J����ȑ�� �j�WV鬾�X۬m�H�|�wư���%�L�Y^�'^6�������L�=p�B�(�=���X��$1�1���/��ΰ�7��$/3�������|��2ޓ]���?��w�9�qF��|�-��Gmۓ{e�7���jEP9�\�R��	�%j�H��=_��7�0��"ӿg�rT��w�߯�	$��ݣk)jIی���8�"qN���Q��9�2Կ7Vm�1O?�r��{�׎�;�y�n\������oGBl-� �������H������׸ۧ6�wқ��VL�(20�$�o�/���܃��>��X/A��W�c��y:��TT>[��C0EW����r+�~����?�C���{K����_ ɉ��~���%{$!�E\[(��c��g��n�X���?�?>��:�A�F]Ɇ�X�R�n.S��9y��,����1� @�;0É��r%K
�l���IfL��:#9I��}��m��;��MDk0wQF��	JFZS��y�b��i��
�5��������۷�sdO�E��؇"*����̵MnEu]���uvti�gWU�(�
=�)s�f�#:t�b�I/84�F�de��m5ڰ͢��eY��5ω��]mu�>��M��#�G]z����?Ѕ`ĕ�pP��)fe�=�Wa���J��Rd��_��_7�`����Wͬ�AK�,q���[3.q��;5Q�<N:_��ɊE'�@ǭ�Q^��/��$Adk��g����󘉫��<��Q	ܘ���,�zx����5_z�i��]�x�ʼ�v���_^�7n��Y������@#���&�޿�o��?|�X�d���deM-\�P�uw��x��?c����S����gFLo�JqTjc�K�1I�Ԡr��@8�r��j�<~���"��c�&*d�t�����ã�&�
LjF�;�1A��Qr4���� `BNT\���u������p��E��G��OMr� �ؚ��N(�Y�dM}�o����5h�Ԇ	fڻ:��	>T
�������h���d��V?�Κm�������Mo�[zO�R�}�Wx�r�d�{���r�vW�)�����8���&[Հ�����{�v��T-L��=���mU$Uu��߄'���f�~!`�z�ʝ�*�1�����|�[�z�L����iξ+@1U�Aτz���Q��0>Gן	��^��Ai�ft��O�)R�npTM=a��T��Y���F��	��3zh�����H�m%�o��װq�+�ɞ�S#���T�5(u1שS}1�h��pp��q�W��/}��6}�j�O�๪*�;��w������ZUU�19aR��!�x7dZ�5羹���СK�`�+`� 3�ͮU��,��r���.�,sr������#�YFu�9��D��(��t�Nޕ̹B��^qln.�jV��v�D6>���CSC�b��y���𮫯d�U+�T3���q$�puu|���ó�OS�n������O���x��
|1D89da���<|!ok�͂A��a���8��SZQ��"3܉�������eTk��u%Ӭ�|+T0(Ɯ�e�hijՑ���Nc}�)˔Ɋ�N���G?R֧d�)�ssL�}8c����ʘپ�=�Q�)F���k}R::q:i��?��O'��3X�������]g�=�X��]9�)�#N��~(p���8?�����:�?R�e�mr<Tt��G?���
<��$�\�S�4�km�����%!eO?�t9�e�<�ȣX��jmC�>������9�Ք}pTR�������8.N�pm�%��݀�*l��2��̨GF��HR>��1�	DC1�<�
ò�G������&	L?��KfR\S=�G�u׏�����[�09:6��i����s8֖�9u�Gfo�!g�?����U�/58�%E2�ɐ��W9�~�H�"_��#癕�0 f`�z��R���J�c�E�|;�&����j���]��[Fn�߹�V��_G��S,g��۸`����pDs��HS2ƾ��q
��B_^�w�HB$�8��|���
c�7
j��`E��Bes�����y���eD��)���N]�W�,��ZŌݯ�Ԓ�b�V�*���txpHlVѴ���,��-^xV��&(2�"&		?�(���X�\��[���{��ս����\�/5��-*�����y��	��6�N��5k�/���K7s�4��I�{?��?��$]��$����rՠ�`*���t� ���Ρ�ŷ%�K��n��Ѝ譊 �/(�e���hE� �ő��'�]�{,J>�9ڏ��G����t�;��O�`��dˍ�����@�B��itN>i>�\y��>�>�tC�T��d�A�	���|c����X0g�fC3$<��g�'���DrE�s�r���64�4�)��}:qn������� �M94�Tcw�>���s�75:���l~��A\á�r�d�Uⴚ�Y3�fvM&5���#�se��9M�7�90{f�94��`�̆�Y�y0{fߜ΃�3�y�i�h٘��>����}��9�Q,[�L:�d���gP��le���@14��3��&/��D���e��~u���/��R	:�1�y��<���r��J�qC*l�B�����r��z����g圞Ew�1CS+�5)AgV��k����DL��K磉�m��k���
��9d��dQ�'B*y7o��5#p������Nl�*�{�ZɲJ	�/<��J��ݥY|8l�ˊ,��o��n?�%n"�����T�1�m�st��f�T���GK�$;��>Q���K�;{�J�C��Ɉs��t4T+��Y���~,�}u�Ô�/���4�E�P���J�� �:���#���JoY���g���-u���^�\�K�U� �c�ԃc�M�=�C��ʺ��b��*�u2�!:ݵC��
f�]��4��� �������N����c��;P^}(�X��^K"�T�Q�k�|�̵�ql��O����K�z̖_;q�}n��?�a��T�$!׆�oR�-�W\P�68bB�dߑDR7�F�Ł�iHTW��ѹ ���^�B����?���oÇo�;<��#x��ǵ�Ñłe@����^�0Y�J6���ϡ�~ϛ�}5���y
Vi!@��h���&��\���DYؑ��� ��04Ѝ���4��ni��ކ��c���a�n�p�؇G18"%Q�1	eq0�c�8�Q�f0kr"V��w��������,h�hX��b9�F��Y8�������ڶ�f��s	�A�Ēj�G�Қ��+��(��~x�b^'���8���;K�����E�$	�LI��[4�*GNAMD�s����я:q�\�$Ka�_���S��С#�9�$�dV��ݥ+tn�P��N[�N�y�c�&Ӳ��K�>ȍ����ϥ���{��0K��'���6f�4�wK�,(g2tc8HB� �����+�&��h\�ro˵d�r�����g֠e�$,����dťx��?`�������a�D輇�j����s�M%�<$�8e_M*�i���G0a� &y�,$�mV�H�9YOpY�^�d�fG��#0�D*Ӊ�U(��Ȍ�x@/*��za�y=�����x�k]t�CA�1�Jո��?��v,.���X����\hϒ���W��u7|��%]��Sp��?��dg�8C^�4��h�ҽv���;T�;�kwn"j����,� �����r���6.�����<�s�^Vh����}���ݽ��PF�,�g�z`<�����J��Xq�=�wd�SB%jλ��3� �K���>f?��j��19N�:9��j�z�uתwPv%nz�*��UY�dt��y�SP,F�x=J�������#�:`d0���^߻t\�'��Œ�[va�_���0���t��c3p�=��$����Ν�����۶nW>;�(���O=����z%�� �E�_4ɉ�-�Ѝ��@C}�~� [Z����6�:z�G)��j���ǡ��Ϗ�:�t���[�W�P"k�id���+:U�N�B�С��f��7W$m�w��}̡���]��ꚧ��T����L?jB�O�ԨF{����O���?=�2c4��&���Tg�Rd{<FB���@F� ��d�A�a�������ںJ�E�U���%���
�m���cd�M"��9R	�$h	�Q�OTz��h�q�)Ji�(��ß�&碹�QБ�%s�r|%SO�@X2�Q	"bu	�3)�89n���}�g͞������#
?p#�ӝ�1���\Qe kt�$eQ�ב�f�t���i����zH�qR�r��sb�B�s��ז����?��� ����q��Y2��W�O �F��R,����f��I;Z][�dRΘ�x�c������ŋq�Ec��X�n�����v���ͪ���!����vu����	�:P��q.yNALL���b���V�e-V��{�a�tu��k�EU]-�؃�p�y�d($�q�Q	W>� 
�3���9KGAgN�\���� 5ȶ�|��N�o��rFq,*{������~��?}�<�V-�1}��7Q��p`�+��.ߓ:S1+�k�e�>��������T�uP}��d3T���0NO���f���alt	|��'{��bO�Բ�6��P����(}��bO(ϪK_����1>5�qT����b���l��Y{�1��^�o�iy񀇘g&ȪaXEA�eWNw��ۀ�U��P$�!�F�?� ��0і� � G1&`l�T����h�9����L%���Q͚�L�m\s�mV��8㪟��{���u�J���r�s44�b?) 3({�ƛR�K���S*��� eXwx�Lx*?~H�1��Xΐ� \YR�[3?�퇨knE/9$�HT�y\o$��0dB�3�If%��d@�u��I�nٗ����uO��ΟիQ�$�XL1д�涿��_�Cwǲn�v9f)�!��i-s,1�aeҌ\6E�s������J�l�l���v�5�C���ݘ3E��8ށ>�
��G�(�b���:�![W�XF
$�ye�cb��V�ŭ�¨L�?�B��d�s*�1�I �~h.��Q�J��I�R������8��v�r&�(�qL\�����bɇ�B�B�He��\�0�f�.A`�,ޖ)m�=1[�瑽�%}F���#�ā��>:�љx�Ί�Ha�d��|gTF���̛7}�=E�]1�X��j���1Gsu�t�t�>�����!3O΅��3�j���i��Y��k�P���[T3cTM$:K��Y�{0;߰a���������٫V	׼�:��$<	G+��~J�v��j;��2A��+c*>C�[U׀Ç��?�C�#.�:�VYΧtkB~>�ޮ����C֗X�x��~��H���Ŵ��8u�\����D�7�4wt��ނhU-�m܂�� V>�,�r��q��|V>���`�H<�
ff�ε���\�t܈��g �c[E����df���ٞa��DO>���>��VE��;����h)ݧ:_"�a�V}���BYԟ��\��w�"i�8E,��s�'?a.��M2��#,������W1#���N��&Vt��)]�K���;�
�~��$y*�b?�����%#�NT�0��a[��$��s A�nA�̨�O��z	n;�;����HD�1,��@_���h�6��~���5GiQ=O��d'��m6 S�8�
�d7��-�����-ss���R��}�xԽà�QASY�������4x~�s�8��@$P*�h,�v��G`1�G=���$�L��q��%��Ƃ��O��]��R��{��P欳ߢ��6%)�"6(XS[���K��9��cb��+a`Z�Ԥ��B�%�uZ�ID�_W1H�����+-A���'"Ȋ��
��C�67j;��W�H@���aMt���H���k-�<���(q�&u=h�朱��B���!��cda��J��x1(�7%U��\cdr���Qp�=�P[ia��V�ȁ��N��|�iqr�񶷾].Z=�z�5��O^��@����\����P{�d�Yv�Ǥ�:\y�
�cx���q�iKu�?�ܳx�����ם%�����& ��%v٬Z���XW]����2Jq����ut�����|�|�;�(�d�<�p$����3e�b@"};hX�:�%��Eˆ[��mmM�5;��3��p������������vl߹[��јD�CcxM����~��3}-s��K�4t�9%�0���;0�[����ѡ�����_n��m<v����h �M��N�.�O���R�:*%׀�`<w��=\���u�K�kX���ى��f�1� %��͡ѣ�w.��D��u��{����j�sT����$+Yue�w6��-����`�0�q�=�{�V�k`Wqڂ�8�w`��/��܇3�.�M��lܲ~�QYi�:�Gԉ;vH��~��j�ڎQ�c�j�|gU6}���x"I]g�~ci~0Տ�۶+��Z2%3���jDG�g��������ŗ�i�dr�(-��2j���=�ԕR�~�Jd��y������y�b m�:<3��?\�Kf��2�Nopާ��a0z&�.�������t_'�Μ�)�Z�� ,�>���,���� tfLY�U:�V�vnݤ��F	 gΞ�U+Wb��I�ıw�6̞5�gM�Loöm���6s�N2pOpM�|M (s��+t�Dʽ��8��Ӧ�z48����ʔ�,�V���l��xU��!WǱ����]���:|�Sߐd�Q�C]M�^[�צG�t�qޜ�ZM�$&��rT�#g7y)fϚ��nU<�(gH]C�$�P�o,��t���޳S�a����p�M_�+/�*	Q��l�S�{B�
.�͘���؋�ʉ�w�^�Y���e֬}E���e��O�$
T5��� �[�����ͯ��w7N?�T���/c�����\�-,���=4��v(��?�~�M�7t���ߏ{Xe��7�-��o�z�1�W�,�a������9�K��l$C����@0D^�	ri��K�T�(EO��D6�E2��E�;{&��I֚��Lmm�U�B��V�y�9⤧c���:�44ډ�7#��Ⱥ3Z���Fe�H�fI�܅��[��I�S8�G�����k^0�Y���p,�x������-���y�de-ֿ���$gbGp��-�ڰ��Z�ˆmliñ�bmf��Q�ftcq��ƑN�%���S�wɜ�′Zj��l�iؿs;�D��!U	�s�F_������Q}�c��ݿE�&�y��8�޽�չ�3�Ӎ����Ο���@f�/�E�u~t����u�8v�C�i���QSPCT1GY���3,g�b��*�$���@�ѧR��Pm�<#-ƖZŉd���W�}�|b$��lVcF'W����7N���-Y �|��AA%�+ &�#E��\&k8�����(-�X6�lo�����R1@r�����̩���h׵�I���n���p%{�={2���+YVZ��/rޢeX��v�@��\�^���6��Fo<G(�&K�&�la����mO�s����o9bg��L���|R���<�$3�:��J#�=�,F��3���V�6��+���)N�D�zٶ�������\����M�gx���E	�Y����]x-��� ��J���$�v�[qݵ�5�V�P�˩-���}	���Wo�"f̨šC�����?<�V\|>���7��*��}����J }��$�o���������gp�W�"�+7XА@�W������R��O|�S��7�͟�,.��g��e����ō򊊗5k�d*<u�j{�r���G~#V�|������{	ګ�\���1ي���(~���]�"Nw��sTWE�_?�6���r�w���	���W����Ќo~�&��850�9���/	��oaӖ�:��x��?�[7o��T�?=�0.:9n��K����5i`;��M���*5\�l�0���w��;������G>��x���j9�gu,լ7�i��23��m�S}����O~��iŊsP_[�mr����=E�*�*7�@!P2q w��Q\F'�f��e����z;:Z3�1�<�N6y�����8����B������F�����"�<`;�WG�{i���������?-&:��"�X�\��qS��GX۲mB�#�u��-�@ �}��u��Uȯݼ�Ɍ㍉` �8[>"�5dFj�%*Q��E�d�$W!�*��ȍ���#yLn\�ƺJ-��bl'IV���*�f]ԊH �~���Zښ�6�+W=&�F��aqLM��P���U�Yv6��`/z�P��a�"eI7"�v{O����9Cv����%p�SK A^��c���b�IKq�)�a��/"QS7����6�5OE�,��гG%`S�1��$D�ǣa��9D~q:3_�l���C0��ղ��u��Ĥ��a�hѩ:7��ߡ�l��X#"�º������OSG�e�p�͈H搖�3f���6G�XronlR"f���:���#w_��N�����m�A��%�Nz����o������:�uCTb*&��5�#��|��fɏ�p&_�O��PM��4������!�b�Z3���� �^�sD�	[�)�ylRA�R��t��v���8Xm���<Ik&��J��(:%�YY�:R�hgY�"�� ,�x�Ȳ:���z�x��XByOY�t�n�B�X�-b�MU
�M���n�٥mƍ�d�y�K%r�}�dD�r�3Q�'� �ݨ��c�>�|���a���g��*=�1�Ʒ�rg^�ᛆ�9F��!��9��Gn,�o)8��������}k�(I�Y�c���� �-ύC�
S�z��ߋ�	�}�\�;~�s���Z\��k�[��o~�_�Eq�����t����ŕ��|�x��]��'��s�;7�o���8��N���M��A�oQQۀ
�b����'����.|�K_��s%��*��E�li��6i{���Οގ/�V�}�Ϗ�PD�0�?'�8]\˴�6���].���+/C4f��{�����*�t�=`�m��$���z:�c�J�|�٧�g?�j�F.]܆m�ڐ�@�e'�s�ᇻp����e�;��e2�i�-��Qy��ڐn�0�;�TY;�{�~�r�R<�����~&�m���+�����{�zNY7C�A����?�������ߣ�_��8~q�=Z�ɩ7s�*EP���U�$�a��Ů�$Ps���EhoOc�+kq�����g�Y1�L��൸8^gy�go�!�0�R(d.ۼyù�H��o`�2`�Q�h%�K���B������F.�<��#hTn��y�[�6���N��X�RVVK��e�e�=��T�p��(I=��#�6` �񅀇L���h>+aĘ�f2+�1,�#�39-��ŉ�`��ݏ����.XZ�"SH!��DMU=�E�v�V���s$�ւ��d!���٧�0��}�\�����)�')����h���-�ɒ�@�+,w�pq03P�Q:rThÔ�#z�r��;��?��.�b�:Ĺ��m��1.�@{�����K�Ɩm;1i�t����C�G^.��Y>�<?+���!²�%����m�p�)s�~��9��Ӧc�8,ABWo7;��kVK����y��A��#h����s0s�<q�9�)B��j�υ_[[�N�뀙.Ǹ�JF'��^�b���Ѩ��\g���g@BgF��S/���\G���9��+����SiT18V�"�(n>�;ȑ�ȹ�SN]�ǟZ�=^*�%UF�])H����g����I�H�'�CE)��v�)z��!��^r~fvĨ_��ؗ��b^�]��|�r��9�.�+��z�w�1JpfE�,�0#&ǔ��r(�9�al�3��rxZ��'kT��ͥ`���}'c
���6et��쳬�%W?qկ%��虼�zk���X:�f��+|G/�vQʈ9���Ht�f�$�F�ˋ拙8�^��fZEiTi"�N��¥��6��Ȑ���a���ݶMn��P�[���m���:~F.Ɏ�q�B��8��v����y�
\|����[�-���ظ�w��/�O~��Z��O���Sc���7l\�D��CG4��O=�8���J���/`h�_��ʭ�ޫ�BAL��׼���gdoO���֩�ِ��gW���@msl����Z�P�JǴ4L��V~ub.c����r��v-�9�dIjپu^x�}]����=�����;�9����
�{����o9�%�X�`���X��#������_�UO>*�-���Z�������]~٥�`������v�c}/�ooG�D_{�b�n|�#��#��yܽ-��yu���Λ7G3�-[���*���$�~�o���[��8��d�b��_��~�~���� ���7�����̓���a�j�qb����K��*���GNT��_?��V$��N�ֺp��&����m�di{���lIb����|��;���e���>������Ff�an"����,��2�c�"g�n(�+��	qs;�E��ƈ!�EŘ�u6UBq�����w$h,�W��|�QB�Y*U��L�.Y�輄�c,q��4�N��M�K�s�����0:(��ӧN��m
z���B`^0FG��1ʪR�0=<��Μ�-�Ytaۖ����W��W�O=���G�{��(�*Y�9�-G�D�Ӳ83�#G��Li���{t���hk)�X��ѭ�n�-r>3g�m��3�Ş�[�i���}H˟;voAg_N;�l,Zr�ܻ�s�e��m#f̚��\���x��t��*����a�\GX,EUG#a-��AZT�.ҩ�r�)شiSQ��w�:g3�)ׇj{�<FF��}t�O��Q��b"Q�H��� p� �����mo�[��Ԓ+=u�WG�:{�5@`5��?�:���lC��4�Ռ�t����bFP�s@��Qيs��X�A9��V?��}��j3}�Li��56��A�P�'�Cݍ׶����<�em�5hh����=�P]߆��sL.��@o
����[L[��5�����v���A�� �|�8i�����9i3#�ε�4�����R&)�%�/�� �]�e�\&A��ң�:T�$d����S���-��^��|�(�K�R<��#qJ�-~��\L��|��Y/Qߚq,c�,���d/��A�=��H��-سᐂ)Y~^ AX������������.;1���qxq�i�����D2�3g)�����]Ԋ#d-!��l���秞�6�rSs��89s���,Օ���d����� �<�T�4�bT���)STfJ[ڦLRg�j�Xߠ"#�	QǦ�3��\�l#^��l%�by�0B�u�0��Vy�I��a�Ν
�[8
NZ���-ȥ���W�I��ӗ�ȑC��!��J �p�,��%N���$�d�����S�?�=����ǟ�=�L�k��֢ן����.�Ġ[�1�a��J۬u�Ƌ.��������݁�?�.��b���Oc΢���/ߊP�����Nׂ���>(A�/�x�n����Ϸ~Y���m3���L�0����y���w��߬�ڮ;�����i ��1U�؋�Rc��94\aO�N���7�P}�~?ѡ����o�����:9����ず�2\�	����`�-��Ė���/��ı��K�X\��MPtXz�|�u�J�R$�Ք�Gu�2���������1�ĀW��yۣ:�̲8{f,GsCQ��Q����zV�r2ω#➈�H�"�&bz.F#��NխH�!F�}g�s_���⒨Kn��)31*��k�n�7܈��s<������b85����@P�"�YƯGʌ���qy�~�s�A�سC#c�5m�l����R,����p>��Υ�y����Fu�W�z	�����#9�}�o��.���[�{����٪��f�ڊ$MĒ�3g�l��/��eϞ=ꤹ	Y�9�'��as��T��=����`@�Ϣs�����U�T�k����=�T�I�^TL�F�PU���d�+�J�!����:1d��<+0��8"�;�%S��VެYκ�iQ��!f`�(�qʂ4����^����-�`�H�o��v�:������K�Z����E����,X|2��g�̛1FGIbX�+W֑#0���)P�2�h԰l2�y.��D�z3� ��P�G�_�b���&��D�� �5�q���r�[+�f�Ѥ�i[f��Z�+�u�f ���}a?�w�~��y�a<���Ky	��z(��Ql1loZ��z�D���mڋ������H4c$�}
Z�h��2��w��GCSU��c ��5�9N���>k��Y���Ｄb֔�C+�z�m�ڞ!�#���0eR�n�=x�><����۾.�<��Spl�M���얽q&�n �m�Ѵ���h~/A+��}��T�\K���+�����K.���ԩM��M�{@w
{vta�$�u�x��O�>�����X��W=.P��GW� g��߸qN=u��'�ūtJ�����YsuT���WAx�	^�"������A/�s�!h ����H2�U��Οa�������G��Y����=�8����^�a�,������&�/�}r�/8�\\��k����F�\;L\CЀD� �A�c�����3F���p��e��0Z��E�:묀/]�)���.�8���g礮�.143�5���Dg�b�m��r��K���}�h>��#���wJ���0��6v86hs��2�rm�Bq	�Uw<�֋���:���
��a����f� 7�ԭ�I�lI�scɄ��qF<��1�b�}8B�)��I�A6
9��:��'�HC�PP�S(�R�Ƴ�Ӎ���q��UIQF��76����=:s�kU%0gѭ`99a�kSk��g�u�f��C��2�\)Q}]@�Ku]����twJ�٪z����$���O��߲�7����S%��SƤ��J"$���aR���z��by
�:�����'~r�m��kߋ�}���,Y쫛��L+4�^�a���l�y�-Ǧ�[$zߎ�� ��Xq�%*h@'���Z�G�A���K����ϓ(~�4�uM�:�2GN`��~���J�C)F@G�H�;g�<�8vKT��C��+�+���_���D��0i�����ƴ�������%!�����2q�-YC��F��)KVG6lڎ���U��%�rm��\Cc�v���D����w���?b�B)	F�0�&MGP�h��[�h�*:q�(��1M�j�L�<�6�f�1`�K�`��53^b���eHl���l{}/��ۮ��l������&F�2�i��5H�U1�-/1��P'�9/H@���J�C+s�ni��u���������Ş:�Ɓ䊶Λp�^� `�\���z+�<'���$�Ϡ��^�[?.��"��wX����e�$�Aj��[$+ݲm�d����O��e�������a�k��CJT�_ڞx<��6�Nl�9ZZ�d���I��;�,��Y,[C}�d��cr&�1���k�!q�$J�53���S6��ɍd�l-U�T�!����c��݈1�{Ǫ��˔L>��(����Z9��W��w��
|���S��u/��bG�vr�����Ź眉UO����/U����69���^�Ҩ���$-b���qe�R�Q�\l3[�b{�� k\r�=�c�z�olAjxO<�,z6n5��@�Ev��~�U>��/[�������q��?�2�����x�����t�F���Rɞ؀�We�e}�����wH$8���T�" �3�tt$�/��P���KkɅ+:�)�'�&)��uc�9`��9�1N���x�����q��s�{�!�}���1��c�_'Nl(?�
0�<�#��[��R�5L��1.���kefF#22jX�R#�0x��!k�j�m�v,Y�X�59K$#ΰ$�Kz��WQnpX#r'�rl\L����M�:��c m&G�h�j��D�m�g�/N"��	�}=��D�|s;6��%m�T�R=|D5+��I/���r&�6"38U�r�	�SϿ�f�c�>#����ؐ|Π88VKB8"AmM����� �5M��ϼ�����w]��n�n��g��~X����d$#'p���l�_~�v���R��UǷ��~�%B����a@��j	���]��<̾���%��J6ެ�;�͸�Wj H���"�)@�y_�qϸ�|G�'�S__��O��/���	��F�z��Yc�����̍�ɊJv���^:�FF��Xe\+!���a��("���{12{�m�d$e�$�s�t�D͏da��5p4�Q��Y���Q9V'Y���&tS~W�{w� 
����"&ǔ��ǐdH�����;:���`�{30n�˔��RtrF���,��e��/<�����,����Bg,�����R����|0�HO4T��������:l��l�7�ۇ	�ׇ/+�����������;�D�Kϖ��^0,jht��{}��Uē�R@��ņ�/a��˱�9x�g���/��5����{ju��/�c��Y�N��7����6t~z�O$`=Y�Qj��uf���۫����n�iÒ-?GN�&��ʯ�������(��	b�ށ,m����u矇��݇��}J�)��9�ǐ���$�BLd>s��Ū�h�>�YshB�r�Z� v��EXZ!�k�۱e�.�u��8�{ ;�nÆS�v�X��#?�e�����~�3�>_���%Y8�U�W��w�]����dV�J6�7+I]�� $mQ�:r愣Y	���Ir1���TR��q�3�$�#9��7i`�QY�,�l��s�Ӂ���K3��`�J'���9sГÿ��w�{�Q	(ek���I�lC�<�|����v�͹��Q	���6�z���x�`���X5�"�\��-�#�p�_��6��=����sN�sG���ާ(�g~_�x<�rQb�B�M��O�1~��I�X�l%װX��Z�^�9���\���%ji7�z�޹�&X�]��_'�������^��_��#f��(9����j�A܇*�RI2r�g����B�o��i3�XW���c
4��6��+$�g������S=9KOa0Rm�h8��ӛR����1r����G�5��=�)�Iq:bt�}�Q�~�%�͐���@����4F�^�Q	*8_��b��U�2��T#b�=�Z��H1�q���c��jgG\	{9?��F<Y��z^{-�Q{xHٛ|q�!	*H��<'�y�7J�݋�/��k�G^���dT�>�
����i6�O8�g��AP^㌙�>�GZn&��2�=0�#zQ����D�<�$�VH c>���3�dT@��0���#Jq��a�Z�}X���:��p����pRǋ����Vvr�d�s����M��J�O�l��Y��Y~&R�g���/2R̰�U��aƁ�ch���R�Z�]����3����l�U�+���'X�5��� ���0� �_c�g�,?�>$��̓mb��/�@��޳;
��k" f\���V��̛�.��ba]w͵�\�'��{�y?��ļKt-�����o�>�O7�{���g����:l޼Gmѹ眯h�����/)���I͞MѦ%8�o������K�){�����ֺ����Y�~j����9W���x�d�G0�,U������N���
x(wW�P@�,�w%�bi[�\R�XEM�8* .N2(�neU�$6i�1y��!�߼��_�5�*e񦭻��+���*�������/\�G�xR�0$�F���Mhg�/_G冧���4���b�oh���E��O�G�t:���c�	�sx��C�������g	\mlnCzpD)��bK���0�w�w��Ż�}�.:Yl���|�&	D�x��m���O�@�4k����6�k���e;�7;��8V��h��s�31$��Ks�~[Z�'�b�������E/�e��X_��Sj�w��
	�?O|����K��s(���R�I'�����|�������ϰ�9hd��̫��QT�,�P�3��Fᰕ@�B��4q�R��d�7k���cQ}�X܈
d3��0R锞Gem��ʫ(|�e|9��3��y�$dd�X��Dl�J32"t):2��Nٌd�ڷgFdwՐ�=h�j�%�
�V�NQg��ȡ�w���'?�[��lz�5�֫�?Ѝ$���1-O��F�d�r�)��m�22Q%��)��H�UJ��ඍ�=7I�02����ND#	�6;���}��?�!���:�b&A��U�#(��et�/�x_p��$��a�s������;��В�>/��*ƉQL�k�C�'���B9ԁT����Y��lW��ɮ4�  ��IDAT�����#�3'�f�1	N�G�$`�F�f�����m2e:n��pԘ(��v��X����&����E��5\��ҋ�*��}zֲ� �:̮7��ؑ�{���#~���{$ @��lg�Rј�^�^�hǀ��w^�P�s0Zc��昿�+���7~���?����+����|-_��k�XkcǶ|�#7�O��-_��8r�<U�S�����5�*|��O�m��;$�'/l;.<M��갮|�
<��&<���/ނ���j��ѿ�G|�������Z��t�޻~�oq�]w�e�'��|�����4O�(o��>�Yͮdl�ڃ��N9�Ző��4��� �<�9�%[G�6���/�
�}��8&v���0Ϟ"Q���	J
%qow�;���_!��p���Ɲ�ĦD0������J���'�S>������:9�#�S�!ɼ��0���;!{�:}�G�l�\��e�ӟ^GǱN���M�[K��%���_龫;Ƒ�x �h}R�M
Ց��F`�C���uÍ���b߱Y�����cu/.Ͷ�eMRS>��f#�f}X�R2�\*�{��uT���@}
x�g�'�=1�����O��O��=ʝK�`�)�3����,�������rQ��S��:������G�P^u(?~ʈj�m���A	6B�l�."'�=� K��n�Ƣ�X�af���HVS�dq�9���)��i�&�6������T,�Ǡ2�^��d���}ԁѡ��(�9 Q��c�zx|�J�m��`��_��Lɤۑ��cS4 GD�@���,��F֝�4[����_���͵67H���/;_2�9
�#r���(�I�OG��@� ���Y�
BZ��y�t��z���W^,��\-�N�5/�]��{B��^[���;�����X��%����V�`H4\S�)��Qy]��#cz�H���\9�]m��kk+�X7)V���i`06�E���Ft�/��ܔ
1��(|���cޜ��� ���* �XHg�)�;�<�B���������np
,�Miݵ��W{�F�2nU�*[�va���\{��P�-� ���wy�-0�G�Rց�?��f��3��uZ^[+*��٧r�g��Y�}~�ϔ�~�I:��W�i��lJF&=�ঠ��U'� ������?b�kk��A�gd��/h�|�G?�w:|� fϙ��s/^�u�߳��V�O��/|�������ŬYs����y�?8�QY]�'_��W=�D'�Ǵ���O}V�/���R@�2���R�&�zCd�c�\���H�ɚ+x�ì�&)����p�n������~��۰c�.Y{I����J4{����C}����]+h�P���7���
��Ū������ӏ���_�2��5Gw $��G?�]���E��Y��%��ޱe�[N'-���v��Ok���F���+��8fBJ��o�N������:�q�dW�ut�����F� C�N4Z����z�y��C����ǐ�4�`B冹�r?�-��_��|-�sy�W�iTG���y(�����4ug}��'8�"Pn����Й�2М_E��lb��3��?AI�*U���u<�a���`?��T�21�PI�\��ͺϣl���?_�`� l����A"3C��A6�w�R���@%֔�VY�RJ�eO��WA�����6UC�%1�z�,�;n�`y� ���tVAx�`He:��r)�F�F�("M���&)�Kv��pg
�ըm����~�e�S �͌�?�+�X�o�Vlٴ�@�ϒl��$�3���FTI�~������c���fa�Z�ĐA���Tn�&d���k���/E�@J�p��|��+p�Y��֯|�v�z�qDĠ�z�-��f��w��3�\��Ί�nƐG�j�%�����`�=7�R����Ց��&��z{�Z�VW�h#+�Ci���������H?"����8:Zqt���:f��%��fDb	����N�����ɰ2�AY�Q�I*����5UP�Wٞ@Q�������������@פ�S(�6Ԡ��"8�_��7�]>�j>ʳ���������\�>����ް��Z%t�ε{<p�?�6���َ���ܵ���s�ZD�� t���hl���~�hH�Zj8%��<���(�ɿ�� �r�;�����Q�c�{4�S�@�I%+3����r�C��^x�դ�ɘ,��N8X��صw?�8��p���}oE/�ۖ�2@�rt��)�9�K�|�elC*{�ŕk$`Y��~��~�l^���'��0*�k�ۡ�d��a%1�)���� ,{).�xH2�g��V�.�2�;qX�_]}�ڢ���(j��t����?H02Il�V�:}342���Ftu���NƧ>~~��G��S+U(��>�8%l[��-�$B�Q+��D������.�U
��q ׮�p(�B�ع��j8v,�F|��!;����
��u�T�����dE�[�;���#(���'ܼ��N�#�/��2k˲��%ި���č�?=�s���h�r�ݛ}�Q�o\t���}C�#7K�4���������Z�x��X�����."�(XM-eOIl�H��t
��D�g�y��A��,�ΐ�05�sit�-�[%�_BU3C���ϻZ>��֦Y7��x�R��A�A��J���gFh���԰E�ӝ´i���Z)�� :��Q��Sf���S���v�_�?���{~֩������[7�������<ّ�D�c����ӟ�$:����X�-S���O��H�J��-���o���X��;6c���h�4�58&��V�����[��������������]�GΏ�htA0
vT;�e��Vi��2�*�J�c8�BD����R�A��P
s�O��E*K��A������_fń#�uu��}ȣ[���dV�j#��s$��xZؽ{�d��He�X�p	��#��թ �u��^R�UNq��9�_�>�_�^���׫}���s��9`���ʾ����k��a��&�j��rY(�>�[�W��J���˞�����_ǝ�?�;��u�����]�(��Y���Lv$=���p���!�X'�=�{OuE�ұH�5�V��1`������\GZ��Ti0T�+�N�B��p/����k]]=�={&�4�d?�:Ӗ���������H4��F*��+����s:�l�Q�Z>8�F �b_�T�{�v\t�i��3���/��UN�(-�m�/��yܕ��&�
�lke�rL8�e�5P��������b�����}�"0pg����񰂷G$P:m�bH,�d,��}�&�$��AN�'W�(Yڂd�Jj�����$��	��	@8��M�8Vy�j�+w	ߋ`8�K��Q�-A	a*vt`������U6C5�m�o���fQ�\s\H����Xܛ���7*xO�����8�j��O�(w�������N���q9�^yV�;����j�?���w��cw�����8��cV�R�r�K������6G�B��1B�#J`ڬٳ�q�f1�B"�<9�V�3�򣨠p��e���V*����c$x���%ƊTX6N%��D�r�#CE�=��:��ټ%>�m��X�	j*B���G2�̩��Σ��G2��ض���T���J�A�@��<�+nx7��ݎ�v�;��W9���=N��xm�?*��w�w� Wb@"�j�0�H ����������g�y�V|��?�s�+�?'Á�U\沷����aē�j48O��Ysfc���@Ea����*S��n�U�~�k��(��ͫS��`��]�S��Z�Pal�������ث�/�Rf�\�0�L�� �/�M��I�6n�c�Va�g�pQw Rݭ	3g6`��VTTM���l�����c�V�����ÖU�ެ�	{c�Ͼ�-�������^A���U��OL��o����:�l�%T��������g�9V�?�c�g��9t:ÐUz#�-� ˻�,��!���أmZ˩���1>(db x�*D��]^#	���+�+�&�#xO�=3N������ʡ�.���8��� �?��ق9���]����Ǉo�+���y��#�K����җW�u���T���s��RU�R�WR�9�3�ɑ���W�8��j�Y�QYk��]�|q쏀9�B�����OX^�}�9�����*����d�?Yh�k�'�W�}o>(��+����He�bػ���V����|�&�c'��\���SϮ!N�(~�^��7S��dK��+��7�����E}6':���zFr:7�����K�'zL��OT>�������/v_P���>��;p����A��W�:9�h�����s�,?�1���s�{��@pG8�d��
�K�Y_׆�X���*uH'�=��
�<∘8���I	+yU̐E� 9�
,G�|�˚B:�@���T�D�հ$0�\W��a����h��Oy�c�*W>yș����e���&�TԠ��1ټ1Y�C�:c�����3�����ڌ'�� �{���F=O4Z�4	�kk�ݛƒ�����Q7�N��)_�4w�-3)��/}��g+Y�2H44G���{���k0���%�a6��{�3f�CGu4��5qM����x7-��89Ό(�Ѭ�����]�tc�V�4N»��@2�lް�*�hi����=�I4K�Q1�I�q2��I У
p�q��a�r��RS	{�<L�@`�xi���-_D��i:�`y��}�ʐ�<���< �p| m�x*n%�ߓWyR�dm����Re�u�����ms3aJ߾|i�w��]����gF�A�}��pa��%
Y�m��F��u����� �w�qw����N$B!w�@�u��ȞȲ� �B��'d�RE,�yA��)��q�'�1ol�OmEC-�\��%���N�u�:f��Y>߃��QJ#Kb�@DeZm˫�X:v�G>��g��Lt��kN޴�֧�J!�r�rNf�Y%��	
q%���[�.4�A7�G��%QS׀���,��y��ɧR�z}�����	�Drz�o@���B�CFƔ�8���>�ik�m4�R�/�M��o��;�ⵦ��Ҽ��(H6"���2��A�Ni�{k�r̾"�c�$����	���Q����M��-�����)O hUl'�fQ�r��x�e��1���[1-EE�*Q�N�vխ�9ۉN�����}����lNԃ>Q���3�멗�g��M,���n�B�$��r:\����w��Ο� �������C�ئ��Q���tc�,<��P�ǘd�v0��Ū��H���&�,������iɔ�0��E6������F���_U6}V�ɞ�~�� K�O��77U��SOU�I6G��~%cٷc��	
8{Oz[��y�d��9E�6����F#*|RK�j;S�G�D�,:{�%c�����̈��̙7W~n4iI3�5̒:3��@�ʜ�;*�#��*Io�1��o��`a�jL��1�t�~%���`?&O�����
J����r9���R�)^�#4��=�{� ��q�a�l:�w`�_7(Ih���y7k_�,2J�BŬގdR�����jrs�����g.�ϯ��M���:)N�]�Q��7��"8*��-�5)���`̟9���U5ĥ�/D��Ͽ�*b�J�}e�d)������5I, �����L޴]ry��&�U��p��-����k��u=*U��y"�ĸ�F�D=���W�.���D�>��5As���R�=ѡ�\r���H�f���x��-��}�Kx�4�/ū*d��\��A�w�7�y�����BmK.���ؑ�Z��X�А	��ޫ���`ާ>�y�|MYU��V)Xۻ:Q�<
�ʀ�$I�e�5�'��J9��7�1K�|�V$�\�}D (�ĸnjk�p��1U#p3�5�K�83��,_O��1:�������V Oyu�Դ���/�%��Z�WzC��ن�S�U4Fq�86��������by�$hy��:��>܅���E�jPj��6j�_���U^5����K��OF1�1�@�.��&ߜC�f���s^�O�_�9���&�S\�;A�Ҋ��2g6�]��KY�_r�����r���o�Mq����� �<����z%��|�r���?������_N�Q:w%��ps2���H�k����ܘ4Q��X��Ñ{0g�t-�_��t�ؐM�V�3麪&�y���8*5c�,q�3��!lݲG�v��k���z�Z��e�!eA�Nx<^��>�KEFc�\��r��J�e��%�P���D�QGK�TiわUV��gg�_��q���.�T7���J63<0�!���5�#(�kqb /����h�1q���m?��b�ң��K�l��8|�|˓�@�{��d2����I��N!!���V2^�Ⲇ��=��̋�	Eb���#d�|i���p(=����dV�̘J�v�S?t�'/i��'/]���!YL9d�+���E(�h�r`��\ό��&��;zw��iKN�ʕ�aH,���S�6��UuX�a�8�$*%�!aP0��P�5���`ɓ_��!�8�� ũ�l&�H��f�����:�w�v����s�P�_��Ė��9��� �7ãc��e(�L5��'�K_���.�ϛOb)���4kU納�L��o��f�|^��A4V4��'�"�U��L����J�U��UG[�ܨ��RY���Hx��M�Ӣ=aچIU���i�6GmBU�F�ݺx��
���H��]�b$=���*�p�S��Ъ���ɌیT���dmQ�t���S!�Q)�+�ICL��y��2P�q�ެx��>��ce��13mb+%�~s���/B�_��X����}��W�8w�݌xZ�N��U��$�Ŷ���X�J.��(X�2b��ت~�׋e���g��o�1QV!0>����͌�z�^��[�ޅ(�Ə����&�NO�i�ϭ�h-W��G	E�F�a|�^���.Z�������8�ŕ_�(��U�]��e����X��Sa����1���K��f��B#r�3��yf��,tL�Wa�\I��z;u����~��݈M��(�Ecc+Z�bزm+2�v��NuBݒ���"�|�8��.�SG(�K�Ú�^C}�d�}�Ɛ8�dEFFe��fn�ԌÇ�*XΊ�� ���75�����h�<IEC#��5����Hg/Έ�;R�'�yW�㝨kiQC�Va�8ef�Q��e�z	��mb��}���m�#�������cÅ�dr��CYL�7O����G�{�IVV���{+���ꜧgz"0���%�PP֕]w�uݟ(�*��[QAA1��� C����tO�\Օ�}�9Ͻ��z�}�x��S�SU��}��s��|� �8����!?�89��D�� �N��8W����2lh0k�()������$y:9�߁�W���x�N����0`#Gz��A�+,M*|�V��cسgT���ɋs�
�oo��$)t���ȠԱO���qև�.�������xⱧг|y����z��^9�h�KG�����p�s�Շ�H#��ۢT^1(H7g��4YQy��re*^��Δe�E�d�������G�)PZe�"��%6f�s%.�#��P���*�W&0��r���y��M���ِ�7�����W#|l�e���s�D�^u$���w�D����'���� Y0:��dv���2�9�u�}��T��)x�>8h�e�a��<܎�[�7�5b0Km �����k%'q��"C4F��v�~�ȝ#�cs?�O�M�'h�KYeBZ�k�%���م��0"�'��e�t�1�ʑ���l�Q0�	����TwѼ��S�L���M����N3����G�(�Q�%.�}奣О���tKo��\�!H~k2�zAWp�R�n�9���Xq�fx��N����/8�nC�6;��&�R� u�Y�[�mu��0�����]�b���R�J�x�>z��K������h������i�竞�폁��Y[e��C+���r�p<[��9�B�������sV���O���\;�d3���=�b ��%ǲZ�:I!I�*�hb
�\���"��Vr��Ys)�Тw��<�{P��qɍtm{�J�c��M�9T��N�g��O>����qKG�"�D�` ��=���q��CR&�ڡz�g�i��y��!��#4����tx0��G��L�^^��>�A�۵w�ǲ�K��w�~76����~i�X�ڂ�47�:<�ѱko^{s���?xp'�}�y�����o��]-mشy;�9���v�����ދW�\O��&ƐӮ�y����^7IIe�{�����XQj�ȥ���إK���[lټ/���x;ң�gG�<�7@����NTi������sX����3��OYq��D,.��`�Nqv/Ɔ�����ǹ���� ��'�j\�݃ɱ0�^�ĳ		gfM�׳d>�4�ظ��U�M�}6�r}f�Q�~V�X}l��
�[�=��R/`��qT��#(��[��
�%�KĥY�����M���^�N��)�"�ɚ���-(e0������	�Q.-��v��%��C���ũg��կ��PCKu���>�'�x�W�(���g$?~�}�I���_���:n��f2
���+$�����ӓ3�����ݍ��#dD��OK���q?��Gp֙����.��/����z���.|�[�`ݺ5���N���5�\#��'?����o�Q��}�����>�яc��Ÿ������!��8v��,Q,^�K��Ħ�g0h�#����E���
���Y61��ڬ��&z��ʳ�a :�^j�Rܶb4�s�n/Hi���i�{��+�_`�ctX��P�Z擙�ac-ovM3���/��o��7L��P�۠�<,���W�s �j����P�a�c!�9d+SL`-Z]��S��:� b���.C��y��}����7+�a� ?�7ֵ��7�a��b���\�6k��@�R��Z�ڦ�9suվ��p�ݰ�� @E��O�LC8p�aW�>��%�g���Ԅ4C��^=[�5�0���k����ۨ66�ctp�����$��ý}��b�{��o�Η��� k�l�	؊��#h�������/��^��{�IN��llĢyZ�#�A8�	�ԑ�JJ8BJ�opg�z2��Ū�oa��bd*��[E�������z=������p�8<�f2A?y���Z����g��l޶�.��6R�3�~|��;�a��E�3RcK)B �}��`�T�x.~�L�*�qYd8HJ����T���$���%C���t��O�:r���|'�8��w;�ʍ&�o�.�F>-i�$	���G"36�%�io���$y�3�$<�Z��Y�������� MK�sφhmiA:��=��z�f�03c��M��gw3��[R:L�+���H5�%H�'�V��V�_�X�o-��p�V���P��.]�F��S[^>g*�|��}�_�<�Q-�1��4�U/*w�9s3H�@3��w�$b��'0�O'�c����׾��y�n���?��)��Nt�]��_x�[y.�`������Ia�<kE#hJ�����x���I=�k9��g>v� ������.:g������~�#\w�eX��ÉK?����>{�58v��;��u/V�x,���$����� 2���	�{��e��'>z�TPl޴۶�å����ػg?#Oњs��wksƧg�7�K��1wwQ����2�Dm�*�2�-oe��/z����4�4[ɳ�
I��P��Pd���\����p��fX��!��z�bĚ瘬�iP-Fr�L�B��������E�r�w��\`�ռ��U+W>.��R���Ԫ��*�o1�>{�Y����+?�K��K����ػ��|Q�Zƍ�e�Rey�䭔4���(�镞��.�����߻HH�M���4aҙ$y�	Qچ�N�&������W�m]=��H��K
y��v�L�D8�`m,Z�C��$�^S��6nڎEK����(jC��$0:�����i�f�5�ԅ�HH��Q�Ј��w��X�~� �؃e�=�]�`�om����a����TxW\uv�܂d,�Y����`��c�Q����1lܾ/�~Y��6o�0��$�r�|͌�^�^W+&F{��S��gFw'ӯ���Ķk���ϒ��'.?E�q{G'�>�����?'�7�N2Pfq&�R�pLړT$1.��!��X��'�w\���8M�D���l&!��u�>���H�w�t0<6NL��6Bʺ=ݝ�/?�w��8?�Bv�x���E�0%��[Z1�?�$
��{\�ز}��.�9GB2�@�0���-"�8Z�cr������)o (!_A��i.&���B�0�����DK�MА�A�}�(p�ZUK��9�|����(�0�)����o4�C2��3���\4�-�e��<��}���_�芁OEW�H�>�~�L�����ظ�E��^�lٰVZ�|�<����;��x��U��⋱}�2RX��M\@�4ײ�Ȩ{�'q��T�f9�v�KH|����T/��#����@x2�ukcٲNl�̝�j��oк>/��Ȫ�{'�x#6�? 
'���_����^���V+��p�H�w�b^OɈq447�㟸��j�گ��=��O?S�q��{09r�ɖ$�$RSf�f����XS�s�f�F���i�x��Sx���
r�/t#-��U^[���|��[Q�|��R.�����ӌ�2P�U��w��L	���"
CA_Zi,�]++�r*��n"%Z��3��Eiy��`M+�-j���J�������ZG�x���V��@�^G��u�jщj��o�3�l3�	e��Un����=5��M���ȃ���S���$f�Q�%1D6�y+�(O���1#�K�L�|��ڎ={�!��-}ӷ�9,�-����a������)���,!\.-����u�!lڹ�<���]��������
W�`jM�x/\,a�C
�Wmݼ���	>=9��y�x��p�E��w�?��N���p�"Oы��{���$śc%�>�2"�25f�pxm�X'��8����w�9��}�xm�vi�^>��[;�p��G�.���}O>�^x�A��ݻ�����.�x�^�>!��4��^�|��%ʹE6��[��hN1o~�.��!��hxϽ��{I9�����0>�9����Yq״�N;��y6n�N
=�H_�}�����sϦq9PS׌��q:N���!)��Y�ddq� #��~*͈������h�5K�En4��H3=��%������?.*Y������c����F�W9b�;F��-z]�������G%�&����G�˽�6(�2I�t�qؕ��?~���LD��u�M����W^y5����j�}<��W�Is��U �c��[w�\ػwT* ����ʳ۷�(����陏={ ��w��	������q�ݿ�>�۷o'���ãxu��޹��������	����/�A���A�m��87���!�Bw��[��� �\������u'�0_(k?�ѫq�W�7p��o����ں�>����
�\b$��n��i�3��Z3L��Ѡ�I�S0���0#0�L�yC�W�Z�!Q0@���sIv7� �"=�I�2���/�
9�^6�xL����{^��X�%'-�J�z��-�ɰ��#J��?�YLns�׫!֏�R��̏��+�,sQ���Aٖ� ��̀���1w�*���Z��V���Λ�D��O�d+��n!��8Ag��[����$�	�Dƃ�'^U���tJ�����<��N��fr�D��W%��u�_���I�5ױ�NJw0����1�u?�꛰x�8D�g�뱷wP��#�Ѣ�"�0DJ����y���u�낋��y{U3j48wFc(h$:C
��P/n��6<p�/�կ܌�n��,�����w8|X���k8B^C,��E�#�0)ZV�Q2\׫(sI�f5�RYV����F0OX�d9G'�s�A,?qn��7����۾�m�t��B�82:���i2��җ�C�5&>S��&�+�w�̈́����cЄ#�7F�3:���}4�X�h9�dh� H��C�=# ?�j�'��H�(p�2� �|�~/Fɐ _x�����0vKT���.W<��+`Rq_���[�';��'�PЇ������p-	�ֶF���Zlش�l ì0���퀗�.�4M2c��G��,V���K��U
f��
�nɚ�"���~;wȻ���r|����w�{�2e�r�t�
��A�W
^$3A���< L1������lǞ]Ø��g�	x�;�f�^���{�u�=.[�12����Q$H>�JTw�)�03%�9�֮y�/��N�����S���C�?��UG�L��(�O�뮕�z>��@��k�u��y#�\�� ����hRD��]�F�'Ҙ��a9�a�f2�EǼ����o�Nh� p���_���r���K�.î��O�ܢ9�"�=�f��I%IƼ�&�� ����r����|����J��^�P�t�I������J.wPass��?�H)o3�B�"Ĺ��j?��0r*�4mF�c/�]�����l�� Ea�
�7�ڲ��	c�e�<$������C-�ϵ��Sh����GY�%���>o�e\�im�}UB���d+Ĕ{����l�a6�u,I��6�y��q��*׳���#R@8���K�$T	�ؖ�o���ܴ�Ə��	��I,?�DR6��MA<�d���A���֭n��yS����n�Cp�����ǁ��e���@�s��
u��.����f�νؾ��r�B���"FV����1Q����8,��e�9w(�D:���q�6���HK�&\��È��w�]�����}������[���:�&�z�r䒼0���� �HB�V�t��K�1+�X2C���<�$�u΍NQ,[Ҏl<��@&'HB�w���ӟ�y��o�ߎO}�:|�×K���� ��Ο`+�`�Z
)	�J]�Y�j���((5n�z7�>��c	z=n�"Ԑ0��N��a���Q�.Wm3�>q�q���מ�S�n3��H��8�ۏ1����1��d0�{��(2d� y}A�rn����&/�+5��q�e���Ϭ��Y+O�ƿ�pol:,�*�-\C�(�4y�\�� Df�2�u"�ذ$��*2�5���ެ���T[�PƁ�}9!�E(c�V�ס�aܗ��`!��Oʉ��^|.qe)%�K�8Nk�{��h��6C��U	����8�Na(��/'�����x��''-��P?�F�0�Ͱ�\HL��F���%ዤ@h���� v9��I7 Α+Z�hnW��{�3�!ɈDV�gv2vmn�H!���ƕ3Yr�� �)I�C�HG#b�st�fin�]5H�г:)�Ze����`ҺF?&�&$�ewHV�zI:���+���#C�����������N:$Bk��й�C rLj�A2�&�T�
mr��-kL����݌Y@J#�P�Z�1g!��Y+�|��E`�:�^�:����"*��%%k�茮J�r8S��	{��,Ԭ��*��-X��|︪&gS�z[u���]m�R0��u����f�y�R�*�[%ʻ4�^m��͛W��u�U��Ŗ����>�� 9���[)Mu�`Q�hf��;{�R�J��E���^��b�n����{$o���SV����؇C�F"'^��2eYΈ�^R���#����l�0��FT�+�j�&�X�9�ӊ�$ν�]n�C��`���,I�0d��U]=Mh6���f��è%�T��btp�=�4n��p��IN�����c]��w�"!�VT�vaQG���ڙ��db��2W4��c$0�QRS3 E�i���?D���^z)�]�F�(���8���lڶ�ƚ5�x�9(������۾������Y�y2�Dw���&���q ���w��� �F��� X��;���mh�>j�����\@ {�yc���jz*B�Uy�!�D�V�[�L#$C&�R!?=�<�*3)!aJJ��;�ϟ��;�hn�����M��׭���8O̳T+�p���Ͱzi�lUXѲʵ�_i��O
�T�������z��{�ئ�m�^�}u^��f�0�&�T^��9�:@�1 *��a��n��'-ü&�Q~���Cx���i.kH�\�-:>=�L֐��B;��81�M�4U�mY#.�#&u�N2��ϐ�DU��lZ�8pS4��S�O|� 99R06�g,�4��n'�!J�@�)Hk(&%h�>�I�GF���I�,�y��ւ��T*��Z;c#d��E47v��>�_��7����;�����k%��3�A��&쟘����\5G"��&�l,>iS![KqN#��q��5͒��>��_p���G3m뼳�:��~+�7����
�kd攏���'�):w�+`�|֦;�=fӎpUo��+�j�mHr�f�n�b��)�P�H�<�^�X�Ҁ�ʱZaj��4p������j�+7��ˢh���T����F%h��>Uɷ��ǵ�e���
=!7/�l� OԫJ�87��&��p��%�ֶ�&S,��+d��L$.S���]X҆Gȓ����0��JM�a�'�+gz�זzdvP���)ʠ���\�S��|��FHq�t��u==1)�˕A27��]�_��Ex��M��G�#/������h�#%����#���^�ޙ�i�:}�%o%G����y��l�E&9-t�\��\���듅uۿݎ�}�����@�7�8�%�7<�â��d^n�P��!�P�;~%1���^pU@6��t&���x��]t��$@�)d�����M�����a�� ���W]~�D8���I�A���7y�:2��x��g`������b*6��%�POF�t*/-t��
H�b�� t�ϼ���[p̲Exu��xr�+�E/7���lJ�5��	�Ba��BP��+[/s,�b�#4��ޝ,+����j)?�׬#qfWsI�̒����2�<���5y`�>|�����]���v��m�A�;�@���F6!t�y���tӨ渼M�3j��/d*� &�;�E��t��̨*����cC#��_'�tn�ʲ �v)z^���ʘ�8յb��cI!O"ӎ�)���a!7j�n���%+�������'S�m�6����>v�196!T�:�]w��{~����cㆵ8�����څ�^ێ��Q�}�\����dZV?�S�f&�E�K�-J�e�Vb���?�
���PH�m]�=RI!
f����1�{ >{�Qf����jG:C] x����^G�]V�q� �+G�J3o�L��r�\W�V�ڧ�⮆>�[Wͩϱ�+eպ���\[����[<Nu.�JT)���;�<�S�9DYd����+�C��z^�Ê�LJ�K�?+����x8���4V���f��D".�2]OI���Al۶]]]�Ahcs��]�St)ᜪa+��>7�G�d�`�^&&S�2�-�T2*�m���g���I�Vf���['0��'>v%���"���ո�{��Ʀ�tF�ym���xuLN	Z<�����Rx�n���yk�1��� <1����F��8�Ɔ�����#u�L�����o܂[��m|�#��=L��0��(���Vӽ�ѵ;D�I䧠��s��799.B�K����p���_�	u������y'�{�3H�t8]5����r~&�Z�q�Ò��p�|���Ni/��,v��!,_.z~Sa\��ϐ�7��	���D�t�#����r�9��%��I���t��M$<���q�}��{I
hj\j٥�=X���gX�jX�l%Q�<�B�� ��@�ε.���a�S��|����9��22\s4�l@�:c�����yg��w᷿�=��o?D���M-��ꄻ�%HY�y���%O�$�P�(î"��j8#��E��}f�ǜ��n��02� (��"��=N�0�$�<ff8d;a*2��P�Dnz�nG#�zSjB_ߠ�ʹi�յ�a2<*�k�a�o�S����\a�Q=��p�>��G�k���TL�6v��%#�n��m�Ž�I�xs��~����>�=e,c�2RaQ�W�
}�����K�����&�
��?o��8gν��0�:�t�����ǎ�HD��UOF9��Q`�L^��2v[�]z�z��� @��	��-���9�j 7�|�Q��n�r`Y�2�P�ϧL���Q�V���;~�Ҷ#o%��*���	�Y߳�:�ty5�VV�4�g�Gq[�>��
ԼfN^��9n��x���q�Oq���
G6����B�3��㡅���d�������kR%Y�[�||�g�\���2��A���k�mLfCf"K�7 hs�`��e'�L��sIX�]H&"�I���:T[C�t��Gq�U��/�����hi�C(���g���=���Nh�-�k�n�G�$���	ᔎ`s������ؓBzt�QO��5W\���_�|�|���H��c������n�]w���>�@s[y$�����Y*޿p13A�X�&���+�˳c@a��GjŹ�[K;c�s/8<؅��H�p6�I��L$&���<�����z2\8��7���$d$a�D@)Ŗt�`�K/����Ź�\����	v�+F>'	g;]k4+5���i48�
��K���0	����)ŋ�� s�>GN��p~��9]�k��U�9�Rj�X��
`��2�S?*�{���*�ڦ��5�v
��μ���0�M�l*(ˈ'o3M��C�=��p�9�9��_Y���$h�8�O_�O�`������ʳWH�I��YCB⒟�*����yac��l
!?�|�Ǧ��K/r�Vʶ��<��hǺu[��?�@�xh�E���Mc�����qr�&W����\�m;�a�>��b�Fh=�R$�Y�%��c`�)'��`/�;�DƤilݼc�1�%�G�7�5#��6�A�}���y䩳1"Cr!G��!����OO)��n|����_h���[�_�p�������<u��"T
�=dE���%��W�����E&)�����W_�B�0�X4)��ˣst�o�-���U�.����`��/\LI�0���x�r�n;�b�U��/!�я ������c����m�9�?��2�N����Q������uH)tVƥ���ɏʨ{�ि�t1�%�f �=,˝�ta2 ���a7��e�����%⤱�sY$�	�����[zk��lh�_~��#���ܵ�$C����1��C���tZ����0E+?���F�=9:���~�.͸��ts;l�$�q^g�8�4<��u����&e~���Ck�w�
w9ϗPm=y<砫��<�"ҙ� ���gP���4�F�$�77����� ��C-yޓc3r}_������������-_����o��O<�	�Q,\|9Fn�x������!(p��i�s��!20��܇�{�A(<��7�&�8-]=H�s�k���ȓ��^�v-�8����-�25�=+Z�K\�ǆۦ7ף���w�	��kɋc0[��S*?�"��ꐊrȕ���%d6\C<==I�T#o)$�s٬���|eC���|�P��DZy���f�.�kE��Q���f-��0���V"�ف�rC��&Lb�`���hX��}�lzk��y
^\�
��<������ H@d�'�����O]q�q��ڇ�[v��!4�9]��DpX���w	��������lݴ�����?�ŋx���������׷���#K��g��J�/���#�ĭ7��X��2l��	;"�Boi'͛�Fd�ǐ"��O���K;X�$�#q4�2�����x��W�{�̺`ؼк�&����xk�N��o&�`������X�� �Z$��NY��J'=�lR�"����#9dՀ΅�ϸ|^�D_��z�����6G���X�m]A��%DaAZ�ٜ[�-�9�Jj��`"q�]l�C�[����ޜf����E)�u~T�v��̡W���>+�	�[��<o�I/A��
�]��r+k%�Nmf-d�6f?��7���*SˉG\z�2heA�y�`C��uV��H ���O���e�Uf�b#�,ߔ�p���떅�{&��/BT�tH���;)ؑ�A	�דbf��tB��ڸ��0�7?lf����D�_V�\���M�{�(tn�!/}j2���{�,���k�Ķ�o�#�~-�_��|�[��#I�އ{_SS38�g>�8q1y�6���I'��K��t���aYTg��xZI���gQӲ��7M�2�dj���4]G �<�Ç��3�㦿�;�wwc2#e6�q2\���
��s/�����k��CG�LM?���E�M��A:A��&�̹��%B�����8�4���7mí��w�|B��sA#�ˍb2�1�W.�g���	Ͼ���݀���}�y�/!AƇ'���`��`����bߞCر}j������ݵ�@H��9ܴF��H�lI��87���,୉�i��q{�@a�qbbL8
��e���Ն��yG�)�K�B��Q�V{��"d�c����*��9�+�KsӬ\yQ>\Fj�.�܄��󊕧��k?�k^����U�?4�Qwm҆$��S����$��>�rJCQ�s���*�θa6�O��"�B��\J�6gƹ��ڗ�`~{ ��q\r�b�<?���d$Ng|^���#Gs�Kkw~{�[���9gt�g�<��m�T��i^�8��/9�����)-52�i�E!���\�	i��7�������R��Y��}�&3� ��Hf$�b���hl��{?�^xy-|�2ٜt2L&RU��J�MI��o���0?-���j�RM����S2�W�a���)'���>��sPlF�3�Y�d��g�z]/���Z�O��N��(*��J�����J��Y� V
��4K�0�jh~�\\)��О*�?²���J��f��H[���mE��rS��b *��[i.^�AB�����T^.�K���ʛ�g�Y:���
��D�J�4y_|����B�Z��G��������T�.������q���+�SyeE���|�����������iX�s�p/���/b%	6���J�z�Iنp�����(C|f��,$D�uݝ�?��<�}8��E8q9)�P;���]yꩤ$c���{��xb�DH�3K�˩�}�ߍ��]XB�����7o���R������Ix�bxl
g������i:IngK�xd
vo��.��D(4�q-'Z*R!}�ɠ�{d�g�?0"=��X�x�]� &'gd�x�.�azܫ�<s���x�ȣO�G���2����݋$����,�Ã#hnlŪ�_��AǼ,b��$<J�r=F�3��Se�~�6���IШ��p�Z��d�Df��F�������EȰ�����x��T1��էla-��m��˜�B�Ô�9z�6]��+O_��O��e�a����D`8C䕳��$�5!��X��RZ 9Ғn�ǐbt;5�n�`�|Km�U�iv���IQ���t��GI����[�kΉO_��ݸ�{G�%
5Қ�eN���)�T|	���w�����^�����7u��I��@�������-���n�σ\x>��e+uтF�۷����;t[t�Dɀ���K��2onk��`����,�#�:���Vq����o�����Q�G��s;x(F���0d<� �1��k��[�]�&�v��W+�\n�NL����zsq�o<�]�j�[g?�cl�c��'���hb51m"KǮ�?��_6�I.S���]��:ʛ�T����
/��$��U��<G���}���x�G�*#�B�<-:W+�����Y*�:>�ޔ���);̺��Y�n��:���e0y��1�H}}�p�'H�����	�^��q�*/�d<O�΅�~���X�$W�ecY�w�2�on>�i�z������{z\��b-�~lh.�j���ؽ{�p�����k��1�;��<�ȟ�_=��uV���>�
�p_]�5l�l"̦&��Rw�Q�ǲ�=�P8�s'�676�A���}R��3o^�p�V�r'���Lʩ��Sc�$X�?���$B�=�ęc!�F�BC�NR��R�O���fx�<x�ggP�ə3��E�����0�%�����2��[P�F������Z��l4/�C��7fsؑ"����i�e8���u*�j�x��'���.=��p�5��܄;��/����g���MȺ|
�Q�CVs"�m9�3b�_�w��v�^3��a��h>��g��� 
;�#E?M�>�׃�i� �w2X��'#�{���`�+YAU�w�~z��+������\�{U_�a�A;��Q�ٴ
�z�����D>)�Ű�"x_��lX31�')b�~�1���ش~i�8<>$�4>�K"$ܺ�ɛ\,;hN�2e�� D�� #��Yyu�qmHĎ���t<CFp����!07x�		'��L��{́&|����[�+����R�d��N㤀=b���t.u@*K���t����ڛ�L�y�뎻�y�nLF��kj��� )�U���KpӍ�#K��'��ӟ����]h� eD�p����x6o߈���FgW6n�"-��i�]�t-�s��Jkeln�[i:��1@K�y�3�J�8��fJ�SZ��&/M�tx}���13=F�:D�\�l]O#T���,��ZD���������z�s���;�$�n�[���n�/�TxW]|�E�.�~3�L0S���mG��;��U*�w2��1U�G�>�޿�.l�pVj8��d*{.;�kEt?.!4@�84φ ��rP���N�8w��<���\|y�mhom�[o�C�<�F��t���053% ���mr�w������ۆ��>W@`=W\��׭����mR��X�4y~���|�4Y�����صe#>��O��{��G�Y�M[&��F
��Gf����������z=$ ��ؐa�K�k�R���)��xw{�3{0F��Sr/�ɋm
x��t��"�'*�~~��WOG%�����֏��j��#^�֨uTSƗHCC��B(�:�1{W��朧U����r��R�a�h� 	e'�+q��P.=�,�ՂE�;L����Ò��$U�n�[x��.��8x�	���sp�Y��g_@�����2[�.x&��{f����W���dT0�]�;��q2�Ô�}Lˀ/�-fp �Xxʫ��bڬZt�(��;�J� ����J�RC.,�\��ő2E_� R�/C {x�_�җ�*@b�=s*n�wl4�o*S�ق�b�p�.]�`�v��TA�	4�Pt��gh���z���cp�߇�?�G4��`��3 �1�e�l��)���D����5��i+N@s�C�����ޟݏ=��9���u!��#�8�T=��S��惒O?�=�����o2NF�[��=� ��޽�ګ���|��O���e<������t�P�-簐�92��;}��$���wE�]��S%�g�Yî(W���r�������ה�d�*���E�������ږn���Wכ��_۷�Sg.}'�Df�^Z�R�ڊ�,Nd���$W�̷�j/ݎt+Q�3��p�׌�E}��S������`�CW�̏f�^�	��̰�e[�k3J���F3�8t���ʷ�Y�si�ϸ�_o�T�BB�
��u��X$Ң��s�6Ց2w�1���,�YcS��	�۵�)eڿw}��
yD<>��;�L�ן��x���$:Z�pՕ��?�)�ǆ��gb5�z��`��U�=�k��0N;��D����}�g���-��BrB14��K�x�C�pl�$�\��"�=>'��q�o��t
��Z�g.��hb|DH ��kA�ᝂ����TS�E��c���֏�Ȍ(�LF'o#
���y%�|
�u���Sk��9V�"AU�H�����L6oVah�yrC�� m�Uƨ�~�;���C��wp�Ƈ�HE146��zf��04:��?�K1�8���4o�<����4�1t�%��OK��C�iS�C�?W:+yj!#�)%"t��nS.7��/���odf�HXA6�8�#$&������.F#WQhU�K1�Vd�R3���U��<;©�Aq=�-�w��u��S�E�l�q�nܜGP�lܱWI7��&�gn��=�<��#��o~CϪ���օ`1�~y��������y�,����$-Ygh̗֝_sIy>.��Ҷ���wlǞ}C��7bjj�t�c,?{��,_rY!���>��Y��BxG�ߍ�^]G�����C�Z'^z�o�=�����,[<=ݍ8��e����d�(�)��{EĤ�pKk'n�{����yX��rR4��0C�+���Nf N7�wg��������U�Vp��rfyQB��) k��܏'s&6J)���:��l�ţ1�I�򼈐!5�H��=�Sv��|�������|��S���H� d1Tp�W�̜p.N�Rֳ�<�RE]-�>����[h£��J�_<����ت���އR��w����(K��/׍1��W�85�,o]�rº�
��%m�U��Iǥ]��/�/\^W��V�����AB9�֖.��p������:�Tg�y�ݪ�Oʇ�GFuׅ|��ᖯ�k'BuAa�rz���s<OX�sh-N
��kS���&q�=?������')�C}�^I�~Ý�b�,>^[�g��2:����Ix�Iie��b͆������`���)pSi[w�񞆜́�׭�q'� �k,��$��5A:�V���i�±(�5�������)�Z�(BW]�7�
����!lw܋\����W�@�rfo�3w%c�ϊ5K�yV')�R��'���C�F��Sĥ�28�v��гp�<�V����~Rklڴ��8�"Ylߴy�qr�9K���:ģ�r's��/&�t+uS��f�.C�Zi ���J�Q������$�1�y_�K3��p��-#�hRks}^�[�WY�e�3�{ke��(�t��=t1�$,�q��(f.Elk��ȇ��W��\��^�x���D�����mKY��*	��>0���id�뢈hT�����$z�9�,�>�/���S���~iR�6�61æ�r��3X�ь���2-O<��'�@��ܭ#/[���������ֳ���Y�G
�|�o%�v�łu�Һb/�nc�vžx�w���!\v��x�͵�~p�,�%g�UⰘ������p�г�R��DD�ϊh|ȳм�>ǆ�]��M2��+ωK�m��X��d&zܡ��~���}�oz��3N8���IA��.{7��(���ҕB�4�BN���EC)�"^-�Њ���ʕ�u�������zN���5��1��1���sF��s���U@e�j(Q�W�����^��M��P 7+�]��к������s�r��l4E+ɔ���8v�ᩰoN	s]|3�y��3y�AR�\��%Q9n���6�N	��˲L��4���!����@KK�dd���!�u��Qm"��;���8T~�E��TQ�/��?�ry䍈��a���&,Z܃X�����zt㗿���o>�y�k��Bchu��7m'Ex4�G�y125�8&F��h!/~��B��������ڸ	!RV���K
j�,�Ǟ~�n�����^)�Ӥ�~���BԪ�qy�V�����Pmf��&!O1�4����&��Y!j�/:S���q����Q�ѼIrɓ�3O?	]����~����Ec�K/�Ɓ�}8v�
<��?�p�u��zh��NF�S��9��sƦ���eb(#o
=#ew�5�R.QЬ��ˏ��HI���fB#�Ԋ3�
���r�VG�J�\td�hqŵ\��T��L	��ܣ4�Y�aYq��VH�|�^�n��ʌ�a�a��	�(%�c��F<��Ә����L9��pМ���9��?c.�4�Z�3��D�QCy��rŠ̋�(Ҭ�����y�M*C��'��7�K���z��/ï���=4���k�s@�E����$.8�L���$ٺ�s��98���4Nk�W����j��0�`����yص� �d�z�x�rt�'����p56�����Y2�kh|�#����A��y���9ͤ+����^x~V�����b�%�ǜc?婗�EmEC*VC8�虛���/�.�P� �S���K�PW߀Hx������7��R�����{e�Cןul��]{�yk��[�����|V�W~V��r	�^��l芁�|d�sUF�{��k�e�U�yW�١@�Q���������7�}Ӆ���RC�j�*�q2�xR��G���PxҢ�scRRܭkɢ4Yl8,��<��5m��x�����4���s����Վ��~���зm�*�m����*y�5�&�}�[jm�}����J��8���w��6�aR��c�Oؠt�z����e���L���C��&/�?y��]*��n:�������{��m��H�p�����=8�wƧ��Kk��(S�v�7ʸ�ƢHE�ƺ�����Uʛ_��E���/zfj�/Uԛ��뛔&�$��)o�pߡ��R�(n=��!9P�Y����%�"$���p����j)�x�LL D^�W��U4���g?�6���O_�K�?��j46-������ٝ>�ӷkn�YUq���b�f<ep�7C]�w�0('�L<��K����I�I�&מT$G�����pu��+��ն��&��K>ڭ�G_�<���ƹQ�e��ߑ7�HD�x��ǟx�����t�^1���\��M��W��$c�қ<B�}S�'Gz�QP���Q���Ŭ��(�}����J�n�I^�o��/~S�����پk�lB]K�9�/vB���*��� n��E�:��Թw:ÑS\n������p�bNҚ��}b���1�=Ћ�]�ho����;��I����ؓ,9��p�g���.A�'������7h[���\��LS�Zۻ���d�;0�Y�\y�ּ����yI��s44[cH�e�f�Eo%���+6��d|t�d�3�ѓ����t.��;t���G�����'�<��Hc��,ӳT��w]@yV\��-У[m��V���B�V7Ա�)ZU�[�:K��j�1{��+,;�Q
"�|�e
�Dї	{_��sɘHxK 2s�f�d����:�۸*Nw�)M0C���_~��%�m#
8�����Z�~ �O8����p�g�'��?�N�1��a1ln)����h�+���1��a�񡍼|�ML�$MP�ǳ�?�yB���?�dʆ'�xNX����y7ڛj��{����d,IA'N>����"K�dj&�y�Mm蘿���M�1>��w�^���?N��1��&�U'ew	��}�2��j�O��F��M���1�5Go��1���w�6�iB�˭WU*B��ܸ!���L��@[sn���8��^=k�����O��#Ct�<�Agp�eW���{IJ���߃��ڂ-��h�'�K��c��`]�;evg$
�SݪUJ�� U�Q��)���JN�d��B��,QD��J(��{cէ[(q�U:
�>X�����������d=����I��H���8�X�d��H��v�{�+Η������sO?�?�s�H���f�f�p�
�)�+�j7TN�2,m��Y��]7=s���9�/�'�x+�<+V��N����k�}�V�5I�3)�,dճ.�U��i���{����=~��)����4yr�8�$&Oݩ9If��\�W�"��� ʑ�l.#������ͦT���p*�/w����S��i�l~��@�ֱ��_S���CӘ��s�2F�Li3�� Yp�#-��T1���^#�-�}4.�]s-����?�ًk���N�kL�r7�
D���|q��ٴ�L���˙u�*s�s��K-p���yyH��%�u�Ŷ��a�|�j��+���mn���A�y�Ս��y����w�;+��)�D��_�yAF[���@e�i�Y��)�,���9,�՜��Ԕ��6��[��Ң��Z���M�Y�}�ž}�0:>&���8r��8@�s	��� :ڻ0o�"�O�P؅��f�����d�J��3be826��>u=�߃�h������uo��?�C(M���#�J	�-�|��W��/���� �ں0>1�^{S��
�lF<e ��������G����ٹKP��W����p�y0=:������5���2��t�W��CW]��|�C�����@�!��}����0��)���@�P���X�h�%[ɺ�(5~U��ql��R��0ϐ���؂:�SC}��
c)��NZ,eGl��t�Mx�Uذi>���15Ex:���Q��v�%�a˞>z�Ch"#(��Ѽ�d���8%��$R��`+.����A�����
�H$��T����69+$��d�B�N�_�h����*�s�@��xG�ck&1�)W�2G���b@�N����Z�92:i�␚rfdR�N�A  ��|9�|s������1>έ�k$���.v�����t��؉�C�+��D􋑤ƕ3+
)����Z4�W�������܇��o����Y>����?=Ec�(���C�,��3�eRBZUC�3�Ksc=y����>RMI+^Ƥp��T��kh�oD�\�\�I�K��T�qf�~�q4��!��	R�i<�裨o�!Y4!�9�.͊�" В��"�Y=òwU6C��ǜ�T��K#��9%�jy�f�]S��bJ����cu��7���|)o�CRO�bfZ ;9c)z�Y�ǡ��é�|���}Ͻ�����~��)]3ޣr�6�e�rf8릔��5��f1I����}��ly��Bwj�w���0�B�Z� ���T*�։����ceK��K_�8���~[��S��m�֬s��?��bg典�A�P�Z3��T��Oܪo��&���<��S�\���̫-���d��^z�O��`C,�U
�=>�ۮray�yK��PL2��=�w�<��s�8����ɻ� �)��]N?8DJ����x�ŗ����ѾL#I��'���3r����j9Ԕ�q����uX�r%�w��$���i�v�s�#�s������74��{~������_���>��|ɞ�X4���,�y'��U�Qο����{��w�(�,#��0�<L�����1�����h�L'�hv1:!<��}��p��g㟿y�oۍ֎$�(��d�8��!��y���o�T��8$�bz���ڑ&�&)��	���`�	�Gd�H�R�Oyjl��O�A��Ŷg���V�BK�[x������ ��_�2^x��ܱO��u��A��p�O�Ǫg^F������s��O�#E�$"����C@�����H�^0zs+	�0��ǥI]�����5`z���2��n2F���FQo�)�
�|���5�Y�}�V�0�4�xw���s��(��e����U���=�b=�58]�,�q6ĸi���;h����SO=_x<ֿ������D��'P#t�R]���i�0_���_��F�[�rcDR�z��'��_SK���f�pR�L�"�E����4�,�aAw2i���DS�l?0@
�y\{���{)�˱���{�4ߓH�G�y�1bH�#�� �%�Pe��=�n$�������R=��q�y�r#���A@�<u���3�uqs�����.��4r28�q��Jk�G�[���q�5/��dT�W���V���#�� t*��\�����
ƃҝ��ƘF��g�o�������`�4,=X����ÜVf��P�C�B)fz��2�T�R��g��+Ƞ�qc]������L"��N�۶t�����gk~kX�h�\-�:��$4�:}��
�gy�s���f����X��e�0Een�ͭ1���2
P����*���/9f�w�c��BY�[�Z6�.��ٌe-�0Jĕ��翪}a���"��p �211!���x�+��g��T�,U���-C��f����i��m��"#��7)d7j<LC1�L�:��={U�?�!+���r��-g����y�i�Ne��Q�i�ߨ"5���zq5F���������_�w|AF���t��ޜ�����8���;��\xB�����#��6��&@
�%�,�����~��9aE:�~�����08�}�c^O;�/ ���_�կa�{N�֦�dƤ�%el��Q۠'믅e���vy1<4���x=��-�@ѩe�i�(���
�y6^��%�nf,���{8��Ex��Gqұp�g��G�HFa<����f����'���ؓ��hd3=7��ٵI�Aw��� �����^վ�U��4)�D8�hC����|�S���G��|E'A�ڕ�-�T�Z��\�ٯZa�67i�=!�y��T���hbQ�eTe�0_��>��v���6�I�PM��L��"p��y�'p��B^m7M?)i?�4�$�g;l��f�&�3���ӊ"XWz�ˡ�C�}��Eɋ��1��3�v�Lp��&�"�X�����Lq���#	�� ��>��=fN=���{7^��/@oJ[f��ǓQ�R�4?�PL� �t��s�Q�vGFR�6�kb���33�q9�G��AG%�@*�j��>?� )����q��q��^�Q�,mC�8u�X�z=F����>������T4,kU��M�g�-yn>g��&iE�f9��{
Խ淅�[��|c~a�ߘQWNi��uӸ�%$e�+�c�e2o�C��kYi�*�����'����h��X�z��t�~�������GO[��t�!�U7�T�("�5k��[��@i�C�շj@6k+�^����R��fy���{���JB�G*���J���B�[� �/	�i�җܚ�&+'VH\GΔ��}�D߱Pa�׳B�Q���\�Y:���؜�R8�aZ0c��X�l1z�`��C
m��b&2��O>�ƥZ�Fci���(�5�2�P�WDf��СC8�o���k`��������p�Gh��q��R�L3������ ��vn�����4l�ER�2��`���y��Hhz�d!�\)un>р����i��T[x4�4��㇏��'W�R�q�!�%#6�&ለAH܆
e������3���}t]q�\��_�%��;
��P���4H�L� �wb~G�9R��.��E8}�2d�N��E�N���D+O;�_��^]�u�w��uZ;�Kۄ���ܢ��x66s�$&/�� T��pASK���DB<��V���om*]4;�&�_h����fC�W��Ў����Y8Z,N���S�1��o�c��S���&��3Q�8�n���e�V\}�54���m���s���2���-�n%uF_�HY:�N��dϐw���ܯ��4�;�&������-/���p��<�q�ٔ #�p�����w߇E�9��V,�|�6�E������2)^��l?�ܯ��������xs�^�OY9�������5q��I�䡹�����9ˇ ]�v>�h�4�����>�V��h��zE�-Z�;v샧�/J��H@iTcbLl��k��T�k�ai)dKgY�쪾�\��T���5yFJ�@Z��&	�Z*o�拥�Q�yk>I�߫�"1�56qqI�1����u(|C>K���t%��%[�~"����_���k�8v�5��B/�CW�B��(�k��EW��K߿S�j���!�K�;�B�ɗ�_P���+*�⹊�1G�	����ǋʴ�˝_*���(BŻ6��4���E�)tk���Kj�9T�J	����&�Y��E0�t&+a��P��Cdy.eF6Z�-dM/=�X��`��t�9�0�MOプ^(
���o�_Gg��&R ʡc�ӊ�I<b3��/~k��n��×����Y�o��u�8U���������hMM-X��-��w`O~Uޣ�� eε�^?ӬF��
j��e�|p`X������=t;�8|��������8p��&������5��r/FgHs��)�]�3�KȌ;D�P�w��;��0�0w��f�k8%����5a�mM�&�1���݊��xȀ�ۃ�z �#�hiiO��q��%���W����������������g�y�Z�{}�wj~�;ڤD�;�u��}#d��y�����ܜG���E9_�Rk}@��Z�G�y�u�v
ZyAYX��ӎ�s�b�qUF����N��:��>�{Q�%wc70�$��CB1�� |L'$@p @�	z7�܍��ؖ�dui�Zm�����s�{gggw%�������ܹ��{�s�sL��[K0�Ր�K�mo}7����������(J���dZ�&D���܏|����^yb�� �|�c�Č(��z�<! ;�B:_Q�J0ƪ���&�q��}Z���/�09����Mrm1<��>�y�Cx�/@f.�׾�5��F^ε( �tؤ�%a̱�i��p���Ϲ��x�܃c�sr-!58
���r�6q�Wi�g���"���СC&�%�7�=����p�8����#���?���HX�ٌ��y��_���)��G�+dB4�&W���A2O���02�r�vI���,G�õ�C]�u��}�֋	U\���FO���/R���D:��
6�n�'��g���e-[���K��~58<^��tny��ț���&������k�}�Z�N��U7��րhm��''Y���?��jVw��V.����v]�����b4\C��ʵ�H�z��h�7�⮖������\��K�$�-7։�;*w��9�^=�;��=�5O���I�i7k�R*b��|�(�8
���&��xva^�q'{p`�>�/� ��~�(ģ�ۿ�[Q��aC�z��ΰX��l}nT���3��,n��V�亟㑇�>��>�߸��<�D���.�S��f��T5�k��G<y�Y�Ae=5;�ۧ!6����U�~:�HT������j`!����g=�"�ҋi��kF:�WW�&¹"��n���l�
˧ޒ@(��G���-=rH��i���������x�A�i!���v�h6�>4��Xg�]ZS	�ȫIn������G�H
����_��=��o�s�#p��gZ���/������G9'�<��G�mm<(	�4�t5���Q��P7���i�bޮ%�h5�:��\q,�����і�.��Uk�-	���i�~�պ�V�j�W]+?��ϱ�g��ʰ,&vkK�v�0�+�4;��d�T�\Ǣ��f���㦅�ʏdF~+sg]���Sh�� ���jB?y�ӓ	����F�'S��:`L]t���9���<o�=/��s���/�y�z�yj�3Y����W��-���O���CcSx䩧��y� �ߌg�s���� �п(k6'k'��.�$�>1�� ���~1Bv#��>�����Ұ���r.�ĺM]x��A;��_��-QL�����^��*E�9U�x���Ӫ��^��n!��&�m�<��nY�9!��}C$�Z檷+������Jݵ��#��bA9�INU1�$Øz(�Գ�����E ܲit1���]��߽��w]����\��x�x�]K�m�G�RNd�O��/�� �j�}�o�c�7*��^��n\�ދ9��՗�9������]�-�z�>��i���ն�i��K����^�f�����D��������'ƮQ_�[��_,M2Ɇv�k�� h������ZiTT��X5�>E�G�#֤9�^�ёy�y��4c���5���e��W�n�L���n^�|c-��T*���rڟ[sĲ��wb\\��l,eab�ˮ�(� eO���6���GG1*V�8-u��L�Bsԓ`�$���/e�S"I2��ׇ�ьh��/@&''�~���^��k�RȦR:���X�r<rk�þOh�1��ʾy��P����|ǰ��b]O�˹#PBڈ�%����(�&f��(R�G"�Tf���"�.?ikS��u�T�i�ET�bn.�MX�zrz���"��8�b-�a5���g�k�Q�l�kU��L�J]��*k�O⟉�p�;�\Y�/����?ρ㝨�Vnj�1l&�)��7�%Zb��	�G��Lr
c�Â�"��| V�h�Æ���˼<�(j^���4~�����@!9'V� POHt�W3�SI���p��'c�I[T�NMqt�zUS2�y�W�z�`�cXL`���ɜ%���o@�F�s1��.�e���%��`B��C�����s78^��/��w= ˟���JG���٫@�kqa
��w:�w�s4�a۵w�R(k�F���
X��u�iC�L��� @�s(�<��d̽.45w�e��yl����洐`ƲcרӶE��U�!�Ly�
�FS�r�ɬ��I2v>3�Bs�ZGA[u�qX-�3��C���m=�^��}U,��0^�(&����B��'Be����
�=�O,�jᦻ
?�~ɳ�Jf�V��s�o��w-Ok��Ďw���N$�Z���#��j5kU����*��͇�l�J�V{\�mnN�]閮�TSz��ʇʐ����S�Fĺ5Y�~��T!�*�P�O�2p�G�hh�S���Z��Q׳i
@����}3�=���$�zj���(�2����JG�J$Uy5�#�7��>8p ��8o��V>8����M��qv�ʵ��b�DJ\�4�����&~��ݚ[[DaGLL��mALj:�Ҙ$y���{0=9��cg9�����c���==5��"!�Ef�'5�������u\��q���ג�|Ny񙱛N&DH�Bn�����(��I����ԩh� c�n�5&�|r옜ǅX��G��.����,�y C����k[�S��2���8�S����ħ?���9W��b����}:���%Q���g��%�%�mwދ@�^Ļz��ъɅY����ȦX��Y眎7�����7݆��Xy>L�O���!�YTR����BǃU]i=��fy��۪ᴺ���G�ǰ���6�s��,�%�VU�N���U���-��8�H4���P�Y�O
?��u���oG�`n��.�t�@E4cY�眀��?d��p�����"6xq��꥗�_�*ʲ �\�,s#J�/�Do{ ~�ho�j���ݥe��8����6e���5٤�
kH���z�{p� �-�ƿ���\��'�]����V��&�����|H�Ȧ���׼
�o} �Ez~�|��("?���o|ݫ���f.��S�!@�,�Z-9v�5��D�z�q|��O���<��7c1[��閯���U5F�&q�n�[��pP}�쪇ZVy���,;�N}��'�\?%��)��y��ː�ya�����hQ\
>�OU6�ͪ.�ճ��S��ږ	sn�@.j���&V�4	df����	�����^����Nϒ>�[Xu�K���V�Xi�e5?�{�}�R��q����5�c-�ڽ�\m+=��H���'�v����r��3���5�]���d���j�ѱ�{��Ӻ���ķkI�jͪ�8�mM����B�^ͥ��<.�B��9���~��E�ݻG?c�yfjͱ��y�+�w�}J@���k���b��z�*��>����^�H�d�UiK�(��i%O�5r�͊�H��g�*JG C4�u�U�b�b�3K��f>_@�Ń�YnD�e&~bqZ,���([/�ɿA~/�����j�]島�,�l��� �����▅Up$����������</��t��b�T�BgW:s
�G��_��9<�l�{ߊ{�ُn���Ø[(�=�\n-#�:�$M�G�����E�^���&��Lj���k߯���;H&�"h�*���:۔Տ1�Hss�<���U�k_{�<=���S���k����<e�uR�nmW{��2o��,�Z��\{[˓���q-?����D�X��'��?���3���A0nX�ȁ�&@|ltx�{q�s�C/�Į]ص�Ʀ=�f�n�"V)jYi��r"���d�k.���7_�
t�	��nO��-ʿ���p�˟�g��A�{	������%�ɔ���� {,���=_j��!�dY�C@��p?��v��m+�sFʹ
E����mV�_D����ø瞝x�姡����X��6�j����絤���GGG�z����se�� �[n���4z����S�:�X*�q��׎���x��x��G�7+��$R�5ϐZA��TÔg�!S�;�j�Z6������n�j-f��$�]K����$~ڥk�#����q�3��R��.�|��b���v���#Ͷ�cN�%�I� ���|��������|jmS�h�&9zP�-ܟ$����?4�U�]�{ܜɉ-�7X)�9�+���Z:v���z��3gOi7���7��N���`V���Ƀ�{�9�Q\���sb�e��D�0�
�Q�ڝL��8��sl>�e�"L�S�Y�,�ZVkŸ���
7+1Qv�`�B0�ևIӨ�j,q�|�}baA�z$@SS\�ҝҰl.���XO�Lo9�>�-'��Y������F��s�R]2���o�qX�H��`jr�hD;��<>��s��Sb��eF�	�l��A��Y]X,�#xJ-�k^X��l6-�x� �#bi��/�3v�|_���7�J������pp��׼���7ԍ�ɏ���/p�o��K��^x9~��_�\XԞ�`!Q��-����WJ&v�g2�XW1�Y�Efn�����b~. h���X�Q�u�>w~���05Ɩ�mh�{O�N"�+-���(x� eQ�������.B�q�lI�\�|�2AU�����ҩ1��#��c��O�<Ib�ͮ�@���H����#������a��i���y����JdD�W�
�)f�+)Kue�q�.�̪���<��w�oW���������˭�����7�T��4^�֙0_��2�&7����*�F�o�-.�ybq���J�!�,��vQ��ڠ2]^��t�?��M���e�oBJ,�W��p�e`.��B:����V��g3����x�ɽ���	�K�h��TUɱ����Qy��f�,źq+��L
?��-8m뛕�(qaN@���8b��13��߅/���%���F]�����x�%�$2��n,����F(�A!�'��;�㧿�	�~$��U��OeM���oǳOq��6㳟�WM���u��ڥ�N�)�<��\����1��F˦�($�!�{IC>6̱�m�Dgd�G-q� p`���5R���Τ��Dd��4���P(�Ch(�TQ ��(cc�PR#���:`�
��pXv7MNyZ$�I�%9.�9s��7��$�b�/�;[�##�rK��e�P����e.��%ɖ�a�/�
�z䔥,w�x����+]�u��۞)�^��,o'�k�����}�K���mU�e�2�?��ֹ�zKݴB���S�NABdƤ0�}�?�;V�|���N}z�2��cВgi�r�G��x�{��!�`ᢋ.�駟���S�x��_��ﻚt���+^����+�)͎��ߴ��ߔF��=Kvbh!�I��e��c�t��d�r)�%��5��_�"��ݏu��-oϾ}����Ռc��E͋�� ����&���駼PI:\�:�"��i��(�����p	T3X��"�O��_+c!o�{�� �L�d|�8�� ���K�Y�%Ͻ �\��O<��]t�>�C�Ī��kt�%W?��uho�aӺQ�%m���We�.׿�0��
̔���RK�� ����s���L{[�X����[T�0�Xw�&f���kEk���J"lDХ���׾�O}�}����7���8��}:��1n�����z��s��ջ� ib�0_;�خy���3Y_�Y��[�+���ϗ��N|�Z�a/�#C�E����KTrE|�������r��m����V�����<�l���1o��>�_ė?�I\r~�ơcM��9��j@�^ԥ�qE��¾���$�%t`KOS!O�̩91GC�82)������N�\��Fs� n��l����U� �(�d���l:y��׾�}�o�i�j�hӦfxJ��g&6�ɫat�׾�_��w�ڷ��Z��F���2�� c6ikf��]�ve�<:|@���ہ�61ed�K2��F%W9�v!&�"�0���_�	���Ȩ54*I��
̨B�X��#��3�E���>�A�)�Dsc:N}=�X̥4�����)�*��(����t*�9�Z�U��=B";�[~N {hY= k��)*�?[v�]�|9WdV��S�X�LU����F>��>6�,����In{&Q��]�0KN��R�WOe�(�I��Ӭ"�����D�?E���X��Ev<��L��f�����C*�<��۪������%��\�UW�VY��[}�>*z�Kw{�uO�<6�(V���J���]M�����2Iv�tڮ*����f:�8����t��D��G��_����g�����5#}��Q<8�K�bv*+\�#�
�ё1����vUN�60vO�H�TLJ09Ӄi�RiN�'>�q�����+��o|�r��}�1��������T��n�@bqQ&{	���x�Gd��0�Ձw���X�7���5�Ͽ������#,�7�����(k/�b�"d���Q�E��s7
 "
�t'o^'��G�s9Ə���O�s^�P؇����U���K���~䭸�������r��]&��(
�~Q�MX?ЋB2���fxeP��� ��D�KU2	���Y���H�ĺY("����"���j��=����}I�YSr��`T��ҳ�h��ӥI]<6C9��8���~쿕C���V`7|Y=�Ĭ��kϸ�q�m�e���X���8�嫎\i��w�Y[��.u�1΄_��״��Z6�.��<
ZbZ�O�/!^��g�8=���qX�&�X�#3�_�#c�2�!L'���hiħ��*6�w���|6l@kWno�S�ny�C�w)��~����D[�r�h�����w�ig�h�ER�]Q0����[��VEM/f�����w�&�uZv�;�)Q���z�lƞ�G�,V���)|����������W^�BS M�&g,o���w��=�?��n����af���Ee'l�
H�BO�X�� >���ų�u:F���<�X0���<Z�C��B��ط�il��I�7�"�tva_�ݧ(c$�u�HP-W&�ƚ*X߳�n=CʫQš�cJU�86#��[�[)�Bv/����w���I���c���/��Y��W�C�;�Ā��#���܁�o����cc�t,/[��ݐ�gSA��h@�^�<1����%#a�p�Z�1=����j�B�[��䋕�b��S(Y��^�����e�U@���?����<�
�M��ˈe�&����Ol�Z�[+]f��WS��$~�8|=Z?^LoY2�*�Y���Ǯ���\u��h�;r�CQ�A��YM򞂘qؼ�y�1�(kG(xd�3����L	��� E��,&�M�O �>����HX]���WW���GT�45�h?�p��b�7.P��鶢�H.&�^�V)�4�M����Үc��,R�x�ؿ����c�֓pˍ�k,�eX��¿��oڐ����=�h�]\����|B�>u�?�����L0���G�1c�ϻ�%�|*-�z\�K�*y�Č��+('|4�G�P�kf������<���W���}w�?��p�M��8����+^~��v���W�?�~=:$�i���q���M/G���SO=�&���>�CC��jGG{Dk��JT��ɽ,ؕ.�ٳG�1'�~ljɬ\wƍ�'1+�  �&PYVD���<�f�����=����,VF
s�3H�spf�S��g��tu-�J�dWL��|�JM&��-��6ֶ����r�v�֘Ժ�\���q�5��������(�vY5�bJ��6?���[��Zp�-�`릭�"
�֛oFP���ܔv�#����1?'뤩I2۳����������Ǻ�}h�9��3�^���E�N��oj��+y�������3��羀��v��z��3(s��2E_��^&�W	a"Mm82~���_ŖM�{�~��{�� k��/�sJ2����~s;�o.<�\R�u<�������plbB�j;
3.���yK��u�*��ʜ��>�Yܰ�6�w���"s��n�����+0�ӌ�c��=�L\r�EJ �\�����ty�-x<Q� �0GDdD"���ܱc�:���7�������E;BF徾��o�<"�dg�v2>~�[��������W��|�����ԍq���o��z#.|��q�٭��!Q��T@ɕ�6�u�`�f~��e2�*4VR"�Z��l����Z���O�����]x�tggg�{c$,�*��g~~:�㉝�=G��Ʀ��rj&}n.]\��|a�R�h(�I�e֫ەT%��]�v��~)ɠ^�/-9g�/_��Dn���*Y��kcl�ѕ����Q�����b-?F#ǻu�{r��9�rE_=��T�TV�X
���n�gL��c�}YK84�Όv[ٓ,$#S,�r󵴨�L���!Qˎ������}}��O:	�G��#�'�O�g?��bE2��"�Q�!�C��\'����NO��z��V���h}�e�>-(:'����*��U �(δ�G։ωe��Z�l2���,.$���G�d\��s�ry�Du6�bflB�Uiv�Z��!c�k����+��%&8[�>�� y*�trˇ΁A%����T�Vf������a�ob��w`H�W�������E�:?��^��E:��{��R�k>Eo�_� ��Æ�v��?6�Ύ65Lf,d��>�_{�gGA�����pthN>�B�}��/��mL����� �����y���VK]}�8����������6�A�3]����8��Z� ��!`2����5�e�.{=8��d����X�"��!p| ��_.�}�<�ʲ��c�ZZu�!ˊa��Cye��JY����[,�tw��o��q�r�=ܸM�� \f������D��IOՇ�ޓ���	-C���������,�Ɉb�-%���bS���t�\�Lb[?T�r��Le��{E��㱧��={���3�)[ry��ᖵU�����܃Zi�r*�M�����.Ě��D������bo�iEX��k����Ɋ�/�� �.j�K9��I[�����	br|�pge}$�舯��䤶l���|��� ���<��&��
��9�W��:��y��w�ET ��c����cW�?z ����)�^�8�O|�ø�SI�m���/�1d�i&��x���^�����2O��q7���f�����L��lr�Xfa���/>�{o{��^t�����q��]��������'O=04������a�W=U+�k��ء�u��j �����J�"p���ku��3���s#����ZR�N���}��s�s�5-���״����������b�^�Ejc� _� y|&E9M�?w�}9 �L�m����Ě���#�1Mx�gYS��Vi�뽀��YY�������zח��%X7؏�>���
�M���[�&˸J"p*K��X�R�3(0q��ڣ���?.�h��'�%룵.��q/9�"�msT��*���ο�(sZ~OQ����:�4̄�8Y{_̢��U��('�ב��{�G��g������Ca( ��"����7,י�����i�D��7�i�%ފ]{����뤐-ȵ��qp3�=44������WLC�@�X{p�駫�Qe�u���֖�(�$�'�g�@
�Cs
�ȫ����I�x�Z�H�Oat��֥ҳ��ԃs����"��iAV�L��a�=!�In6o���`��'5��V��0:�sΏ�lw˪_����*Wk��㭛����|�mE��a�����q�9ޫ����jI�˓�̾KM����ɞ�����N�k*L�]r﷈�DjF�<���|=N?S �͢����㲆�hn�cxK��=��1��� ���X0�X܃p�M<���AΚk1�RF��eߨ U�v�H��ydcvgGz�)�{YS�ZX�O�Uݪ���.fgd�th�"s��qNX��O�]�����
��L���[A���&�=6���VY����-o�
7ߴ?����Ӄ������YE!ΧE+	�L$�d=��;��q�Tř'o�o��Q���-&qp�8v�:Z�PI�>?g�\�j�b}�ǽ�>��6��
pZ���:p�mw�z�)�-��T*���}@g�#��'oڈ{��G�'>�a|�c�����"K�f�0(r�*��)T�yص!�۴�-�L��ۖON�,,L�l��o{�;������c���gp��2�͇~�w���9���=�wd�*��[ᨕ�9@^V30��^"�-��z��Qg�׻�K]�H}g�ot��E[�~9�]}kt�7*��	��߯v����k�����*Vy�X����?��fj���)V]��P��s���:Z�V^���{k���v�Wpa����UK���$0C>���Yg���n�>� �Zڵ����Q�=�4>�EY���cOa�c{���Ȓ�l����"JiH����1��`���7b�w�,�y��WD��L' �f�WL^���`_�
��]ޗ�0�1�%I��,�a�	A��G�o%Z�A��.��]�����E����M�P�O`o��!�,�ydD1�se%��l�O#'��'&C��)!��c-r�M^
��Z#�˖񜋟/���5��翾�s��Uf.�q�:�L�jY����4qqL����X�C�861!�nVX�d<��S(2K��YQ�\����-T������GQ�s%�����.�(���Q�Jf<����f2�+�hLݣL8r����^[Ku������WW�רPW[��V�����ꪲgi}�����w@�j
]?/W�v�.s,��vV��(R�	V���X�)�~˭8�`z2��C�ϻ@��.�x���jk��:�Păb)��a�~����{qF,Q׏Gk�	��D�_$38���AV�?P�s�Mu<�����C^�\����v3tU�ZOd�����u��b$��s��\�E)W��hR)j�r}�`��Tr9���\ǎA���}��hoc�奸���S��;�)� �Y$� c	�`Yݬ�ih�5�&,�:��gk�@��DUqO� "��Ք��(O�</��n�Te͍ܫ�`� ffS��ʰ��看n�V@�z�]!�X�a���!9%�4+���V;q��7����߼�=XL����BH�i�MrB�+���P�*��v$,�%�R�L�W->����_���>����h�v��'LǞ����l��?�g3o�x��2�P|!�W5ϳ���3�c�3,p'��R�v�q����`���쏍��o��z5���k��9�s�j���/�$ˬ.4���M�P�&X�DW嶺w]:@�����ٔ��t�Zs�V���]��%�%w}��-�7�G��ˉ�bi	k�Mͼ�KB�.�����u�)���;�u�6�eB��ك�Ͽ�=���� sO��iB=���yRu�2g��a�SZ��[Io
� ��V���I��g�P$�������}*���"������ƚ��+�+eeƣ�B��E�Lc���f�s,��b���Y�,wa���z��8���пn��s �~��(��^�m��b.����af��Ӥτ�&�n��#�+�x��g��o��������x��6���`��!L��s�Yk��"��ji�.�	�8���S!�ԐX'o٬���:��ٜen���7�9��-�\k�J�#(��bA�!]�s�$@�r+f�j���M[k��d�S��d.&�q��嫻j����]G��U��	ֽ�[�WΫ��՚��"�]�*�*6�]=޽����p�V����+]�|�C��iŴ�+�Lw>z���� ���:$�y�����cذi>���#!��?��7��-Q�m+�̪��vq�LKfry��e�g/�3X\HirR���L�a�Q�X��GP!�0[����J����]%s�r�ͱ ���$�89�#��v諈u���ĒmuiDN���a�2���nS6;~���w�̫O|�j�߳7m���Ț�G"+V����(�hk/2�C`GɹY�Q�_�<� ���pΖW 1�T¬l6�6����O1)N�~[�RU��J%���a�d6��(���^�����_`Ӷs�����Q��!t��z"�:�\�����`�MW�b-͸���W�r���o�s_����g3���]�� �������%=cBR�G�9����Rf��˯|��H��o}��G>��~}�}OlZ�'�v��2E%䄗Q��𔝖�t���2-�ʖ���:���KV}+����Y���X��Y�Z��ěk�Yj;����v��Pg *�:ۥ�,5��]�cm�����2��\����F(ee�Z"to�ܮ�  Gz�xx�&.��D	);P���EA��H�I�b�i9qc-)Y�����(�g$_��#=��Q}���X���L�mE�y������vc~a��"���E-�?!h<��H�gw�EH��&� �T�&�ٵ��b(�c�� �����K��TRr��(���X�mM.�h����H�����l��ʟ�o�� �|��*o
TЧV�Gv<ޤ��G���E!�S�qGR��5*-pv�
�<G�>�&R��Rs6���^r8��6���ߢ�������aL�MMϡ��b���2��/f�bc ��7q����s��՟����C����И�5��6؎#�X�~G��f-�N?K,t�g���6	E~���e��9*e�X<=H��2����hj�W@˔h�{~F�n����1e�b�s�D�l&Re3�*d?A� z3z����� �y&��~�%>���V��x�4$d�_V����v��K�Y��Y�PqR��kUk�⯭Dː)��ot��vs�"�F���=�X.�V���N^신�(�	�m����d��3f��1K�e���xt�U�J�J<5<2�+_�\�*�u?�)ڻ��N��#ò�"c\����r->2��m�Z�i���y�c����Q�iK�\s�Ó��r��0��#��*�QSO7��rF�'��2�.���G�xss�hi�c}�z��w3��Y?��a�b��"G
2�{�ؔ�OO�U��*���M���M���?}������|2��'��Kd'd3)wP#{),LM�#�Ʊ�Q�c]D��R�駝��Zd��L���]Oଳ�+z�Z�n�HH�KM2A��fe����C׺������O����<�a,�������܇q������w��/8?��;�"��2��v�=2�o�h;�z���x04�$^�bZ�V�Nd�ύ��S�[E$�OL?y�9�n������̝��/:2����G������4F��+8A�LV�f��hV�-͊�d���6����F�����^-��D�;T���_8�R��J���7^K�Pb9��zr�v�Q�5k��P�kXV�ᄎ�}>vP�2c3W-��R�Z�a[ne/�~��i*�#����p�}�Ţ4��ڛ<�Lo�n���n�>�
�Q$sb!��y�28��w�ua�9t~Q�Lؚ�M
Zu�u��o,{#7<;�5��)P��P�����9��ggTA�ejKK���&�}��JGI�_���?��%�oF�p*����`�7���V��t��y�H-&jnc�b����s�5�t���$�L*���@��<���w����ǰnp<$]�G�-��ڟ}vnN3���	\������at�blj��_����=�@����v��F ڂ�v<����M-�6�8��c��G�[�ǎE��E�y�������$ ����F�V~�v"�ԃXs7����'�ގ��������D)gd��mL�̊\sY��Ӱ5��9����N�Qτ8�_�T"P����/
 �1�h|�g�b7O�S˩i\7N{�M�2͚q<�䫮����%�J�?���a���7\���m7ծ��be���=Nb1-����ce�K{tr����e073���Z�����/�������u���S��##���,>����e/8	?�l�����+�ϻq���W�G?�)�r�)���^��q�>}��<\}�;�r���n��������l�͓���|��·[nًk��g�{>��w`Z�ϧ?��شi#���+�Q����ۅ���w����ħ��ӻ��n�6�����]�v�mX����"0>!�@�m��1NN��b���݆�]�G*�EB,�HЭ���X����`Hk�]�6o��0��|F��i���u���gIǾ�� k��q! k�gp��&,,�p�^(묨Ի=�R9�׭^9��|��kq�g+���~y��GhkmG�D.I�"����H���0��(��n�ie�37!P����.g["�߽������b{����gnx��}c3���ʛD��Uc��?�N�:��L6ザ�^m��ǘ�Z_�>��T��K�y&n�g�lW��|-�]�^�X�����V��~ո�D+�J�3ԁ��k�#�����q;t��Lu��ܧ�����Z�[�|¦��S	�r�H�f/��1��\"!f#�CJ��/B���/�B0ք��y�u��<Z��4�ҙ�)4�"�"_L�k��B��@n�����HD�T�T���4EE�K.�Ё=xz�c8u�VQ���^X0n�b��c��=�b��C�[�c�NM�����9�:7�3Y� �xT=]u�>��-o{� �&��}�C���o7~)V���'U�55����`�c���F���wxB��!-���p�M����C"��y��ZƮ]q���޻^���f0+J��2>̔e���}��2�{����׵/�Æ-��nw�FǓغ�\���[E@?O�;*���5��P�[�]�mH{��@�Rgw�nP���+C�os�zTѰ�KBS|��3��_�Gk$�Zj˸�>_���n[�ڝ��WmM�.Qm�i��5�����R�\u��%�PszS!��� G�RZ�+���"+�n�7�o]�]����ᡇ��������a��h\%�ZzTF����iFK�3���q��D� ��@X&����X��m��F{+�|P�J1���$Gٲ�_���
�Z�w��mho#4�\kK�q�����4�J.��2��w�CQ��;�PXAF� ��*.�f�kF8%[�j�D�bN����1�D���C�ə4�Tl�z:
�"ba�(�Q�P8�y���2?��)Y��S#�U/s�E�������7��`�b�?��Shi�@쒵�B2#k=��c���#�SW9���fh��ۻE���qlb3wܫD3.��4���;����Ɔɞ�<�B�T�m�����7�`��M}s�=�{j��b�]�����`��E�W,WZ�Xo=W��֘��e{�d��7+?_�'��/K�i�l����s�>ֺ��K���|�5R5�^�J��Z��2�Y�v̸���e��2�tV��0���` ~��5]�"�M)�!����E6��g�������&6��5���ړ���׾㓳xr�^���b���ǘ^IiJ�?��t���$
�K��^�i��\�����wzDY����0;9�͛7j�����I����ڕE���q汝�}�Mk����9<A��}�)H��2�=�����%;������+��^������c#b���q��AX�p	R�z�����CQD!:��w�g����n<���H&	����������R�������d��|����%�f� $&2�ծw�HL��C���0#����7�k�����Mv�}Zo˸+W���rT�B,��V�z��{����jB���[��,0*J�� %ψnE�?��`�T�|w|��V�Y��������?�j2B��.��n��$���W��;i?l�Q����@ݡ�5J��q� ���܈G����.��!��wR��&�3_��o㞭���1w�_��q�Y8tpH�[��ݟ����hE���~���
G144��bIr��+�ф�_��&LL��_���[����{����o_�����8� ��x;�6)�}�{X��G�j&�£�������x�'������/|�{�?��dw�o��Dc�F"b�W��A]Ӝ��5�j4��'k�Y16Ƨ���Ş�192���SNވ���&�-����lA���?�t�L$�:thH�Eo}�{D��ٳE��aAQ�|�"@X��BR�SM�n�J�SA 1t��\eK����ѱ�)9�U&�M�6�*��uϗʥ�'m݁?����t��G�>�B�UФG���q[.��N��x��c�J�jӸ���Lz�]������u�x���5X�g!׶��k`���:��#�G����\:���u��q{���j�>Ӆ�^�W���t,���U��2*^���-���8�R�V�Ӑ�Y��EόP21�J��Y�u��떅qҖM���s��#;d�̨U\�urj��oĕW^���ާ:]�<�b:��x|^]�s����f�R��;�/-f2�Q�2���
&�T~�� �o}�[hk��=yE!��w<�K@	�MC���6=�&��rvj��A3o�&� u�O�i���\�����P�2
Av�{��^��M�N�1"�`c�<�}��]�Y�%
x@���`����<R2>%Dcq��+������X�I���f3k�蜜7+|���\eva
��=<�
��� �W�����$G�y$҄\z�X�w�]�TjJ�+/�zPv ��ڽ�����.�����3�[��Ͳ�U�1�ԌfQ �HXKz�;�A&ye{M�k�k�����u!r3ŝI��0�c���^�y�w+ַC;[���іg�/5Yrb{u�z�K�[�5^	z���OiLs�u��bZ��S�Eid酋��?�Óxz�Q�aRFgx���˳�!�Ԅ����J0/ @^��s_��
�֖A$e=���{M"���h� n�������jY�ѩ��Û����\��翡!���A�r���n�5���u�~�G���ڭ�y?��oP(��{i�* d��� �l� �>�<Nm��1w��
n�*+�ե�%��cT����+dS8�]�����Oba~M�禴��d�A���[A8C"��ɱ�Nd��*O!�܁�7�@S�6&ʈ��4����S"�z�ɼ���Tz~�Eʓ2W�Vo��m����E�R�x�]��yf���rj�My������Uȵzҹ"ף[��������mD]�8�+��p��^:V����k��]��Y�����]�jn���|�����Z�Z���
�J}�P��)�1h�D�g՗�9��yP���/��[�R�¡u�AK�\����~��+S��47��a�WLv&�@o�����8�Y�D��BRӝw�U���Obl|Z�$v>�.��>Y,�
�I��
SS���e�"�r�2���T�N+~r|T�aA�ϋUHƳ���=�쒋�w�crEq�h,�ʚ�

��mI�=n��)��=�_둯�F^�s�r1��1��z�/��MmNK���X^,ײ��f�zE1��]b����}��3LЅd����A�~뼷Q�$qY��Tk�� !B�0�A�r�==}Z+��8'֑�hyA�b�FEƵ�mP�0�"�i�"��<����J���5������1�Lk�AKs�6��D�E@���y,�d�*��y+r�i#�Z�V����a��dBK�ܰ��&�)i�i��l'������_m����ZV� .�_�z-#?V��h@C�"s��o�cAR�kd ���3�p�f���{�L�D�d����s9-���o��h�~����S�pm����w���|OD��~H,�P��3�&E��C���M�68��b�<E�A�d��!�+�{�-pxBE���z8<�6��c�JJE�D�.�-Pix�9��f��s)K ��+I�I��V ��j㯪�w��G��Ɓn�wSh���9�[.�bgJ�\���w�q��m ��,��8�	 EV�����h�5lij�q �Eh��em�1&����P&ۦi�E3��}ʞ貓�-C�̤d��̈��C���4�57��'o�+�s[Y+o�������Q������t�����ޜ��ǧ�1N��v^W_x��4Ii��.�����8���l�5�U�j�W�,v'��R���u9@p�ײ�B�)�J"���D�t�fe��P7-P�/������z�L�tV/���br�L�LZ��(F
 
�d"�����8�����Oj���c���$:d,���(�����-��w�s?��v6���uN��=-�hԸ�[D��4�0/J����-*���9�'�	L�kk����8�ۅ���e�.��~N�$��<���f�[B�V*j&�9�é��˜ni'I��S�(���c�D>�<�yQ��t	�|��/��G���>�Y�y�z�q,$ @��M�6��m۶afa�� �)}�=}�r�uH��ܿ�idi3�O�O��U9Ⴢ���1-�	���x��GC2�]��6%VK4ޡ��XA�'�d�R �<����)�Jښ��Kƾ�qR�ӓ��V�J�T"�WRK�_H;Iql;�;5#��ȹS���/�r��|؄Gj��a����"�����w�g�}���$��^?��/�\����ќ�Ɩ��x�%�"Vr�'T�.��̑W� 1Y��-Q��ńڄ(4�<;����Ų$CcR^cv���"i�<���AL�˹U�kY��\��Ɋ�EQ�\�Yn��b=� ����<���ч��)�Ԛ[�赒ʖMNL�4�Ld�r^vA4���jQ k�	��ENÂ;o@�·���[�iB�<?�=�9�3e���/��\zM��26�X��_{'T�q�����)���ȉ��ϋ"�f����ًc�3Y�\p���#)k6/����)Y�~�vp��L�A��M)+BJ���Q���.�᫯L:`N��3F����j�],,���\ݲ��e���u�f��wUҝa�)��ZJ�2[�+mg�ը[��V���k���,�Վ�����c9h{���m����-j�VRQ֎c-�%���/8ѧ�gխ��ҡ�)���k/�q&|�@���nO-ɩ���Z�n�^\���m8�c�v>�[K��^=tp�7m�ig��J�V�`�F����[�kÏc#�����O�* �S��$#��e��K��٭��J�����V;]��3z�d�ڽ�	����nA��},Ԅ8���1���&�~�U�̨�+�Ix�|���ͯMG`⹌A��!;�E2�P�wE�S���ZG�>���齇eqq�g��6�G��cw?&�z&�������kӘx�T�m�1y���d5���g��� ����j]Q��=���kLΉ�%@(��1�N(y���ϣa*�K(���u���M��Sf�H8���1��0{?��j���W�%/?��̤�:��6.X��ʚ.S�Ϭ��Z-.�2�X�b�y�ֺ!��i�G������+矂�5�Ӓ,:�Bw�k��D=���&YS�_3�ð�>w|m,�*�"**;y��2_����W��Yy�Mj���̙��~�����1)�?mV�5�0!Y'�bN�R�C#�bQ���N	��#r�քH0i5&��������&D|�J�Z*��1Ѝ�q�x�[ f.���f������+=�V9��D2cDTY3M���{L�HQ����٥�
�.VД�P֦v8����y�&���Caq.���턃�6O޺��7���7�3��F�zTdO�ֿ��/w#�&�;EQ sP9�xV ��a>eJd�I>.�>�Cf��KE��5\��Y.����
�wP��
ْ�M���įo��5�ك��3��)Y��帏5�_��P���w�Rn�b]ý�v�\eiqۘ�4,���,��$��l�s�Ɂ�r�.k��}���$e���j2��X�3��1W#3H���������I����4[4V>	TX���;���1!���0I�0rtT㜹BA{TsRi�5�������Ԇ(l����uutt��c��z/,maÆ.��y_S���Z�ꛝ_ӣ������xf��4���w��L�T*���>�mw(E�8J��L��bw7*�M�6i��2W��Q�dw����U����6Hp����vzȓ�ɉ�s-ۅ�!�C݋2v-�ļTl�1/����
2��~�*�{0r�M�z<
5"��G��˔=��jkk�BG[���w�ڭ A�j	���Z���U�h�����Τ��W$,kZݴfrȈ5���C@�
r�]�X��EoW�zk"2>��cS�J*�09#s��s�<U�
��F1!������>�4��)����<26L��v�\� ��������z� �K��H�2
N=�n��l֣�n�Կ2ٰ��2,sv,+m�Y������}<�����܆%]�*k���ɾ�����;�.%��o�E0 �bxߵv�j;D���֞�U#���Ɠ��ﳩ,BL�,�pg(�����=̬f��e<FS-kei'=E9����������\$�[I��_�DQ���3I��`�^v#=�ښ��k���9]"󥜲&2���e����R�y>��+��1s����e�m�V(��h�Gs�yP���94�����_�}�Z���]���O��[S�b��[;�}L��%�:m�)����K#��,��(שּׁݼ��R))��eb�Eۃgٜ���UJ�k{?Y�@� ֤s)0'�^5�Gh�b�_�T;��?�,7:�?�}߾p:���8�)Oى��X�e�J�d��<��[f1;9"d%�
��ߟ�F��x������~b[a5%�|f\U�\����6JɗV��ε��"��`�Ήl=v�4R/j�ȸ�(}�$E)��dY$�V<ˌ�ɢF�YT�xƲ�<�`�n/.�h4��cl�0���^Y��Vu��؈4��j&f����܄�&n���� �������Qk���v*<*t'�M�Ck<���7���X%�o_���3���TV��&6��cMX��R���|i�;��|V|�cE�+�������sȈ�@W����>D�mxx�.��?\�����Zb��u�L�a�V�軺��a]�X�q�ElO{3��,���?Ѓ��	�;�����P�M,pK�A.�Me
�,ܧ�H[�S�<���|�O��{��n�:U���M.*%oW� ںz-Ⱨv���y��hkmB��u
�&&��yE�-�.ڨ&8:y,���R�HA+���Lm�Y��Qo�Y�_=��R��y5	r&��rrLL��FS��(�F����z��jy��v�׹�-���HH�(}�����t<��W��ֿ�1�i����c�t����P1��N9��nu�}�ZˍAm,���Қ8�
K�y_X%SNe�Ϥ@�:��F(ъyn:���L1\�b7!qiwĪ���#������UCŎ���{��x����*���;�q�4�ܢ�I����n�2N:i+6�
 .,(,Argk� dQh>�^�xn�uHE���'�|���|����}�1�*i#"o0�A�~aF�
�[�b\�T��_�	�$�j�H՞���E�����ܹ�\����'�ff2у���[�Wz\n3�n;��A���t���L0n�^���XEy.���_?ÛXK��{�R��\&���8�s�5����x������ޅjM��Z�[����X,���ue[��$(���Z�
��J+>���k�=juRq�Z���#�t�ue�mP��k�C^ÉNŜ� !VxWG'H�$�� 
����%c+�X8�	Zt�{�m��y�A�,�a��\�+*\�'�\v(rQ������R&�
�`�����w.�Z��)T�+��{S��ј�&��4�G]�^�F��Ȅ7�A݃��Zڴm��^�-�O������X�>U���s�����7��\�\92�n���҄Q�ݭb	�/ �8��]t��abbϽ�9x��/�`���Ǵ�CR�3�����D��)Rҋ��S�S؍��N84����DGO/��ǰn`����7�Z^��ߣ�G����թu셼 �`D-�rm^7��Z��x��4?r��9f����������w����;4d�)H[>�+N��5|�:9b֚��V:������^J�=�#�Tז�t<��+�����+l��ֶ��m�l-�I��R\�V��T�G�7�P۠�Z&9��BGA_C����hoU����w�
����-�	��bNV��<�j�;<n}���V1T���Y�&�Z�@�N��*�rD,�*h�&��A�ZA�*�j0�|;:p�T�R��E�\L�a��bb��0%k��Q��z\dc�<�i&$�L��kU�/�p�W�%C���P����M��A1��-������.;�~܎���mEYeMY��#����ה��ϼ���>�Ɨşh����J�K���v=f�V��J��4��?�o�2�5ia�b:Ѷ�����3��xװ�Rv�珹�����S*�䝚ifSq�� K��PKc쌯�ꬥDe:�.eķ�v��&E,��딺W�Ū�&˘R76�iɉ7�|�.cȊr��R��D�4M���E�Ǣ���;�/�Q㯭b�ӍK����_�b������ܶ炛���Z�87��~���sؼ~@�3��U=��*�,xA=�L����[�g
��d�&��-����On��>�w?�o�C��f��d�Ett���c=�����9&�1=1�������ލk>����t�G񊗿��?���x�[��g>�U9��3�"�|h�@K��p�닊��m��/�y_/��vd�	��#h�mb&o���05�_�q�e���۱���x\�y;�؁�/�L��ޏ��8±0�,��M���Y)�S�l�KtΖ�P�������W�Td`�]�9,r���sS0�2@�j�Q����N̪Ը������C#0wTJթ>Y���R����\��{w2^�W�>��pe����Zy��Z�l�Y�� �m�W�31����i�;ƕ�����0Qi�j|�ڐ�ᗧ�0����J��7J�sչ"�YŖ=�H_F^e�!���>C��8: -F�	�Jv���ĥV~�I��B�p��8JC���z+���z��ů��W�#�į~z 睵���c����5����yM�+��Ȕ-�ϣg`#���h�E�G��,���S�m�+��W69Ta�n��q�T،G��U�/�3B�߫a
FR�>_S*�;��[�v��ձK/��s����ܻ����_��WOM�����Tŀd6g)ի����2%�7`\O.���mP썖��n�e'\�d��}��~��ھ'�������f'�ZV;���,nY vԥD����J��o�X�Z���0��1A�j/Ms����8.'+ǂ���86s�L:Z)�OY��&&kN]LdW�x-d�ͩD���%�X{WW�(����ڬ	Rl��L,�T�
�	�w�f�Y�	�97���sOw�LO֌$F�<��E����&[�	lN�ew�x��^�`X�`��YB�QI#M���9���9篷��;�ܞ������ÅQ�N������z�.�t��H���R�&''�{UG_�G�Hk�S�45�%˛z�kְì$B���~�=�T�׵���Z�=(�c��dM\G�i�M`����!�<�"t "��O��3YO��?�'�|�9��<��MG�8A/�����C��T�����`�#�?��_��~�]���)G	��'���t�7����}��@ǎ�@�P�����J�4q�8sM�^�QvTI�Ϝ!�G�����NЩ�Z�q/���<Ha#����h���hr6����d�����R"��_w�r�u4:V�;��:��J�eZ����Z��R� T~��.����K�P��k���:��CVZ���n�3���*jZ7-�g���0��SZ��|X��|�+Eߤ��]�;���ݦ�	�7^"Du*�a���23��i����M� (r�hW���"sc�"�t��U@��Gji�.��ID.J�]qā��-��=���`��S5h9_���5eu�P`(���Z":m���vF�HX,s�]��L���2����-�eb���n�������)�a:�YI������j#/��ϊI�>��������5Hi��<��Mf�@2�]�Z[��i�k��WBh�%w�_�b���gE�Ό��~����4?�(�o<�p������ᱹw���:i�AI�8tk5�`�������OsrA㺚��l�cx�j����67�j��Y���AV���bY����__�Um�[���l�!|���Ȝ	"=�BSB`A{�dZ,��fiĞg�6�zݓ�5OP�R����u���{U$@Z1��ƌ��Tu!�U�tL� oK�����ܺK�JER��d�]^$R���t�����Z�:t�?�.���� IS���J�R��{������8W�ڑ��� R�`�K�.�����2�|� �C���r^M��zɺ�1�ON�R�&�Ȅ���=��c�̎�[��7��+/�D��z���;�>�aZ��C#�*t�7���o�"N*�g0�|H�A��-ѹJgN���Q�%�W=Ai��ǩ#�>�\�H	Q���~��w����F7��T+/I{���(����r��-S���~���Qg7Q{w���u1�s���r�fGzh�1�j��Bv!�g�{H���k�@U5�D� ��-{�}�t���ʡֿ�ܻ?���S�k�����JZ�Ś����t6���
o�>���z��[~�]��q��{x*�m�\��di�Gj(�>^K1"TF �K�5�	�3-#9M��0�7^�T����@������u%lUs�MB֍���Y	5G��m�/6��}��S�R!|J:�����sbZ��,(>�\~���d']���Қ��fܞ�o��vl?�{��²>=J7n���0}��}��O��m���8u�YOs����œm"c���#�NuE]�d���F�;�V�\t���әT�[�^\��������꨿�ٮ|n�|�}���o��_~���R��?x���=r�Sc��\���E�@$� !�FvX��*W�M��ڐ��:�V�&�8Wt|��j�֠Rܪ,W;D+�v����|5̡�]�J���y?�Z7'���"��Q���U$6D����h��T.z�	��:G�J�e����H���a&ua��AAD���w�������R�E��
�a\�+"F;��!�S�^u�"8r��1v}t��(��N�sh�ɩ���OOS ��\-�m}uެ�&���C��O}��"�Ǒ������Y-_A�Cď��a1�Y���ߍ���7̅�(�a����!K���¼ҕg�w��z���3B�S��VZ;�tŒ�p�<��J�E)���g����˴n}���C|�~:q�(�+�@�_t9��/^L��g� y��I�$!#�DN�ؐ��&�)?|r������m�'�p�ex� �H���e����m�ɑST/.S*���>:|��ߤZ�p�N������{�tg��r�O�i���Z�#t��{�_�#����V��x������'Dg��ϱ�V�9l�-s}����Y�j�I�s��?�n�x_ӵ�Z����l!&�m�����{������Cl�k�7�2�"p�1�DU�v�&e�!1��&@Xq1�k#e.tʠm���~C]�W]4`��%_�T�K%�����U�Z���fxz�$H~��3�7�r���R�CW��Q�E�8�`���������'�������5}�?�$��Ko�w��m��C���o��;v�E��nx�[hdf���_�,�k�m�ǎY��{��������J?8G���Y�>���Xʀ�{�m�]�҉�k� �7����������a+�~��~�_���4����u=��c������,�+��d���0� �����p���"ZhGe�q�f��q:V3d^�_�U��Q�����H>�Ui3���T�Y�z�L)�%M��$s��k���wݺ��úw���j�ڠ뉓�����IS�g8�;,+��Z%j��B�PMK��� RM��*J�pĝh�G~7�����������]r�N�5���s���̜D��XZ�H�u�_-m29���0]w�����E������#��K�^,Wk�rG:��2�مpL��qLx�1�7��uk�mT�}�Ǵg��������J��[r��?[յУ�,���0��pÁR �h�ۆQ�Պ�ݢ66�`��c%��0mڰ�~���Q8����ez�ٽ���J��x�k���8��� �H���O�����/?�{t����������n�M[�
1��+vу��!m��@g��|F����|�V��ؠeSQr�yo�~����&6H�����&�{j�hM�[l�.����:� b�k��ٙ��=��ߋ��/�}��<Lł*e��|!������J��!c�Z�ի�q�,�-��g=[�J��#N�T�7��se���g�L+R�����z���8�@�	m��[��6�/�����yy��������m:t�"��u�;WGضV u#�s��� K��_E�bƸ��sF^@F5�K�&k;9�;u=�P�P@m�v�S�2�� ٫��#�(� �F�ag������M����z�$�x(����g���t�W3����<}�Ѻ�������޿�|��ش0X�##SbSE6`�E��Cm��#��l(ʏV�� ��MB]��#�"�6n�t����8p�[�]��阥�(��x$���ۿv�C����w���_y�MW��Жݣ�����|��{v?5���b��z��.��49�c�*1-K�^	[^�1��IBw=�����f
��֔!�47��ҚZ>;J]!�ڠ����,��h4kd�+���$��N��v�
�����<=J�5���PZ�Q����p(@R4��R�JҌh�d��ia6�T���s[��y�E��aJ6P�KOj��V�dj[��I݆�� ��/ _�5\����f�cV���:����N��0Em�������t��@K3	v��4�H@��ht_m�0D9�|9�f�wQ��%Ǳe� ue����O��ߤhB��A�7m"B�9j���U�R��T����j|!�N�E���7��#�i��<o����d8(�U���A�!�Q-�gY�,鍟�[���������lٴ�������9�ce���������_}uv����O>+�i8�*%Z��b��>CGG�f����������F���:ƪ���%+�������g�������׿qs߷8�Η8��a���A�b~��{��JFitn�2}�:t��g(��p��k$
�����`�v���MGN��Ov��s��9)�����ݝ�8
*�w|J��X.�a #���I�[�Q6�=̪��t�P@t�tdH��2[�]�I��:X�
�N���%><���o���:V�mvA�JYAO;Z��o7���ƭE5�d2"~pc �⺴@��H~~N�a���@�Μk��pv��i������������{�����$*�mD���v� �����D"�_�����1�HTڽں۩��g�[�D����Z�*poW)E�_>W�6蠇�{��f&������/�E<~�,=��n�����{������k�����6����8=?O/�?@_�����S�]��'/�!'�b�r��!U��
���/`���X*)U��g�=�ke/�O)p Oh�vUx��˶�$k�]�R�j�#B�%6%���*N}c���|������߽����ï�|�L_Oi���τ��Zhf�L���L��/{hxt�ƅ|����s^݋%0� u��W� �`�kX��d��Ȼ�JV�����%��"���z��ٵc����<V�SW�V[63�jE���h7���ǹR�&�%�����5���{���Zh�:��i������z�J�Eu{��Bт�}T���fې%�'x���� ��+Eq�XLP�*����%���ab���1����"��D�4���gBf�9b��(�AZ�8����uȍB/=Qd?�$]��������)�����l-р�"@?���@�('4��7I%��1�ch�KЉ��Ї>Ď'��C�����i��C[brn����3:���+��a�P�OI�i�\S��D�|�n�Dc��M����O�����}���/���مy�0{f���R"������m�E��~��e�]M��;�Ž/ЎW�G��������Ct�-o����6z쩽�^�ə�s�Π'�A��c������Щq����s0M�܂� �"��xܧH#_+�ݿ�&�
�!�F�^:x�ΞAܚ���yTK�Gׄ�`�|�{$�!K$����=�6)6*c ޸�P7{Lp��j��[�u+��e��ce���[���fHiBv
���������L�b�(�d����ym;|�f+�a�K<m�ߜ�PW ��g1Q �J�e��#�@��D����ڞRps���9.|��������^qh1�(�2�~�ȲU ^SW5i�s2Y�@��[k���8i�Rz4�j�����>FV#O���k�ګ��O��	�����>����#gh��}��;y���U{-)��㐦!2�B�1)�#> c�Q��M��Pwo�h���9 ЂX�=��+�{ȵDR�H3(�K�ֲ�M��[	���G��ٙ�K��{�M�O�N�Bn>��c��Rȶ��J��Rs�k������U���+�o]���*`͑��� ��:��	�']�Z]�f����.��Fk��Z�xo����m�­��-�zZ��mM�k�k�T�8IS��L�g@�]��G���� 5i�D�H��Uz����ԓ�� �BY4ܔ���������O��*@I3�ͦ�l�#��D(qd2�D	`��ف�f��i��{�$9%���	�D0�svn�&gi�ŗ���+!��:A��,����8�b#G仴()�%:yj�6o��-.2�(͠II���;:�Ƞ���bD�:21F�[�ny�M����pt~BƇ�[��je%኶��E�!�����.n�D��W�$jG�g\l�r�$R�p��s ����%m�����o߾]�4�<F��4�8�竴������5Kг��R-L�st��!���~����
�`���ջ���e���B���W�＝b�n�M�X�?>�%��Rq��o�L����A��=v�l4��gi��Aϐ`�(��X+(=v��8Jǎ��(G��pbKwQ�	���,��	Q�����.C��6���A����G�D����"1� # #��:�������u������] ֹA|�C����Y�ڣ�~Ʊ����f6�Q�������,]G0��G��h�
D�jrn�t�I�O;j�ylr�~*_��m�N�����_�H�*��v%Ŏ�
W�=t��@��|6�c�TZwITVd\T�t�F�����юQF�J:۔To���t��o�D]Iz��W�k�o$������O����W������˿�t�ko����#�������\��
�gՊI��V�;OX��DT��/ؠH;���Z���-D_��m�߁L,"LS��SR��݇� �l5H+lE���̶����Sw9 Ȧ�=�T�Q��X�8n��<'��OG\�� �j5�fJ���w,���$6[��{�P�\���4�c&��a23u5�~��t�+RA�ս����D�+7�o�������*�*_�X�YL�Q�)p���<X;�10=�p�oF�+ltMD�k&��O�����0�R�Z)2i���{�LOdI�V���A�w�H��jRQ�i֙q�	�Q�s��O]}�ƫU��q������𰤒�9�Ä�r�Q=&����ť�;���UW]%����1�񵯧CGG �$"��tA:a��@��1��z�M�B���F���������~�ﾝ���Sai��OU���rĸ��ln<�7T�ܲ�to8d%��~�JEE�(S��(_�A�:�
K����	;������>ڸ�~b7���,;F[��:�����Ԕ�$����E敟��k������cg�%Y<�9ʇ��h�3���E�q����񓔯X2Z�Fqz��):p�8s����w��PO��uX#AF �>�L6�ն���T�H1�@��^Z��)�%0���Yz�To,@�=�D'��I�.I7 ���	ْ�7�� ���ΙL�ٳ+�������-:){�����膬��w�	�W~��������|?{njҺ��� ��D4��W�5��fV/�>���L���������M�n����+7?��������A����VnI;�Ț��J�Fɥ^.K��>d�|Q�|]Z���]٫~9F_?M�HE��vv��-/Ӎ7�H���M���,-��|���G{��(����Iޗ���ki���hi�J71x^(4���'��Z���Jl۠'�H`�ĸm���P��-�&���A�Ŷi��]]�mK�FMׄ���фd� �#!ղ�z;��dTq��b�T��e�<�e�_ר5"�h2��Zkk�ڍ2�W&BY�hE�s��Cf�3\#[g?�oî��
7��x(2U]����[nZ�o�\����M}%��оM�9�))-�h���֋��Wi�&�_PV��4��S}���-���}0��D����6V*���r�E��o>ڦ��kZ�]�Ul�/[�����ҟ�{��B*�D�x�Z�؈��r��ύ5[�t�9H�&9J�bǠ�=lܰYf}�����:y�ES�m�F�ze�x]E�gF������-�.��?����h�c��}�>�nk�Լ)�@ Ƭ��3�t�>��O���IJ1���?M���$� ��m>fOG�c��(�|!�>�	��{�Ej�z��N�p�g�[�I9u|�>��O�����P�y�
#��C�K�#I���a�U���LMQ��ˀ+��.����^ą��Bmu\Ѿ�8!�_��l�v�:��b���uq$�,)=��q�H�����r��_F{��N
��Y��ə<���l��d3���C0���G���2�K<�?����5x���JbA腴�aO`7��U�������9S��M���W���o�i�k~��aƄ��j"�����8z�� �ke��8x?�]��ט ��Na� ����
۴�Ճݒ����`"�w?Ut�n�W�y�̔�����:��Ku�h7�>��ߤ�Nw795O��G	 � �JK"d��c�f0�p.��q���X�����vWf>T���="��2{���_~3�]/ܯ���~�0mذ��Q)�˳�Nɺ��Gts#d�ɤy�C�*Ց���ѿG-��}<�?'3a�W+EY��;�}y�(}�zVx�Z!�P���&�܏����0G�giYIQ��Y��!����# ���jɍ�k8~� ���-s��U3�-���ڳ��!ʒ�\X����?���h������^� �_Y?�n���7�c����7���ͥ�θ�j�h�5�D��sZwy󳛈�8Y؎I��*�����W\�ZĴA��f2��T�u�J(Q��O��͎K�s��!q�!q
�Ă��!�ʄ�ʳk"p��iLD�t��ӝ
�^�x𚅅����<�c��{�%��Dn�X�+���_u��p��,�����<~r�:*�49=G�B]�^1�	=u�� ��S�xLq�N���$[Zҋ�0?-�"���?��N�mj�y7t�sj�
ԧ�}0�S)���q~f�ju�=�p���=z\+3�L�D,N#ã�������������u����	Gh.��N"��[+�`�Hc�Yq��	�(��R\y�|���8@&G&���p�0��TB`}�|�0괭�_&��P~M�f��F,cD�T��.�������}��s���(P�(�LI���!�Q��ɒ���ATkE��*��	�?H��:'����E���f7Ip_� �0����Σ�xE���"�s�}e����Fr�+#�����y��^ﮰ+���)w�h9�Xlլd�y+�]K��?�Vgn����U�DGpA�m��Yk��$b;mKϐ��_��v��j`�Q�bx���������IM��=d��M/MV��o�x+�
9Î;��9uf�*�i�q=G��`3G�5����� w�����׾���Z��O>Gw��r�ͰM�},M/�͌�9��#Z��A��g��^K�^z)��k�����+K�9J�w
O ���>����*�j!ҁ՟`ۆ�2���&p �T�M�����Q	X҉�؉��^��"�P4?B������3��|�b2�O��SM���,�� [�/`��E��e1�����E��bDP<�0��V�s[�e�P괻/|������c
�N�%�|�ѫ$��O�3�Zʱ�'�y��$�<6^fY�j �bA�XMY��I|���,��K�S��!"��9�vf������s�0 Ą��`"v�b9zs���cT�E��^G��!�.�Kr��q�<�*�51��!O3�Q	��H;��+|�1��X��F�Ȧ�y��eA�p|���&�dGT��8�B��s�#}��'��lG�h�c�a�!��Xv����	�p���%Pt�Qn���v^���ۼ�����)�4/mf�iA�L���kF�^TJjZ&T8 �h�e#�ѐ^�L�c0����Bmis\��2���]��K����S[W=��#�/��i;m۶��H��!����!�M�5"i����q�, �ax������H6F�AX�1P������W�|@���@�}aa�K�N��ܮ ���ubSq)���r�9��ɱ�v�:ٵ�"O�?|�r�1��uJ���dLF�b�*��F�̑H���=�oS�ݒn���oA��GZ��Ag*�P��F�gy����8�Z�iV�׬w�N.o�|�?ͨ�d�����P:Y��W+U���[��8t�9b�����$�O�eYOHi��B�A�X��BQ5�ur�a�F����
R�oaiY@�SsTǎ�
6��1J��U�
�{nI�[3��hԁ�f�_[{����S�����ӧ��.��>�~���/�d�&Ɔi��f��{���/R�*Ty�Gy'Rl�R��CԸ����C�|Ow'�띷ѫ^��so�o��m*3��֕Z=�gq�$ӊV\�!�q!�S���H�$S�^EĲb��*U���uc�>3�,da\�ץK]D�tJ���b�0�AN�BYN�!u�hnJg2�N�'6(ō��|��٩t�ʵj��U$�<ӉS��0���z���!Jۆ���R=Ix��%��ns�"��j4�C�������c=��޷":�4��s��Dgh�H�.tֆW��F�\4��4�P)�MOO�5�\#(lj�Ƽc��
�,�%�;����	��D�$iiG�6lG�Qc�j�S��@z�D�u��������Ը�&����6����0!j�b̤3ғ	��U�a��4�KyIS���b�)�0w����;�nZ�q�� �����a �f\��6��E��LZKkzӕ!I��m�r���}�kD���RP�ý�C�s�JMXG���8�x@�	��x�2���$��w;�ꆩTD��ЋƱ�V����t�����.�?�����ٯ-?F��,G�)�f��i�htj�Q|V���I�38��aF�PZ������đ�'�J��e�=y�K%�zψ�O�B��;t�^�M�CQuX,���LN�Z�^����5dP��P#�k\�ҲV�0�8&ÁO�1�96��s�SG�ZG�X]�*N���=܃f��V��;�opR5ݥB+��Z²V��[���y����Wg1~��Q������ͮp����ɲ�(�Y��,�R���G��:]�_+����r|��
���<j�\g��HOúA�0̀{E&��S�w�Ly��R8t�����<rP��.�C �D:mxOb�+:'P�Q��?�U�)m���i=j<�M��N���|�X��`���L"-Ƿk�մ�#&���|!���	%���1��-�`���y/S�2�IDp�8��6d�"�ј؜<�5��4�����7\L{_���|�����b�5;J�\���2u�tK�k�R�@��<�"��s�i� ��M��n��_x�Yz�ч�7��D�}� C��nPJ�|m�l��a�����G�G?J�r�}BU�{Xe�1��7D��0�ѣ|�v�޽;�c����ӧ휑i7���� @^@p�q�R��_��9r�0����U��R���L���k�Qc�Wы�K	�YH�ScA��W�<�|�~���`�[�=��0��!�=6Rè���jj��8�������0��P����PO��p��1�����޲�F�:��2m�_���I!=�� �g͉�1 ��c�˘6����l�,\�T�  ��IDATET�Z�ː��'h``�6m�&����G��]�!��D�=��b���q\��0���y�B���P���(�͢�$��XC�Q�S���j�#OhKm����n\�� ��.�>/�<$������5�����g�t��jV6���R[���d����7i|�� @��6=�]$f�@u$8?��P_0�{��+���s����!�����5�,�����^A;;d��FK���$=��3TsCMey=g�w^�V��Bw���-��0'�Mx|�I6h�h�<��V#�l3�Cdb��g"eǏM�9�0���q���8ow�V�-���K���T�D�l`����*y�4��i�ګy�ڤ�HuJ��`���/ ��^Y@�V�5a�AER��u�<<�
pZR��չ&!���׀��W�j�ЁѲ2f���NT��>��T=6V���q��җ<O��{��J��H�DTP�O�wU���s��W����qr����n!����@-�'����r�ڡ� ;���a{q��d��*&8ԝ��[)�ض�K�&�� nq��d��k�����+�R&�����#S�����Q��c~n�~������Q��F����F�s��a�S�s"��v�Ư���O�]w� =��~*�h��:Z,W)˶k~~Q4�!��ݞ��ǎ��[n����KlGJ��*�l���mt0a&:�,�U�-�ˀ;U(�=����mX�z�Χg��.�������}+=�؋����.�p����������7�%�n��/�іmk��g���az�m�H��i�_����0�lI�; ^��;�TJ>��	����
%���8�H�����#K�ƈ�.	&g����@[l�<IӄBVȰ!���6���Y)$�7�Ϩ&Xi ��I��&�dg�Rm|,�퉃oH��B���U4�:GG����B*<OJt2�n����ˋl�i���I͈�?j3�8�)�D��mٴJ^zy]��Իf@괩dF"K8C�\C����&��7>�͔q���&B�H������.�����Iv0o{����v�Lr��A�����_@�T��v�-�қ�P��@�lp�!��Mؑ��k6Z00�;��8?6�xH�h�r�Yy���%-#�a����樈�	�1�J�37�R���� Q�x�f�f�z��o��9s��~�	�9uk��Y
,�cnqd���Ñl��g&yU�t��A�֯Ӻ 3b{�zفϊ����G���1��m^��9�K}�Qu(ÿ�������ŗ�lE��R\��#B4C ����T]��箎n��]%�Mc�Ċ����rm1�%�D,"��ohP2*5�_�[�l��uk�\��Y���XX�&Dq��;(ǯ�HW��q�nD@�쟆R�*�ʪAJ�`�_��7Z
!�Vh�K�SF����T�ԕ:���Pӑ�jmO2%��6���޼2��-)k���|��]�$�[R�ιj�/�Eq��h=����U�>[ ��������z��X�'7t��w�do�y�F�ne��_o�~i���S�=z(��g�ޢt�0��"S���X�jx��~X�%��os�ppձ580CK����j�ff�i`͠NQ
2�)d���;aN)(0�?I�t���Ob��s*�m�V�a��kʔ]
{Q��S�ҋ�����Dr���ˇ������)�8� � ��-�P�锱x��y�=�t�Q���o����h�Xl$��	Jģ�c`��k9?~��n\O�7pT�:3|�������_{+�>9F���率n��>��ߢ�[7����O_����Ӄ��O����G_���g���_��+#�'��űLT!C�\ D����f�}|pp�α�3�db��۶������)���C
�P��[��*�oؘY�F]�cX&`�����C�˗�r��=��e-�⣅�!��,O�}�w�J��:�1���*����	� e<�ֆ�	G��J���@G�d�0NdDx1vV�,�~q��x��Q+Z	��8��&1Z	ʌAV@�Cg���4,�>�'B;.�HR%G������$�Lq,�/<$jo��r�(g�cT��ԞD�0bY^��]���L�e����,�}ｼX�e�O�:MW��z��]��_�S�� e�h���݈��X�$`����f!���ŀL�[��щR��葩y�*e6Ԉ0�5�ꭕ�*#�+5q�x&D'�T p�	 5%��6�ƺJ�B�ؒQ��p��s/�Ls���/C�,%�ma"\���� 4   �T:+�Q��;qL��
����a�F��|1'`�b
�|,�DRR�6 �Au���'���y=G9J�Mm�����uok�d��Ϗ�C�0hC���&�Ej�t וʅ����`qa^k1��s�����mRR�A���c���O��DL^M��#��T�J��SL[�����i����`!�(mJq2aѧf�nc���2�zġ��q�_�Pfhh�:9>�I�u��9�A	���#�S2#��t�S�V�Z�U;6�q�j�?������g�kW�ן�i-ϳ�nyo������F&-%��u
'"���(7J�MaE3� ����������\�)�e��Ƈ����������s!S� '~}5\��Y�r�$�0/�l���o�m�Y%�}����+�E2��,0�e?�{�T��_X���q8�����ZH,dH��ϛH��������C�<� &�ȅ����H�U��u����<���P�����:_�H�ҙzi�a��_+�*�@K�f�;��ZQ��De-�O�QOo�(ϲ���sϋ#E�.,U��s]��؏�� B.��T��w�4�e;�:�r�70o�v@yqi�}�a���Ɯ:��_����[o�������k���dV;;����sZ.�٦8|��h�x��0*q(���x}��U���?p���%^��H"\��'efY�@CT-�jĪ�J�g�_�`�7�[e���؟�Bbn��x8�vHX����c=V�U���pm�f�.=#	Y�!����Cܰ��j�0/�\)ϸ ���H؊G.�[(�Ѫ�v@��PlОCOC�u�/6$�4�xц��Qs�J��"Gp�$uc
��<;��]��rI���|���ГO�o����Ӊ��2z�3�DW�qh ������.�z;�:��a�2��&��zU�8Bk�{E\�W]D�Ss��g^�K��Z�k7�;���t�5׋�R�]��fq����Ȓ�*>�Z�Ħ��5��FU�H�˰>A�֒�5)��Y
���9j�°!SյP\\��n��g9�:~g��==�y-����>P_;|���[�L��Y:}�8�{�e1�u�6�|:9�]����;ʠ*O�]~8����c�9��^z�.�����k��<$���.����>>���0�mxl�v��RZ��N��=u���������xcq���Y]i��(�jƁ#��z,)NU��m(�=�yv�T��Z�$��ľ�R\���q�΅z����#����iZ9&�rf��%�d�=��m����=�����s��8�F�������n��Y��8v������-�.��%���d°N��>�4��	��g9U�@��\Lu�ܬ���kZs�n ֕ C��6/5+��s �>���9�7G��,��AGW��D�
�S1�6��=����JGTE�ڠ���܀�\���E*{��YtK���H8C��d��3��]����H�(�'�Us�K�G"�N���AEA���ͩ�i*�V����$dV���ao���:a�
���?�a���U�d0���7r}�o1^�epa8�)�
����aݕ}�t<4�_ڻ�2|��]��8��x5}���JY����cl{�5�5��d�&��n%�.�8���%N����b���S2�����LJ�g"���7@���Cꞣ��K|���,_�d�0�-��IT��Sdw?�b�t�;����_�')���;w�{���ŗ�r �@���|�����Tv��]!�O��5NaY�=�If7+��n�:F����nݟ������^��¯������O������r�zw"�!�Gтo��";Rd��~pl�5����(�E!�K^M����@|�l�����N�:%�y8F�rȁ^s���فœ���W��b��u���p��eJ&24�0���B�lM�.��̬��غY��xD1/�I����G�h|�)��[������ȶwS����=D/�}����; �0moI��ޅG�Qowg�����*D1v0P�tu�!Äd�`~#1(Lk�Հ�%��m<��ؘQa�V$���W-qBX�HӴ�NAWw���QXB�V{6�N�@�O���S'Dyn��e��w�Mk7Е��H����B�v��Jʗz��'�ï}-�/ѳ{2Jβ���%�$h�n�u;�~:r�(�������ٟ������������e;:��{���ɰSG֢��W��[u����eץ�1*ߛ�<!��B}=��NA��VH?FݰN�|��T�ny���ӑ��W�ߏ�?x/��G?��l��޹�f�������N7���숣��ӧ'e�m���U�.���32�2�@4�	kB":��ex �`���  B��|��2-è�1JV�e1^`榑ꬔ�t��������ɗ��f���ރ�Y��H��~�15�7�jG2Y�v\)���w����Ei�^�{��?s�ZZdp����T����g5������x��z3~vem��,Q���7I��Z�f�0�M�>��A�7�0��(p�-�Nl|�#:4`�u�P"-����5k4;� u[��%$M#qŅR�E�x��֎ۍh����ы��L�s&��J�:�r���!s����������i���T^^��LB����{�V�e�g����b%; @���!G�r���G�v��s������-Oge�Gy�V�yQ�� �IpnM"u(�֪%�fQ)�!=ި�hvz����S_oT���Ķ��� ����k�����(&;ۀo~�2��Cw|�N�0��g��C~�G�ۨ����7O��H+�ۨ�r��j?	S��g����e�d�?|L�������7�-�bG]���cbU����? C��ŝ��I��(U�����..������{dS�egU��i���/����`��;���GR8h�A���ӻe�J'�00䁝�%F�!*Uyq���)���C���`2�"d��r2.�C]|��������ԓ2�$6d��5�=S��1;/�aHC#]��+ݖ��$�l���s�����^�/�ڛ��&�<�� ��B��S�Q��сI����LJs>$�G����v�ʈV��Ϝ�6v��'�m�Vzamf�޷�:{i��ћ�|?5ɿ�-罚�E�~��stzd�Q�J��R������I!��]��{�y9�L�&:xl��0�j!is�g e�&��͓�"@k &I&6���RKm謅j�te��(G�eBi�P�I�rD���0��E�2}��>H�_���w�#����P�K��w�Q2� B[շ��G�����^˭N�Z`P�����GX��2�>��W��y��:{ya��XP}�!��(T�"�� Rb��rM��c�6�V�͚F)�%�hq��{��������~��s��`�2�s�~�gO�qm���j̎JIKǦ֔�M~[�|�,�O����V��'T�����J3� �l�4D#cS�z6�pP.�*�Rk�}���v�;��e��9.�jq莖��;�q]1_R�ZԄ|��j�� !��.�*�
�жZ�I�d���@������)�ml3*ұRV��]W��F����k���Ll��±�4CZ95}�*Ȇ���	�95y1�J*���g�gxb��ȍ x���Ҽj&5�S$���_�U�9&��fe{W�,� R�_��_�x:#��<|�-L���萁3G0+$�����ό�i������ҹ����o���_������׿�/~��w�}�2��o��.��r��_�����+��6>��/������x�y oxQ���'�=�MF{%o�o�H��T�͡���ա�����_��e^��$����7"�Re6og^T6zѸ�s�����c'O������Q�ZXZ�h��z�{�����:ڴ�6o�]�������B�o8&)�6F|�_��=65#�N���\�ʱ	1�R�xx6�O���%���<�Nq����5k%�A���!5����m�^شh�HO����i�B'���za�><2"��'}�!(�قpM��U�Z�� �Gz�Ǽ>�N�M��%ՎI`x�0j���a�ф&2�ⲴqtSw�F��EްQ�ɳ/�s��c�4"�����:t선�;>�q�����u;��_��Dl�3�6<��َ��A�4>Y`@����Nã�5�Y����١�bp�(6�MA��tp:�f��� �O�uk�-�F'��}A�����d���J�ZʙE��7]{ݸkU*�N��[h����=wQƫS;ߠ��a^Gj���z!G(7q���b�}k/]|�N��w�g�E���O��_�����tŵ�d`�O��%3�`<��:�.aG�L���������;QS�sG�W��E���B��\zE-u�.d�Ԏ}������ZkV����-��O{��܋��>,�	¡+9fd$ %:ђ��t��Q7��]��\y1�p�մ��h�q�Rz��,Ȁ(YH�qV+R���Q��4�OW;����&ƩR��~I���6#��SO�1`���=�ֵZ����F�* )���i�'��P#��`��`�i�j�4�x����I�V���@>�*�3"V���̇��%��
pd�R���{"{A�N�U��1�>솒�n��R,����y�����q�G���6*a�;��r_,�D�-,�ʔik���J� ���;X/*��8pw����ꠋw�/1�0���K%l����O��������ߢ+��B��Ga[���1yoY��f;�G��z��w��Էv#ۻq�^�����&a޳�U.�~"JS�G�ҟ+�0۰l(�{Z��Hf�D�&$�E4F��@5�V��5� I��rI��kR�̞��F\J��x߬E����(��5��n�F��J4��0����ECI��ˮ��.�U��3����W�G7��,=��E��4�'��X*C�JQ�K��G�1��`;⽖�K�P�G�d,l���ֈ��r��Q�9 Kuf��;� ���sd{�����N��|&����Ex��7.R�!"t����Ąu�S�!���s�q�,���*��Ԏ��9�&zX+;�(2�qM��i46w�*�� �Ju��'��Y�Nav(m43w���#ߺ|V2�-%n��8��h��I�dXر���Wu�Ԡ�������~J$3� ����i�"Dd(��J~���؉G��BҎ�eafMc��"	)��lN�Og#Q���1�ܾ���9�&]��/��e�T��� ���)�t�i���^��%}Ks3t)Gw|��W�����y-G���!��8����߃B� ����NIB��t����	�C�Z5\���3�ټ�1]
�&�ۯw{~���V������LH\�2��?�ں�&m45�u���Q/[-K �2�M���^}��6��հ����y��nZK���f�Jt�5�O��^�\�������4�K��%��H8lQ�ke��6 ���[[���Ԝ�-�b�0�!����R�|�%�/S���Gٱ�bHW]!X��3���d�-Z����)a8TQ崵�(�>W+g��s�K!A���H�F��9��C
[�S6�Wm�l�ع�B���495͑(lCT��2g��F��'c]!�B����A��6���X��\ԝѢ�=K5K�u�8t��	��@X�M����	����[�ԺKmI��n��]��m��7�DC�T��dк����S��LC��=�m�#�����[��vi�NW�5t�k�.	v�z;�؉Q����8@k��?����03M#S�!Pe�8U�
ۺ�e[T���r�P�U*���������4(��x�Xc�N�ŬV@K	�X��RX���p�F���U�JiO<����%��P���6m?O�L�=����0�D�^:x�Fx1A��k`=�.�I�ꨑ{W)��p�h�a`j�B��h]�9�V�Le���j����υ�%ڨȋibD	���S2�R��A@�@��jie�~7o�A��H7\u1��u����C�^���n�?����vHo3���Tz����d�Vr�|j|M������U.���a�`�;�z嵒�t���Y�FH�I����\�zSg���:��6r�kT,y����4���!Z`Gecc����$�/�<%>�:f-�s��J�"1Q�6560��*���s;��"S�q�=�^9�~8j�w c���鋖�ֿd`�Ne���Py�כtn];uҩ^�E̳1�["I�nݾ����z�)F�|�.��E�p�q\�tj|�7�2�O����Y��Y���U&`#2�v��'^�h�����E��h�wHZ_(fG�ZD��	^���n�F%O��G�}x]�Nz��c��t'�g:�ԡ���k/�`�(�)] �
���%�=�N�e����	����g3�a��\ �o�����g۪ �,J]�����z��q��|p�5�8�E�����L�����&���0�a,(m�hu�|X��)��eLD��}i\3��S�jR겖,�؛Y������D!V�rM�r�겁V�
�`�� �"-���=Gi���r���ȴc:_�Sp��.G*P�~��/|��tA��ӃZ�Lis�&y�!V���w��i������]��Uz�[o�Sg��o}�9I�S3��`ъ����! s-��K_8�4ʪ��.�${o�8;�9�|���0t���Kjܲ]��ʰ����M2�YP�Z��3�cP��!�if9��w����v
���r$.ba��>(�w`M��ܻ˞��$3�jZ���BH!1�k.�	V
r�L���ꥎ�5c{X,��[OU�A��%��f�y1Ȏ$�0=?_��Gn$)�c�QS�x!�J�x����t҈�nv11r{�6S�v���Kt�o�֮�ǟxX�<�����u���fN���a�����=��b����F�L�'������ZH����Wg�d��e(��5q���o�U�i>8M�G�&A-R���/-,�`�Ԡ�ك_��Te����/e h�o۱�x�ӳ{� �o#u6$q�:3�[�-�IB�U!l%Fb���D�h����(�9�Rs��+lBa����� ���%��B�7�5+Hh6�N��#�Y���9��c�vu����5g��g@$=�":��Z����Df���#%���Hq�29ɕ⥪4$ K��.6TW ��LG�b��;�Z��~��mF�k���L{w�0����������BZ���N=�|XZ�� �+V)�ktml�6\]T[�J�N{?/�J��ü6{��{��7l�W_������������ ������A�%��,�r���X'�}���кA�u�NZ\(�5�m�Ç��G~�]p�N��ϋ!�g��s��� э)��mN�/�(Ε+�"��Z��ǹ�.k�wZ�ns�z}k\S��l�v$�M VҝKJ��;-/,�Z�}h�#�Ji�Ώ��o�E�w�$�?xH�8B"�b�Zp���Ǭ@^�V#���u<<��	>��|)m�����
�1�=Φ�_��W�Q��!����>��k^Y�Q<�Gj���@*�Q6�Jp�ٳ������O�ys��V�YXd�>)bW���-�u%.&ѵ��ݪ�?�5 ANMJf1��G�l_ ����f����ʟ������-[���G�A*1(���i����D����]ߠ�G�'�b�[��	Kv6���L����L�\� 6S/O�8A�DZ��Қ�Q:f_D�)���Z���(��vqr�#���iK�s��)��,wt�ۖ#6��?WT�p8T�Fc.�0���G�>AI%BqS�F�a���J|q;��P��ٿ�;����?�;��S�r����;hbb�.��
v]t��Iz���h~xq4DL&�>M�DZ��=ө��\=��E�r������6�.���߆���yGw��!2��O�fyC����$hM����w~QZ���7Ɓ�'铟�]r٥t������u�Rq���9��1+�)�zX��������@*cX�~��f���������/jЌ>�~��b�;U�z�uÏ�dX���@�B~��n����N�@�����G)͑$�"�w4�I��R�r����cokF�����}���9ⱡ�#�ĈG��-B*��IWj�h�Ni�/@�R��0���)z����uW_N;_sJza�M."B�i�\�{��� 9�(85��n�F��h|bZ�sˋ0q�8J�Jգ�}�����+1/I��V��?h>���H3:!^����i*10����(�S8��ݓ��� -��c������Zyp��zj"%q�Fj��x�OS�7A��p����<
�ŵ8}�~+[���+����u��_D�2� C&�LK4��l���g�%��9���N�������׀�b8#� 	�u���c�}Q�r����������n���[��/l�R��+���z ��F������Jֺ�w?X�X�A����/��(��{Tuc��S����9�����em��W_B����t��5�z?��T@R` d��FJ �m����DR�rq��QF$�])�֔�]2� ז�E�a(.��M�"[��)��_������:��>j�$ �T)+���T-��b��zץ5E�%��H�%�oM����1��:t�C��T<FI�h/��x�֪���<?'}��S�d1��"����s�rA�a�E�h�*R�7]����L`0�e�RfgX-D7L�X�'����1z~�Kt�e��Si��w�#�=M��O��܂��d3���Q$���t�-�d�5���aTo`���QM�l�v�+�����Y��S�aA�q�,i �Ņe���aCU/�"m�A ����D�l�7�A ��"zuM.r��d��h���p�T��&�I��V�m��6/;�pL3�s�%��� !���CY-���U����J:�	U���*[��!�������1l�+�� ��ܢD���x-827^;q�Q!�s_Z�l1�8^�@h��Aa�
�_PG����B�p��^De^]���j�/`A�@��+`Hj�ܞZ�������mt��zy���<C3��;��H�457+�Ď?)�!�w�7O=��;t���{6m��N�-�ڍ�i���Jœ^�j]�b���u�J=�$�&�)�NO�C����i�e6N N�-���?�U�������c��aY�O��Z��L*%�#�Ǖr��&@[������W���<u��q�5׵�k��I*����=o�gVp�s-�5�^��񴲙y]���T�r4��V� 8�K�g���S���6X���zC6c��E�,����Ĵ쯬ŢD�9�D�~B�jNrT�kE�S��2��7�$0����u����0�$���1�d���dXsm�?��#�*�*���*#	�S�Ewc����$�� ���3�:D���_�e��D�I��Vq�e�rC��Ҫ�*ΐ�A/J^:A*��Ș�%��N��2�p����z�}��g�$�ݜ�W���^�+����3t�5������i��S�M���-�]>19gD�J~\)E#`\X���А�xX�P:�_潆�Q��Ed�0��_;��VͥS�STlXtޫ^E��2�1ض<�¢'�l�ϕC�CI*�	�㔄��v(3�-�Ar�j��|UE!���KӚ�n�$ک�����6�43�S/H��b�ff�Hd��Q;j�I6z%����t��ܦ�������k=~�r�)9y؁�F͔�������77�4�RN1��h�:��u�e�R�!rK
U���-�|I��+5��<;��[�Jz^�CCz�����Q���!�?1�dj������s}#���bz���Y2��	+�g@�@�b(�*��BO���i�F��إ�0t��6��H�"��#��C*2�Tw 28H}�N��j�n�d"ԝ`ď�s ��(���f}]M��uF��;��ya��P`�I�()����LGMO-���@E�Jf��&I�"�����r�(��<�z���#�Xri�Kh��!��%v���|@�C�,��Gj<.Z��0B�&�!~�|�on��\X���7_�i�>C��;�-��'�m|]�Y�24�g%�|�!;�G�k��}tM���J�䒯������OL�t�7�oh6�hi#�rM+�dA̦RY���ԥ;�Cw��k�e��4�`�Q��F#'O�^��h�L;�޵B�*V��U�1���\��gi����x�{kn��j�L���O�3�J����W�ݿ� /&�����`]_}h�[�����oE E}?�m��*�����֢"�N������]��[b �����T�K�3�v����a.ZK��h��4ۑ���j���&e�/���6�s0�r�sK�.HI�l����f�=4vb�m�ƆOQ���_w#��կ�)�k��>�s��`�P��& ��
PY�:W���5�tp�˺��$6���A&Zd~v����z����"2�q���˼A���ϕC��۩�m�IG�DuVH�Lj�5l�r�����g��Fn##(�R���1Zfg�q�v*�x���na�{%�}7m!��#*��k*�fi�	q�*%�jMa�8G���2��.�<��������J���OPqy�#xF�N�����q4���c�)�HK�g�����߸�2q�&��pԿm�>�<�[�T�ela�Ru�s�6�����J`����uwd2��#vK��#fF6����) h5<~SU|����qڴy���ɱ#;�������4������&�	��T�
��J��Y�2�[�p��=�#��'�/�������WG#�6Q~/�^I^@�	���4�[P�����l�mb�ZUB�Jo�x��u��4���1���d;^_n�&C&��3iQ�C�e�}�@V��n����.if�����(��oW&%�d���y����<���(6��ّwf�yM��}�������b���_�^��� J�o�����H�R��V�J�煉i�W:�����{�YrVע�NNݧ�t���(�F�eIc�s��ml8�m|��{1���� e$�,Q�&����t���^�:�3|������:�TU����kY�S@s"��77����x=�n �p�uL���"H�,,jV��'��ʘ��}=?��R�GD�Z`��_Ν��� 4*nP�4����n�h���3���
hfz��|'��/�����;š�*G{���V���'���`_��ҵ8��l;�����<�y2966�2�i�	a�=��5 ��u����v�"��Ҥ�,'�Lޠک���_7a���5l�kG�M*U]1���N?r��;��k�#wJS�� 5,�x��ٶUn���q��-[d|r�{PS;�����!Y�z���/�`������ZD�l��Y��[�0��PD6n\O��NVB#(���C�O���إ~']���E����
�U�˼���r��HL�m�LfL�`��4�]���k.w:�d�����q��������]}�JZZ�2>1�LT:�e��: D8P�Cf`I�/�S����g2�e��7�w��߉;$k��;������a�Gr
wF�1:�Z!.Ҵ���\6-ͺ ��_%����������:\& ��Ă�����O�!?��̼tw��d_�"N�΀���fj �@X�B�ؠ�WG#��� ��y��D��F�����ZQ�������⃬:Fd0����Ju�+�d\P�W<���!�|2���)�F�p�fJ�Q�
�#�1(����c���`�V4!�<�(��G�d�Kp�!3�c�Wc ���"%:LRYJ%Y��#�ǏI,�A����;��&q9tp�X�֚"is����,4�q�.4�,��f[ejA��ꂤ�!&T3�6dP�@i�݁���M'��X<(�6����Y YGqQ��fI67ĸ2Z�5
�̦qMB���0��:����1\���6I�?P`zb=�K��L*.�ݛ�:<��Ľ���Yr�����b�[�8��nl����{�|�ׇ�P'��7*;5 KY᮲�8h6z^�֭��b2�MI}��?#����ePt<\�(RzE�FU��qk��YV�;}�'/w��5��x1�P�9�;��;/U̽�kｖe�v�dO����(��벨�m=���E�5��&��җB�� ���:ԡ /:���%WY�k��)d?�)st6�}\PۄJ!dN�j4zm�H,t�Q�s�0N�ʙˑI{��`a>����^I��]r���B�L�T[5#/�gعs�\w�u�۟���ڵ�-��~X��_�K���V)�4;7M���n�B�԰ �"I���t}-Ȋ�~�K��MF:(�|F
�EJOװǂ�	�Z�$g\��`˭�6F>l0�2d�Xl��&�I�J�DĤ:,
(L6,DM(�uw�dAo, �Sh�j�b>ˌ$*�`b��������Kj���^��ŷ�ˤ��ʇ&01Q�e�P�Հ=s0���9�jdp��T)�PDy�(�\�y�[�(?��o��};)Q���5@0k �����ŏOLU9w���IU_czn^3�E!�r�Wǔ��&q��Y����B��u����ӄ����JQ�L�F9�G@���-��!����nP�GB6�N*7?Cֻ�:ʱ�òn�F��0������9?1.��v�A���l�����̗��#�u�H,��/��BFT�����\��TzV�F�j+��&(ъ�	�-����N�1
���,u�A}��[*��R�rN�����]o������I��Ռ�&�+&t���6sa��/�v]�j��ě5��dz6/����9y��������hs23�uTI����ٙ���Y�k�����OOʵ���<xX�>.�3j������"�c<�����,5��0�� ��W��L��:q�G<��YƆk}	���>�l{���2t�U|�2�����O�u=I�]�@D�ԡd1�D4�u������l���%��˳�R��:�x��; ����bhMq�O��/�1����G�\������!Y֞8�x%��K=�t���>w�k��3�%دz�Edk�D*a���M�62`d��K�	̒ͤ�.Wmb[��� RG뽟�}��Vg=?!v�ƔB>'�D��I�҄=��L�(���)ٻ��A0FgN6;gir� 9���fҵ?��f�5�����it)#�Cu`\O.Y8��Pz?���,�x~�Ԕ�{����������亏�&�/������ȁ#C�}���^��t�uHV�$��صϰ�f�@����ԙ���@t�1��i�g=�"V��L`�����Nج�(y3��W�ɂM��#i
��u�:�#\&����gx!K���U�İ�����kp�M��}OR�d:~W��%�8�r��b�ɖ~Џcan����Jy�5�\zFz:����mr��^i���3bi���)i�7Ig{��w���	��9!�n�@Vjf�G��c'ث	�B$E��NQ
731vB�oE�l� _��?��G��=��#���2�k�E$]ҍ67I���d��\�H�S�ߑ�1��Ms� �Z���u�-�}�w�}262�l�E�J\&����薣G����J�R#�]�P2Ց�%�oA�����HD��\�~�<��3�_Y~&(�V���ޓ�imo���V������L����t����Op� sF�Qsg�-�)�z�7���A8���۽�9��h���S?������g?�	Y��M*r�X@�n�z9#�ɪ��!&�����u�2�ay��������>}�%c� Չ�&���$��uC`���������z��s��'?u�l�`�����W�r�<���׀kq�B#���쯫A�(RQs�����1`Kg	.���u[U#R���^(�_���\�Ñ����R��k�{#m'=h�{��N�Z�>,# @�R��$g�ɶ�`VX5��ǐ���q�9�U�r*�4�/���X� 6��Hy�����y��n|>��m����A2]�s��	ͺ��QzF5eZڷ����%�'?�T��P�k������ǃ{�c�3_�.^��:.��1�
F��V�X���#�G���H��Ax'-B��@5�8 1`�k3��'��Oˮg��G4���bN��� A��������(���>0,�?��TC�(�D�#�1hFO�(�{�H&�6�J�1F5�������Ǐ�V��{��[8��E쓟?�8+�ss3l&�5�9����&4[�ģ�n�zr�@�ྃ�L����Sr�<-��~��`T�9+jT}�q���;^��q�F���x���S?[~�U��d������1jDI�%e��E����G���/n2�-,ZSN��T���`�N�XT%HL�0�(���5%[\��<��}q���c4֡0K#�� dq��n�3�
A�Ğ����#G�]���ޕ�۞�g}�eޕ])���Lg��4K����1��_��#��8�e�s,�l���IM�~S� �cllDJ�E��ҋ�����d��0J�1K.�`+7@{G'�>��=�Չ����ʞ>��:�!���\���	��G~�,JǏ�]�o�"��g�������^����l޼Q���Ԉ�9oݸB�������dl�ע����]�A�H_�n������3n�%g���m�J@d�:�={�J[P�?��޻G��<�ѯͫ����K:�R��gv3s-���,s,�e�圭[eb�?rH����˯���|���+�H��s�&�n�Hz�����d'��ϕ�|@�uNOHA���]I���Uo������<��ۨLH&4k�赘N:��p�$�^@�`���.ft ߐ�{�#J�U3ϋ.��r ��Ygm��?��b���t�-��C�������i�M˧�NГF��?ؽ��B0�q���Dc�,��:r���K��S2���TP�)q�\$Eu���V��a�����`��� �-��
"�t�SI��= 
{瘯�Q��Υ����tr�x�˩���%0���������m�~�F�$��3]q�:\�*6����A�/��n@�`�[~�@�4ʕ��� ��E���☤�c�_V=�ߵ�^lфanvT}�nI5e����}T?CP�����>&e��=�ӿF�_x�� �T;�Sg�A��חD9�C���m��j�,��+d��;�F �6~�Tv0�%G���#�����0
X7�/@C�-}�3�<c�;��kP���Az�_������ީA2z��~bMf�r��g�C�����#}_�2�3�mC8Km����������h���Da��v�f����p舒�uBM��X���e.
e��M����}[8�X"DG����|�ɚ��� ��>_D�(��L��#.Ч.e�H1�,S�����	�����b0�sB��p���j���a)�j���`��5�$wL�iu��iu��j����n��2�<�Tͺ�"�A6��'>�j`2��%sS�R��H�f���Ⱥ�X^�uY���%�u��=���D�5\(I�~~���T�KD}��>��w���eY��������.J�[�n��g�
N1����<�󷝥�n�<��'���!��r�9k�7oA#~;#o���T�ʅ[W�ֳ�Ռ����_�h3�Z!����]��;��>y��.�/�;n��x@r��ɽMw4�+)X������7������������D�A��nΑ��4'c�/�5�>,م)	Չ���9&�zY�K@�y�#�BF��Ӊ����߳SZ�ZeQOg�]*�g�&ؿ��l���Y���;K¥BV��p���moe����OHT�:z}�)%M�����s�~�X80����>a-r�O�H�:L-Iu�xmSi�7F��t{ɩ�ʷ�.e���;|���y�S_��Zܦ%z゙c=G �"���j <77k�5U�F�K�Jc��49	�:�Z��`�R�v%��`�~�WV75/X1��CE{�M��Q��e��J w��\���q��6 �WՖ������	�L�/���y�{�����
W���'�b�b�k�8�`ِ�}	#
ɛ�r�lXӫײ&�-r���v3�^H��8+/�< M��y�v��џKLg�Z��"r��F�cq��,N��-gKnꨴ%Ze~b^"VDº��{zehhH�:B�T��ş�"^h��s�9�yU'o
_M�V4�.28;�Y?��<��泶s�AL�䪖��n�7���;��&pg��p��L�� S��#���h GI��2ꊄD�L�H�V�Y����8�)����{8���xذP"酏G�Z2<�a5��fp�g��TdA�DD�M:Cu��K��v �=dh��T�jY��EAq�6Z����(��1��O<��ņ�F{G*!��G���W�7$ͨ�(y���
FH{
��m&'�H �S� =��e>����26~���͛��k/�D#�q��u˃ܯ�|��>F��bn�%M�����Z:��%&�Z��w˦�j���	6u(t�fv�YcQ3���>�D�����{�N�~�4�\��"����u�dllH�o��r:"�m�n��ܤn�fܛ�N ���k����jt�l��������,*	ُO�Ⱦ����қ�˪UmX�J�{���3R�]\Zy�%G��sQ~\Hg�	�5u��{�V���H�9>||L05V��M���)H�@�,,f�8zO���kB��c2B�2�{���U��R�s��Uҿr��M�I1�N@��IP�`��ߋ@=uL$<�ȓ��cO�TeaQ�rԓ`�Jґם�Q̲L� ��]_��X�r��u@��dYWJ�+�"��g13������8ܥ��4Y۫']9�?���<2md��(�_���4�d��ՠ�*���,��W�����Z�&�Z�*\�����4�Q��tKHq8� ��!Nq5��KԹ�,#t$�k�"�<~�M��QQ{�����^���I����Y�W�3��kL;ؖ�P��q���4=n���՞mܼV^�K��..Ȏg����R�������[��m��������7��R�����S��7R��o`�G����G��5"{w�=L$5�kք('y�e�;�f\��!���@������D��o��1e�S�cx`��~?�o/�����$�>!S(J�؉�;��2lFm�Aa|�9t��7�.3')�y�|�~�s�A"��
�s��k�ӑT㦎+�@v��>�5f��p���%>?�[�B[��M�� �]>�e;O�]��*����֩78�yU+P���7�3�ˬbL&�9q�`#lTT��Yں��fa����PB���;��@oS���eN83Z;z��{肋��� ���j����( 0W���\N3s�et|V�֌�J@a,�D9�s J�$�5�c�Б����̒+*�4��q���~���4� ��:Hff�Xb���	#��ᇂ\�Pz���s�;�=7l���s,
��a���f�r�hs4'Srx�f���D?yn~���J� S����A��%]��5�m����Gc!u�>�br��e���eV�š�{�X+��ԴDۺ��eFf��� ��2ْs1���$o���ܪ��[4������x\^{�2�[U�O�K �&Ǝ��kO���H��H-������<��~���i����}��48�%�y�/��w�J��|�}D$䖛o��e�����iY�i�9.=�aT*�1��4"� ��u�qm2��r�7狤�� 8@F�U����C�'^D(IbmP�,]������!4J��;�����`#
}Cf�K�ݩ�oYM���7��D��@k�:�(��V����@S����'���E"]�TsR�u�ԫ[�ʡ#!�h�p�/�ЎAٛ�L�l�}�:f�5x���IdS-,�|iΌ�6�ԉt赫���g*{dK���ǩ�׻�r�xﻜ����9��'[���]b�Ɏ�83�4� ���ڀ�󇐉Ǥ�3D����&S!i���ѽRq��=w�/+V�Ƴ.�����ԁ>/�O��>L���u�l�hA@�O��W��5�Ɨ������a�G���,�M�(����a}�IC� <�Ƚ`��1�6��&��s���I�;3w\M8Ȅo��M2���a��\A�C�%��U�3͡�+d6re4����ǹ�Ѐbf�_(�4�w^��cq8Keq��Kt�03�3,+���p͸A#��+yp	D�sb$z��Yٹ��?<�Ө�A�#1�U[g��?�s#Q��C��%w(@��;�L��V�juIE��_&���iT)�y�����{�������u�압k���w�.�lX'l|���:��h
�ohLj����o��6�cO=��FD���hi�Y�n8�x�Y�(����ww�S���������QJ8� Q%9X��F�)��$��9�)R������f�R�;�4��3F����zP��ԍ*T�u�I�����5�*i r��!F����Q����yݔ1�q�'��5��B��{�����������f�$Ë�t�5G�ߧrҙj�P�/O=�[��Z�z��iKyࡧ䬭��K��n�^�?��%��y9o��O��?{X�����/Ȣ:�|�O��秞ީר_|�>ɩ�� ��������i{{���5����޻��E#d�K�Zdl|X�5�
�5C���ӳB2� ���4�Wj�ۦ��(n���=F�������a8
��e*TH�#��,��Ş"�l`i&�����Ҧ��3�/5���5ʝ/�������4��%���E���x₮��fb-��o���q�b������7s���L��E_�jےחojn^F��{[f��vs,j����ͥe�eo��;�s����_/�v��ܼ��:�7F�8�.~���a�l����~��ܘ7S%�����@�D&��jv^:R�,�́a�� ��������?ˆ-Rs�a����õ�\�g
9Y�5&�A}������׾&��?Km�����tu���������E�~���#@�@��s�`_P�ٵ�t�AC(�����Q	x�����'[S2:1m�Ӻ��CrL,���:2�eˀ�jzӪ�N����=a�c�Yn8 M����r�y�Rʲ)�2�s`P�1_\�JS4�FN4�k~Q��]
Y���u3�~GW�t��ˌf�O<��L�O��F2�M���,�Z?fب��Y������ڎ�9�lӡ�a�7��o��|���ݙh��ՠ<%��������'d���J>�({��`������_�8{���4N�֯��y�xTv��ED�HT{��~�H\�۠��,M��=�eﾣ���[���<-;v����d3%����y!���B�<;���0ea���:�9�f�ɀ��{Ftg�F�S���.r.u׾C �aor[[����ǨP7tl�:�}^���)��У?�7��J�����|&/#3�f�:u���|f5+���2���3/쑞�ղB��GNH��*I��V�H��W��%0�+1[��P,��/�ebdBڒ-���,uGA||H�A�<�� n��y���Hzv\F����t���Wv��I��c�˕�x����WI�}@�xz�<�ϟ��||LVm��#�z�Kz���ե��/=�mT~:.����Ӭ����+�����z}F�hG�q�Ϋ�7�)�H��6��:p 4��F<5p���6��fJ3��7Ǿ�'��A��,F{�x~�@pP����mw���6����ӑҐ�N3F,��6���ў� ~��g*�����tŒ-�f �?X���f����y����h���q��?�x�W�YwI�|NPb�D���={������Y3�Q�җ����0e�q��͡w�U���Guv��>����V��S`o/���֋_�1�K���O��x88�8q˛Pp�ު����|v�"G�����q-�U��>�.�e㺍j�j�ؓOip^���6�֍�Hd�D��5`�-P0�e'���~T>>9&����I�ڐ�}���@#�c�JL�dK�`��k�R�^�y��e��X,��!�g�&0s��21:&�o� �C�i ��ƄJݧ��q�B��qF9t���}��j��"��9�_wٛX��M�d	%�i-�r����I4h�X������ CB���H����L^��EhނM�'�p�ݷ����Fԓc�$I���V`B�Y����_~-3���� P�3�^�͞��N��2r�/��
5"v�E��g�a��1�;�yH���.��M�%�>(�%}m��F5ب�d>W����f.(��4�B��k�H:����K��p"%���nI�S~�Uo���~5�m��<6<.�^p����;�p��m�iW�yp��5��(,	5�7���Ї> �N��=�q�Ξ�����am9�B�����;�y���O�S���C�J1D4Z�{���<��3�_}�Fփr�7�[��^8�L���a��ټ~����]p���F�7�������h��.50R��f��XNŦ�3�P	�XA@�Н�0�����V����w�+��~�:�&���������ȸ,�Q�6 B��x����G9����n���-�R?��:�o�M>�;��BF�����1����5uօ{� ���d=�TPn��n���4б����G�T7�d��a�13�Ci��ll���o�3��`���lـTI�ff�>>Y�IKn�E�Yf����Nפ})����s�Z�~u/ f��q�?���EB&@���Ġ�4 Iu����@�*�2)Ɠ`�;;;i�!��'�]�ܺD.#n�@��[a׺�p䭪	�3�fѠʓi�� I?WA1'h04���/8󓮝{E=�J4�/"��{ �k�򚗛�-=nnB���8pP6����ZY�����ell�I2�K.:����4I������l;�{&1�<b��Ё
V1Bd�=7;M�����哟�]��w�Q�n�(�?��t��&M�3��� ��1�B���/��  C���E���t�M^�4XH��.��d�Ή�I��v��y	�t��½��3��^��ԍ�[D������I�L��3��7���rԡ`$-��@\>�7 cWŬf,vQ�k�6�^	 5�.�+l�do�+9V��/���.�l͒�xJ����±&�����̧?!�n��펍s��I���qЖ������8�[�`��>: �"��"�lWg�Vjj�Y�	G%�/s�3����� �
����hc5|Qu�P��R�Q	��,.�z:c��0���ՔL�{������}��eܱ�L��j��AjYT:�o�� f������n����!P���X��ſ2���������t��MQٵw�:>��:��<��iK�&|�}�`�bN�%��ڷ����wq5�y�����b�\�(�+��Oȅ۷K�E��������80$�k7�=�q����u��b?�?M�L%˖G�Ϸ�YbP��Q��$���E�9]C�Y�8g�9Q��*�T/����u�H�����h��q�����:9��CH��~A�~*5(�?D>��?#��ǆ'�9naJ��<�a���/�ߺ�� �㻺zaZ>u�2��~�a�b�y�� ����|�8��3����#���� ��/�\ AF+1Z\���$[, u¬2Ȓ�Q�[Q�	8<��e>�7�<#_����Ig#��q"����hQ�Α܈3�aC����A�@kR ��@;���:y3�TAYUx���u��
f3|��fx�e@��@8�Y�g������K��.ؚg�yAn�Q�\s�f������CSp9z���\?K,����[��	z��/<Y3�>���^��h���m��/^��(.���c������>��ʺ��`��8Y�0H��](�ҔԿ��;���<��C���G��iw<,Ⱦ8�����S;�%6dafD�mU�!r+v� 1$�QQu��G{����Ȁڕr{��^P��~ͨ繾�` I�FCLT�i"8�L#fᰱ�Pr�1㛨�f��`&'��SP�!����������v�0�����&�:U�)U�[�q�}*����*5��ቘ:��R��l��1� �@��ĉa���M��QC0���Y�Ӹ��S��*tBp�E;�+^Ϩ.쏪қ��'�J��ٸ)@S�ǃ�+I���fȃQY�����#�H:�y�z��u��A������ �!�5 a�:� ��>r��}Q�˨�)Nu֬�����]E.�1������YoO.�`��HC�@nR3ː�p���d�i��!�Yg鴹5�����,�P._�?p^�܏Y�@,(��I�c��}�v@� hy����n�n\�B�dtl�փk�9M�O�	ͤ�tS�Ob�3/3��rh�>Y�jP�:��\ͨ3pT#��-���x�����p�U�։_��iiь%9{�7���
�����.X{UrP	\?3�NhP����E�������fa�f	�����麁Z�9�M�$�cj����-�6f�(3�Z��ƣf\
k(���#��d����2�p�������HF%�'��z� �x�[���e��(�ڥk��=�ʞ!���VA�CIB'W�$���iA�*�)�Ѣm��(Pi��DE�bWݬ�gJ��ՠn�����6=r�|�Fv�9��j�+ȤB��
y�<�䩚�N��W�q<�"�hx8QT���cz�1?�u�s����¸�J���{����!������Ao"�>?12!_��w�?������`�����X�^�=��,۳���rG���Ϋp�/w��ܩ�s�9pاP6>�?�����Gy��w��o�K��)��s��7�^h�`-!�oפ#�IׁCJLW����Qx��h'�����3�����[���5����_.?��d���ٲ�AR�H4����c]@,
\�_l F���(9֔�Do~	����C}*T��F�$O�u頮�T�[�qX��>�3�l�&f���m��sl��EG�\+��p��'�g�����������o��U�f J���_�Űj�j����Igwi�j0�T�13�9 ���@�r���s���*U��7��w��9t�����4k������Q�W42���1������$�eVD�8?�����q#�G@YD�?�3r䬨I��� )[��t|��Q ��v\���D��k� �A9�mAs�����4SG��(^�}#မ�%�s�lp]�@��P����P޵ɬc�+��#����s'H���p\�Z;���lk2?1+�)�/�i�!D�T'jyF�4�~���fD�Y���h���pl>�|iҟ���M/���O��qނ��)���`�F e�B~Q�[��a#�6��^�i5꘰P��w���9@V���PDX2s���=o�6^�y HY,H�P�#'*\ϽX�rv#Eҳ��_�A����	I&[Yr������v<�f����i�����v���`�H��_�j�Z�ā���E�>v�����[Zu� �����C>@ ʹIDc���=I�% �ՙ;��B<��k�
�j�Q�R;�FVg֡x���Ŷ�2}j��?_����1�!W�v�`�bYZ�)�y+h����#�7�<~�o���Ai�u$��'4��l�ZNA	��bt�Q.��'��E��~P9��ҮAg|���-R�k���S_��s�"���h��-���d~:��Ws������t����O}?�g����?��N�o�#�������xB2?��]{�K5W hHbqӳ�tO(lT'�d��` ��������Aw��Ts�ۛ؈7EerbFң���OZ����P�Ab!;�-��G�� ����Q^�:h�k��R��D��p�9X'��3<�5��F����`�Ŕ�յ��8*���X���9���|�7 �M�3�b00�_]�:9����l�mut9�� 3�[���9��0��,`Սƻ��e�ڵ��:D����h0"�B�=��V�@��C�����l��tn()�|˝r����(�=.��X0�LЄ���P9��|C�R�����J?0�a��+W��G��n�dg� b�g5F�tu/���a�# �eV͘A�P��R�Tɩ�T�!�^9#goY���Ha�0��k^�Cd!�>-��k���ޛf��%���icA���Ϭ�H���&8�(�!u�(�#�By-��D9ev���}�~uZ�n?��M�3}L�n�-�V�H[I?o�i&(�<�y�����K�B��������	ȩj�������L5GcU�s�4���/mb�d�4}])��~]�oKv�� O��l?o�$��y0� �IHNP�A��f'�Q�.P֠sZ��<�p�1�L63��|��[7�s.��i������k.��*W �5%;����Te|��m�p�=q�k:��9\�;ٲ�%��MF�iDb�STK����aٸq�|��]+�z-o��mf�ft�;�%��9��5〮��:h���R�2����,m9�{�Е�{̃��'�6+@��TÍ�����tT%PI�߲u�x%Ud�x.��z_�&�P$�qXz�"�:�D� �1��|�Ba3 H}H#x�4��P�b�+��z����c�/��c��;l�	ۜ`��	]!$j5��7K\��w��r��Wh0?��rqO�����=��[�����ڂ|���L�L��=`��@��7�����w�M�Of屬��M��\�d�x�{�(Oc��H���~v�B�P�w�3�����q>n���A#�P?�W!���իeB�5�/j9�Z�q=�����з&��@8���F*���~yh��Y�:fd�p&�<���cBb0q��
�w�9g�|351�Nb��}����I�4�>(;w�f�d��<d�j�mK�#>0�3SR��	�
�&؇��a�3֠79��A)�Hv$d�,ۨAA|�p�0D��Z��d��0���C��,�TMv�r6�AI���<�'�h�� �qz��"?[�Rc�X��5�r�7zԩ��^+��>K��8�sjI�\p�A����1~�E������{D	�C�e�nz�5Ww�6c�lTUe��57�zM���? ӓS.�JX�"U�F�p�/`b�C]M_#ՉѻN+$�X�������M��)��֞>�G|�
���)��
��Tg����9ÞIg�k�f^������6�����.��������T|���"��z�*�h+�reH��UHE�Nra�2��y���5j�h��yn�\��D�Ct��_�'iJ�ؒ�Q�$+�}���k�sV���pQV�j������ww��t�-�ɇ��	���v��Z�����P!6s��8c����%[��$'�q_��S0z�����y�l;�d�,w�{��?0���LmP�z�af�]U3��ڲ\���0GҔ�O����B��"Q��z��SE�<[3���d�IYn2���G��S?>�󅁶����c�ە��1" �2��GK��V���FP��Q^��k���c��
F\���;�9���wv���u�qǟ���h�����З�c��%^��	;~����fPL&4ǈQ�f�2�0'�&��M쥟{�E�n�
�d�6�W��z���Y�LQn��^Y,�5XL��ni|6L'h�`�>S���A���?��;E9.۶�+�=O�1�xB7��jܗt����ҳ�px�̳sF���HĠM�}ԤAl�6��|Á�d*0��J@��Z53b-�&�y=�CA���V�6��\�A9'�Ͳ<�y43����	��U��<z�׼�=r饗JO7��06q�րx~������H���q�hD[R25��x�f�&�/2w��%�R�8*����FK`�Tk3˦�D�udy��%rxco�Ը�߉}�E���w��� xr$��Uh�k���x.4v���ɽlݐ�`a{��E��eu����j|RɈ|���L���;"�òM�:0����%���<3�L@��:%�
IKKI��7�i�[�},��%a�9{��u��M�&�ɵ\iD��������]��s�����ƍ��j��NH�f��:���R�srh�Q�Kщ G��z�Ϳ|�\}�er�}����c����Qck5Kb�V٨�36v!���z!'�cѳn�@gN�O#�����\������k2��A���^"�A��v�Z���4�����1^����A_\��z�p�w=%��}r�k��5���wP�:������'��4�z��}296$���L &�n�
�����^�&��o����SY�j@%�(��N���2�ٖ!�1Cq�5p�C�)��@��y0�vC��)Q�����M����@��'L֣�>_̸��V�,kH�f>��Ջ��ӕ�OBQ��I�V��o2$5��کS��*\p�Yu�蹑��9#y����~�
\�Sɯ�D#�L����=��a��i�d�1��Q��m(a�D�����H���,��_�����/⤝WY�x5�5�F���*�;�2�R�%�qh#�cFr���ֈxka������8(T?@�Ҭ{՚c��~�d�h�������'%���f^v���}� �\�1�F� ��]� �BPK�l1�O��?�2��H0��_��d�p����bR�V�:��@ f8O��<�{z�9t'���O3tu>(�Z~�Y�P0��`��eN�0�MM�I�� �z�Z������R����ب���S&g'��%!.�����?�O{�1}�Y�ܶq��,�ˤ�=�N�ʍ[f�\�:]H���"K�~��Q�Q�F������dv���a�M[�L=rq�DB�k�����%8' )Q�(�3�C���(��e{�HV�������KW��52f�詪�.�P< &,�e��C6oZ+��ݏˣ�'�'��vu"붬�cG�������,���a��XIs�ȲVg��\����`�a@�6JN�7���6ѼG�� ��S���3�qL��6�$����lDWH�_����#��,u�����ɇ5:�ށ���_�F���s�o���c�?%�LI�S�z�J	�<��i}����7��Č��h5�s�Q��h�*Ő%kV�ȝ?�Q��'�{����RM������fU�:��4�ҡۣ������\7�����t*(�0cޖ��o�EοD���=������dz*ǹs��ܿG��_�IJ�y]���ӿ�I��Y���>&��,%�p\�{{$���g�Ҹ`s��@����5��g{S��5{�:*b�B�LWՈ5�o~���+��cǆ䉧�&�m�%Š��l����AZ��r�I�[n�ɞ��J�K%j��6��U�`���n� m2�	F�#��nda����^���D5 K�a��,�����bt�$A��5�XA+{Ĉ�~�X�i���o궽����σ��_B/������� x�����{9���W
�՗~�Ҳ4[N�WWZ�}i��F|�v�и^��T+�(�׮g`4|b\z:�LƀmJ�D��)Lw���*���6)�6ey;�v����h2	�D/<�*��Ԙf�a�I�݇v��p�G��50FK�8�A�t�F�ճ]X��p{�hEA�jQ��a��}��j9x������m��:�$��I7ġ�ı5��;	�=zG?K��+�j������l#٬N�'���4Ni��?�&ɖ�LN�����Ɛ�����P�v��#F(����v�se��u��Aw̪P��ؤnh"}��r��A2�V���YU0��$�L6p�.�̜~�4��@y�s�Y}�	j���b�hZ� ��d�N�iS�����9�0�0�.�K�i7������x��/sJ�V-�{]�W\�Zy�{�&���@o�\��wjƲ(����d׎���S�S?�sp����F��"���L���\6��� U����_��l�To���Z��ݬ���!��`p�O�2�l�y�1��9g�-�gI���>�rW�9�z[��He���=�>��Q�9�[��!�_�F�__���r���?��ulY��-;v���f�K̀V�������?��M�s��������jND�:�M���;��vI���������ほ�5��C����܂lذA.�~�ft	������N���<'����^��K��M�����}\N�XQ�8+@������ryٟ{z�|��׊/�$7�~����S�9���5��>�_;��<7F9m��9J�a4��WM�C.�h����U+���	��?~�ճP4�׻Dq�pS����YE3�d�tE#����`��Q�ٗ�"1NЌ�V]42Zq��!������t�.>�h����F 	c]s�
^�nK<3���5st�UE]�����9��v���6=Y���Q�5�JS�w^9�~~ �z�)v�i�Ա�Z׻���X^1�-�Oj����@o8.$0��Y��#��`S�;J	�n�Un��;v�2%�*"�'@<��"+"�SjWú�sY�G��l�a�x��A�59��W���<D��#��ے]2=�ր������UW]%��k�&��z+�?��Z\��}�H�t�}��
A�k^����y�x���|�����y�Lk��Q�n�s^v��XP"!�p`8�Z���\����k�B䭏�Qd�]�G�Z�Foּn����������4�����(7X�|��p���[��M�����ɕ�*J#���$�%I�����ԒF����\�֖���s'��=)u�\�e��$4�h��-�c�m�H�̃��/��r�j����oX���"��4Ш[u�r (��CZ�%�����Ɛ��7,�+�u$ }���hNh��g�������kF����gٸfP>p�{����Ѭ�c������,�q����R�bx�X8�e5HCp=a,����@O�?�����@�g8}S�5�:��h�Ɍ�����2YfYS���u��1F՞q�kO����H(���{��ٿ_F����G$L�W��m)��F����ܧd�� G�>��+5+�=�����db�&ݱ2u�0��`L��Dz4x��������D�+z���L�jf���Y�)�,3�)9�H~r��2;7/�6����HQ�bY�]w�%7��5����Eo�Jr��[�W\&���;,�]ݺ�7IkGH�J��S;\�r`7C�)狆xG��?�w�#ܟP��,<�aI����:EK�
x��1ޣ�-������@�D1��
%9��J�Sw��g��/)�⢨�z ;��ɬi^Ay2�*�>����L�v��0Y�@YQ�uP��!ڄ�:(��eA��k��>}M�Ђh�^ThK���p�Ñ�"��V���U����ߝ��]F��4s.'�����T5.Ų��Rǩ�t��9�W|�[E�|�H��$��
� 2�~~&���i �0�U�dr|B�b��i08�/'N�mT�A��.�>8�.q������<z/`��]F�k��]n�ס��χLߣb{��~��|>�=�>f]��U%���ׁ�:�kݺur�e��B�y�fy�o����p��� 3�?�5��q���v,��4)AIU��Z�3��P֪;�|���?�|A������X>K0H9��4��ŝ7�j��hnmf)�n����iPeB$j�y��5����mWO�#>  �H�r���SzD����'o�����-C�G�%�����9���
,�:�.���sb����6��@�;�v��^��zd�D��cT���%S;?._���Ƶ+����jy�\u��埿�O���(�ȇ�׾�}U�v`�P��;K#N����nubeWw�E<|�B6C&�֦f^G���`31���@LZ@��*����.�
��Lg�t� #��
�2I�335�����f��;����cc�~���Y�ܟ|V�AX���?�����a0� @俁bsI#��~��{!��)�@{������ ZP����D,�,�Q}��D�}�,�f�{��n�ZY���#2�ۧ�z@�zu�n���&��?���r���e�/��y0�8���3;�s���0����$d8�15��hF���ci�DQJ�QH	#Y�)Ⱦ4�>?���.�ۂUF�h���vPs �Z�aR"*&Uݸ�Ь�9[�����Gá9f��cG�W��i@Í�}�e�u���YH3o\8Âh�.oɰ������J�t�Χg	�*��{�pl| ���?�ܶ�v�:�K�ʱ��7���9u�|i����r}�W
��X^�`p௛�WJ5���u�L[���EE�1�^O�U8��b|���W�g�7I�GHd/@�}j�xA�8���#Ң�i����G;�5���>���X@v����'�oS�&(0�.Q]?\p�>F�L���o����g�}�`�t_8׫63��)��Q�:c{��_:� Y�k)UȐ����$��Av��w� �S������a�afzR�(Y�߲eJ�;�锣G��`�H�ـc�x�j$��U���
�/eR�V�+t�������M�2̈$��w��`tc���U�{~������S�`�f���c4�~C�A�2E}x��G�4ԍL�����Hⱐ�g��o{����?�亮;Eg~�M?�ǎʿ��7e���rx�n@8)3Si����ȅ� 8~&d�IS�G�seނ;Fd���8'<>������b�Ҝ��^�%��0�H@�U0�a��BoNi��Ne%8���e(x��v�ʕ��keӦ4��׭�ݻ��?�ӿ����/�SO=#�<�����ۥ���5��Nn��.��b�J���WM�"Yր���E����zݤ�L�b2>>�k%/��m�n�j����e`�Kz��(��X�������q{������y�2��XȮ� �>�)y�����T[L::�ȼ ��?�!���r�2�e,Ue+'��*`4P�H3�Q � n��R�]��K"��� �	����� p�wؓ`�3��Ս3���`$��&:Ǫc�n���hv!���W)����O�{�Lo����X�PP,���ĺ��Z	�+����̚yϸ�2����T��ӾTkM���T{�;�h&X�E���s�=Cޛ�7�5VO*���d�u���q���0�myN���+d��.�i��+�l�>����8�@��J���	*������I�I��_�������ft��f���G]R�
�k?BF:�3�����+�U3����
T.��@�W��i'f����BZ|���(@ q����fE��5�����ͨ���<��ݻw3�K�� Ne||\֫=M��˚5k��X��=ỳ+j\s��8��󅬀?��$��s�h�2�A��s��wP^6��j����W�&�1�S��H>  �	R�6���5v{��e�g�,����BJܐ\���4q�/�Q]��!�+�X�"2�"�Q��2�k,����l��oQ�J���+�ҋ/Q�|��tU����py�9s�"�����1�l���(�v˚�J�PoE��귽U�x�)���/~V�{�I���_�w=G�}�q9z�t���I�J��[v���#ǀP!`�����y~. �q�s.��(�.ʸ�Gv�7�x-�(k.������0|s/�FU���B^��)+��
Y1�QZ\�+΃�5(��Ip����רs픕�rӭw�]w^.���"O=�4G�n����w��O70�~~��g�N�P���KJ3�yijN�~��&�0#?�3�/���|�Iٰ9�`-��bF��:��ML�I�`�<��}j�*r�5W���̨ƿ*lߢ�.-�=�������;����*Y�z���ʫ�p�̤�E3���M����2��^o ����e2�C��q5,Vc��>�r�,g�!a-�s��+�+���9[̡s����J+�������0�s�O^��{��#�X���k8n)��2D0�\w0��C�2�Z�d�����6Œ2�5��Pf�t�������֐M8�^����߱ 8]`	�M��m9�3��3F��%�:��疱���[����t���W>l1�#v�����]u=��S[��I[KB�R�b[�|�%w�!XM-��
8�r͌�Z�S�'&�9�0�UB�1����Sws���o�4�Ô	.2��ep�������Z���� ���:���qNS�w��d���:*�o|�ٞ�������Af� Wg1"
;۸6Ι��5ۤ�U��pYR�W����`k� ���"(3������d?C&��l�k��!��܄ �?���׽浤�<����?�d.@ s$�4�7ٿO��dfnT_kNb��0��R;�tq�ca:r 2�ۺ�@̓l�` (A��:΃C_��x���1~n(�A�j݆M���ˈ}w' f���%7��T����x�{5�y�%[��?��Ҭ��]?�C����)j�u��eQ?ߑix;5�#���fI����@������c\�6n��s�ݫ�d0A>�F�8�2d�N8�ӈQ?�Zk�\�<������8`0�ϐ��uӛ�(n  ��X�[�y�U���ϱ�s�5W�����9'6����V9�V����S���;���/�[�|TVm�&3Y)U5��e�����;�J`Їӯ��$!YXX���ɡ��$�)��W81����d���NKk�I��<�����f3Y��G#��:�O�������FVɟ����n���[�f����I��w>���b`�ſ��@�����^]�s4RXo�f���Tث�ʑ �Y.�΍�H��ڢ͂,�����G��`���� V\���w����>�ӈZ������Q_n.9����S,�I?5������R�W�&LJ?��P�@�WB�\5cz�;�k�����+��k`�3�=E�"oʼ��lN��,?��h+�Lϟ��F_��W������d�\�n���{ٹX��5��4��r,ʟz�_�/�ɢ6��ܜ��Ao<�1�E��7��4���]����.�lV�Ҥ�$K~
�p��rj�`�)�re�+(��7���Ԕ��e �}����f�C�Զ��Y'�=��ڸn9rdVJu�q$v���(��ٳ��{��^
���kǣ���ǚ��@`�qU`{�X�����w�E"&�n���n� >����8��c�}N�+�Y���l�YG� �����&�9�y��J/@FoٴV.�p��w�|�ɧIq�ȣ�?���r�Yg����+r��ˮ�;��]�p`�
��`̡��ӓ��n;w���&d^���c��t8���G���h�QP>bfӔ��E�R��S#�x2)�}������%�����F���������eeq־����5W��;n�U:Z[�W])���n�Z��YI1�Ӭ���e�իWs��.H��`��-��8������ģ,'��������#�@�Lj	Id�!�ْc6�-�<���詡��;:v}��^m�ԙ@2�`���e�^"?���+��.]~9|�tu�4��7��
���g���+�"w��$u��eݸup4I%��k�@-�e�P��$h�e"hCu��8F�ǥ��]֮�Dހ�C�253O��.�V:z���qY�f�|��}Pn��F�֬�{������1����}^�q�5���!��q���G7��}����_ҙ�^��d5XF��F&%���
d�3F|��in�m/�k�p�J�3@�h��Ao�d�>Y%T��%�q��^�j�d�/���a���r*�_t&��Yrx�q4���U3 \�D��BC�- (C�Ɖ<�0�g� �|�,25Ԙ�7�2;*X���x�qԤ�`��pT����`��䆨�b��f��7��+�����S��~�,�SG}��d�n�ᘵ�s5�D&�zݭ&r?8фdҳ2�����	�/�J��6yh�æ�Pz.W1��n8tϑ��o�5�m�o|㛲�K_��|�7���jDN?*ɶV�B=;��&d�o��w%�U*�%�4�$Y���Yr���La����wwtI����Y�}��>+�tҵ?��m7�Q��o�$a��`�lp��A'�_[kJfƏ�	C����/Ȇ��`"�,����t�,��n��u�[��ѣ�����r��Q���F䎑+�����M�z�v�����:�����Srp�~�z���{� �\�ƾe{G���3�iV�-qJ���Og���ҡ�AX~����D�XG�q.3�Ζ�<�k��z��Sq���\���s�٧���/ٮY{�N;ٜ�4+�g���vuq��y�r��1�p2K�]�(tyQ��'�V]JÔl]�h�p�c| � ʹ~J�Ny����ܝT?ù��Ȁ&Q�m$ɑF)��hi�r�ߌ�����4��`nzJ.��r�n��}�cRÌ�>n��urbdN�:{妛n�7]������ݎJs�C�̓���ҡ����U�����F���}2������8'��?H���?`��16����8g�'�O��z�X�R~��7h�_�/��ۏ��os6���p�����ƛ�#C����^�|�5&�A����@�$y��T��)t�f���/˥�tܶI�������S]n�k�P4�lz+7n��/��z��4�5q����~x(t�2=0e���QN��O9N|��3ju���&:wTʝ�@�����#� r�B����S(��@���"�ȂK��K!�6%�/�d����������,φ�s��F�޷���ۺ�	�@ 	B �@xzH �M/!!	����ӌcp_��z�����J+�V]���s����sF�-v�_;����4�����u_ł�p
�A�ɨ�ݑ��,Aa�#�T�cZV���;�]�A�;[����=��z,ͬ�ރũ��9�GO�Vn<�hU���D��prB�Z.5�/ۄ_}�͘�>��\3�c�j�����܋���L�d��oZ'`�^v�� ������qCG��G>�Q|�3��������$f#�9��c���>�e£�������F��.�
�r�/+�/��� ���L���v��a��x�#�jY�t�ؚ��	�@��0$W9�yL�WN�jZd���)�%C*(Ukؓ���J^�oġ���o��������7����i�i�1����:��"&��,��H�q��mjIJ�ԉ�.�(ٹ��lZ�/��f�쁟`׮��9��g�H�N�N4�dP�����Ȗ-�$�š�`l|�̸;�R.hVkz���fv��Ln	H�P..���TS�5`ٰn�j��MO��+.S�����l޸I�Rܤt����hL&M���]#��Xznz	Db1
ajW%ױ�Hg>�
H4�}	r2��Ȉ���(�gC�D���C�FF�Qa�^��K�u�-�,)o�k��xFuݚ�8qr���#Gɪ���|NW����c�sr�G��ӁGF�ʓ	v<PRR�Z�0b$"I4I/�\���N����7��J5@T�:t��4�!:++d��Ljc�7ްJ�{��ŁC�f�z\~��X'�ƞ=�0r����=���_�Sxr�#�ƒ��i�5�^��w��ɞɠ!�|5� -�c�&�8��U3V
4d�P���N)��T��1�q&8��Q1VCǎQ*����ktO���Ƅ�e�̨�k `�������c��Ѻ}��Z�0�X�z��@-��]ԍV��;:�P�X��W�����T�� =�ܸ�BzLmY�Nh��6�L�.���3&#�½�3���͈&��KIxF�����[Y���k@�pC�-Oֳ����;T}��}
Ԑ��A�i�D����`ܩ����t_t$ͻ�������_J�c85�U�U�*���1��6�?�u˾"�����ɰH�+�|th�=��C��?~��Ӷ�k�)^D7�ً�
!�'E�b�����S����'>����?ф��gwbՊ�j���W�n�?�>���M�~�Lq��+�1�߶wtbp���\'�HI�lҳBҙ�؛`c�j~pr˭_��+h�Ev���G��,=�AE�k�Ϊj�HI�@�Qnb�P��)ƱW��%pH���׾���]x�G�u�8r䐖���ڍ��v�ɦii"�!��ɴf���$��4
��D^)-���t!!p�~[�R2*�_�G����]��.Y��MQ�!�܂4�,ӒBu~!�XS�8m�>8U:�R����44Ĥ�%Ȉ��̜��f� �G�ӵ�a�M�q�<&��(-�M�������%0$ƺϿ�W]q%�gR�����CX�n!%e�74֨Xi����uk�;���1 ����S�g�ٳ%5����e�L�ߐ��m������gYwAK��?�gVʋ�wǮ��y�~o�A�ɬ,up|x�v(��K��v�z<����Œ�NN���F{W�IPG�2<2�_y�d�� ���Q��Q��b�dvQ�hg�����::z;q���Ka�%�#=;�-��Xz%���7߂��a�JFΙ~f�y��������GP�o��w�s�&	�d,��+�O.��b�<���薠��f��J�)�Аl� 3/�/{�m�@�*�����
\cV' '����u6�Z�ZDK{�<�\�ܗjP�	����U�F���%�p��^����
vU�.�� t�4��+:������Mׯ"ycWZtf6�C��`4��/����T�m@s�r��1����a+�����~fj�O�L��$�	��c�uu�<)g��s�sU��?>��3�`�̹}Nep��lrt���O 3A���ieN�9'kFP)9�ٯ'�;�qTo��]A�l��
9�Se�|���}N^�����AXq	E�'�+P6A1�>c��/�aא����Ή�á�9B�����_��{����%�[��(��!����&���h���Y^'NsttL�f3S�H��[;�䳻d�5�a�_U�� ��A�cV9b_�VT�/��ܐ�������?����η�?|�+_��}�u<��Ƿ]�A,|�!r$�E;�s5tw�H���)���3������Ԭ�}��)̤g��߅�M��5�����l�B�������{h��"2�5�m�*��cg0p,۠HY�g��S�~VPa)S��ߔ&2��p�-�5�Y�V���>��7�ǣ�=�e���u��_B�l�g�z���r����\���T���h��^��ة���ᆛ��X�E��2��i�1s�q�ˍf����$��,�?#�C��*���3oH(:R˂r���f`�'�@���rӳ*aՕ�4�c	�h�*�hP�\.�����{���'��4��z���4���k*q�����*e�V��G�|v(=�r�h���ѿ�\�|Y�# h�Y秽��]���Pؾ��'*l��0%8ҽ�S��>(߃�"�[�@���F|X2��5�e�eӔ_lU��W����:5�����ͯ�����'��Y�(��@&K(�c^Y���״L��ա���),<){�)�\�;��.ttu�;w}O�3>��������g��w��d�̦敂��1����,�' �����8�=���"��X�v���K9tt6Jv9��%�ɩ�!H�R0��~OQ��|~��r��S)/2��~4��3J��ݳ���G+,4Ǝ�V��/Ж�KP[�`��G�cB��w�ga����166� ���U�f���'�������}���6�)h&sc�� K�j�p�X-;#�g�aQ=��;3u��y֝�����G�8i�j�i�NDGs���C�{��vYm���$�����Ri,`(��=�y�[�M��� qgM�g9��q�3����+
�7g���H/���
��w<�\�ͺx��q��g��%U5�=�"�I����|�Z��
7uR)V��퍊!�b�)�����w!5=�U�������8֏��� ���Z"�� ��?��o�L��Li��mW?�kg���۪��Q�ɤ��[)��=)���iE�fq^;��1z�KvY���np.<icr89���0�*��T���B��DP����Ġˡ�nC6����.�\��\O<���^�Ʀ6mلG~�R�����-C�ʕ���2�N���Y"��/�V��D�=�8=*ƸՒ��{UV"Y���L)��;)gdg)�)�`��9yҙ�h����2O�$fϊ���us�:}��Xvd�Tuk�t���7�4S$�l��SCi
)q9ߋ��=I�z&F��f�k���$\ѸK�m��U�����w��;�� ��vW�D=�f|���J ᚹz�u<]v��'�X���3j�QuN��\CV*8���14�w�,�ќ �߳�q�L!%�E�l['Bl��ɏg����q��W�?��Ϙ��h���Ù��,��(���3�Mb�x`Iz(�B�:(s!���mbR�F�*`���O!Mbt|w��uflb�?�.��Fu$�5���Y�;�&����K��t~tb�\u����a|�# �7v����]���*5��LnQF�x���f���8Z����z5�}�z��(�p�3Ǯjc·se[��N�Ì�����6������Cc̈�L�:���I�c˃���hml��؈�:{�5��=�1=U������5�:^L�r���S׿!Ø�U::`:���	ؤ0��%5)�������]2�L��g�gj:�mm-��T%,��C�
�do��>��y���Z�k����¿�}�^�'^�8��^��s���{>��EV9����|��QI2�X��O�uN+G^)�{���1G����G�ֶcA�"I| hr ���y�p��\6���w�Ǹ�ʋ�������q��>��d��z6�:CDm�qa���_O�e�ޫ��� ����)lf�u��$i��cyb2j�B%����Wm����[R���W����m�d�@Y���2��K�ނ|-����W��*������sӦ��p׷�FKg+~��O�D�HV��ڨ������>O���Өɖvd%f���I��~(�A\�up�lBf؍��ᘙ��9O�O G߂���HLKB�����]�DcB���\��-�|~!+�"�97�A~��h4i��j�Q��e���*��=N�]!����dF�*x�Z�&	��Qs�-/;�{�QC{��O����Q�����p�\i\���dDk��Ѩ�����`�RO�,�'\����h�_)kb&��}�LV#�,ˮ�-�I1�a���4��p*�}�\� �Y��>��U��`d���o�h��[I�m���ıW���R"3Y�����+V�П3h�k��)�>T��~z�}x���+Aay�Q���W�:&���-�2`DvW�`�Zݍ)	��E��my�R�����>g󯸲�s.��f-v<���!��@TQ�s�*�>��5[����A�}I�R�J�&�Y��4�l]�`~|D�|�8y�����س��Ԝ�߲v3.4)Y)U��F�!5qA	��'Q\��[��#�ա��q����0�ňRg{O~���� 9������/���މޕ�qztԔ���@�p�D�fW�f�r��~_�GMT+ � �b�g�*꓆	(g�N����$��N�#�y�r���8���y�����S��s��{��c�Wa0x
�}����Ne���^�C�������̌��V�^��Q\}�5��m��ǝ�d@m��kyS2�U%�m�Z��+�I����Ɔ���c�� ���g�!�̽������&��=cW�3�z{�W%is�ۖ�ۉzgPX���d��G,S�T���>��|a�ܭE���8�Cg���Eq�pt�A`,$Y��F�O�}��Чv<�DK#��с���MT���9�V����N��mm��?���Y��Y1�MH�]̧�O�	`��P�L����ظq��/�ڻ1xrH���Of&QT�����I�b��AQ�i�_�U�ԏ?�S�����o���̋���y��k)�T�ͮ��u<��������(T��8l��M�����'šR��IQ1���D���I�,$`���<�T+��A^�0}YT���W�T���%%w4f��=)���L�a){৥|㖁�NfgQ�H��c���N�>���}��,S�^����fU#j�g���!Nڲ͈Qv���J��i
Vbd��q�؈"�e�� 5�Zۖ����q��j��]�����s�Q�D�E161���CI���g�ٽ[���Ï�K_�*r�]2��v�r0���2NQ�te��5��. ��d �l��c;�8h�1c(X�����ꂣ{H){���Apv�>�l���GMD�x��bu][����8�@���n�r\{���>�:���i]���b�s���~����>=.��m�����_���2ZQqa;!YRc��B!=�Vq��E�x*�KG�[VΓ�:���qU�{�,��A��Y<ւ��	�����"�<�ln�W/�ɓ�r(B����FU��Sc�P\PIЛo�[�^��|��N�~��(.�a;�Y�#㩝;�b�s���t^��\Y���K��M�?��p ��!�;�F6u7]%ںZq��m�����~�����S����BF�A@���m�*�E�A��HP��k����b��������^s=�zd?"L ��f�;�h,fڡK�/����'g&��2�4��2L���õ�������
�c"�ܳB�K�ⱜ�d�O�dk���s�c0�����>�0ԣeW�Z���CbLG���h/���yq���FZ#%"������H���ݑ.���ɑ!e+��Ќ��o��(�����ถ�9[\	%ѳ|��&OON#/N!��+�S��C��������O�F��q��+N�]������#z�5�I�ߩ|�=��F�e�6��1��
� ؂�gn�\��*kY�*�@��Z�3c]�?�2@"v"ʬ�L�%v���,�8#*E	+ȥj�R�v�zQ�_1�A8�3������ޡ�cQ^$�G�Z���߯���x|�N?����33�%_=>xS�4})�E�`PG����n��ؾ��iΨ Eت`6h�x��ϑ
����&"�Y�m$�I6�)�<�2�J!��&~=k�o�h�[	هyU"��ʁ^��-"�ZU�kn��mR�a�Z��[�x=�z�����z+���º�1����r�/�QKJ�z���kȠ�s��8�x���X�v���<��#����1��H4��C�10������>X�,3\�Bp|ө����܏�/����K�rn�!,�H������]xRr�)��������>��]��y�/a���:���mسg���/����c���׾���lۥx�+n�׿y���:矗L��/�� ^���T�R81�{.�B���[s`JK)�bUz ȹ������o|�m����%�<�h�)�ĩ�2�~�*|��"Y=��w>wǗ16>���n,\C��#kz�����8�ۙ��|%�}XK�?�#ۯ/��;Ŷ[,�\��?{w�}7^�˯�Em2X)�uY�}�b���T��g�j��W�4���>N�������A_o7��G���ӧ�%�s�v�
������:bJ��/�ʠ����~nۋL���q���碚1�~��_�U.��!��*�Y�i�Mᾢs�$�k����*�Ҧ�������D�F����]s�Z1\%���uvnG�Uu.Fی�Z��MO��9� �|1���.-1�h��R��\!��g���=�Y��ۑ����4�$@sSV�]'A���ʟ2󞜝�F,l�E��d�V
�;N$�Q�ʆ�sR>���3צQ��(9��u�$��{�|�r�?oIeW-�9��#���Ū(�R�͚��C�X�a3�۩T�:W��)`�筗K5�a%2����e��q��?����ǔ*f��ٖ1�U�����h�t�Ji1cw�Z�^C�s��
j	�lUu���T���"�@���+��}��!�+Ƒ�}���l��+��L
�L�hZRW$c�^vl���+:�e2ZVy��$'���(Ū��0;� |�K3wb��-����bsQ+,��D�Ɉ�����c~_��CgO+����%c;�",�O�رc���i*� 8�A\Mn��8tz�MA�"N3,[����(���kh�U�+T�����'��{������X�Kd��TU�X���(JeL�l^�.�=��\Z"PB���.�P����Sش�df0|� F�B[�����W#�pl�.��D05|Tň�NQq��y�c+Ҡ�O�B`/-3C�F�b<�����8g�F!��$�nL�05=��]H�M��%�w����.q��u�xn�Uؾ�IY�9u������$@L�fѺu-��������|*��r�4� O�GŹ��������sf��=�� ���/2�����yn���$(�l�6]�[o/b�8ڇݍǶ�B�8c�q�h톋��ы�S��|�fL8"{'f|�>Hf��d ��h+��Ը�����:ɾJ�<�n݂ɩӈx":�"�:�?["Uo^�/��;�z��q5~>*�m޼Y�%G�����$�u��\eB�� M��sl�v�u/8�N�ܪ������3A�s)�l^�b%^s����#�s#oG ��Y�c��D2&���cʡ������ҭzC��zt>�N��e�Z���� ���Iq���V�Y^���GT��P�d��Ƒ,{V6�m�z���g��".�����gǓ���5>�1Q�d)���ŉO��~g�r��%+K�,�r��DU�qH6N�6G����g)J�Hj�'v<���M��|3bHڛ����+��Z$�d�=�`k���P�Wu>�S� wA�t[���z�<J%Z�S��ԕ�-h��:?f�v�(���c��@}�� �+o���ZZ��xrzF�⠒$�0o�)E�d�l{��)9\ش�"�����GR.Td�8>e�~�rI�@Z��f5F�S�H�3�kWGo\l�pZ�	5�>-h>��
�ECJ��'������q��ʹ9��H0A�9�?�^}��T߽��G�id򮖋5�r�C4� ��c��iz~^�C����$��s�[ӣ`��P�LTT����g�bZ�xD����}���Ls�!*��'��ǰ����y�܃+/�(ge'��o�ᵲΫ1tL1	��]�Y.���7���[�H����mـ��4N�S����>�O�:�f��(�8�0�@4����F��)���q��FYT�'�ȇ?��
l�YՃϪ.AE���$~�������t7�����,[wq�>��~t �/ڊ�{Zɐ��d��M�I���ښٖ��·{�T6]$�Ϲ�O���p,�s���x�����R��'O���'�l��a�5X��Rq�Jk��ONVq��g���bqLU���f��X�b&=sO��E��&gdu9���ѣ�����V'�(�Ū.���������W)j��(����ӃmW\�?'���oքqϞ]�p� N� ����u���}w�Ρ����Q�����7��RE��#P�+���].^<JJ����Lp|Ԇ��NU�8s3�b+5 �!bј�`� ��C�<�	*�L���B�Z��X'��"w~��H�	�4�P��Ł��fAN��d�y*=�絔S������GW�2�����A<���J��̜ ��l�MF,&֠�_2���f4�$a���5%12r�ƨD��Rn�$k��s���Y�N�BYt.����$�Z�`v!���G?���O) �<�dFb�Z�B(~#_��MZrg)��7h��<4~�=�֌���,��F����G�J��eD3��HF�bl���#g��s��AR͞��{Z,S�� 6��q�a����1�#�?�<�=������ν8%�a�M��0(�|D�(j����&ѽj�����dKh�c~V���wf�9%�	��&��}@w�V�q�'�'�$�]��������)l޸��lشQ�3���+vY�TZ������x�/��I������?�����)3���C��d�㚖�&�	ئ��}�q�T�y<��Q��Z!��-r]s�ֱ��"�*�H4��1{�|\�:7�`��!�$������s4ֳ�,-"�)#珥�h,�ɉ!���^��]���q�|��� #^6_T��=��O��V�%���gM�!�`Ҋ�K�������7\��z�{7̾xPI]�N�>ԡX%��������PN��N�k 6jga�TL���	��Y��翆7��
Ժ���ȹ�*��v	�5B9��-�}�K_��Μ�`�5/Ξ�1�Qmo\�Bu<{Q��|�|��O\��V��9����w�6V� u��N
�qm�_*O�N�8��gKz~|�vD�\g�g�{a˥I>������#�J�K���M��}(r\�=q7޿��k ��"&K�L�.Z�eX�LIEt<nr�����,�3��>���+Q��8��$�g�k1��If�'���	}m�[��J�+�}v�|���P��H�h�k��1����[Ӈ���F]�F|F[k3r��")����j2l�5�(�J���譹�I�&%P9���k"VEB"uru�C�J�k����@� ���u�%�Y�QO��^A��"b\�H����)�=[$r�S��.8�j%$Q���3�I)�0LF1��,[�V	6J�E�f� ����h\�<�74󱜥e�3r�lt�4BM
�I�4k�aNP�d~��>��<�s?>���S�1�DW "Y�Ï?�-��K��#�d5s
���
�S�����T�3�f�(n�oF�G~��g��~˷�ޏv�Q~��6���W]/8���5�����x�{�60S�rC` �]�w$�xv�.�/��ַ*��W�;{�z��9.� ��O�Z�}L��Q4��k�l+;`J�����~�jV�+V�|FZ�,�d2�c�������t�]89t����u/�qm�oc�S��	�]�����m8<0��}�����`4��a����O<����}�c��>���5h�X���Q�������ګ���=b O�#�q�)	`v�����1C��S�Gv��ezA��S����z>��Z/���߷3_˧,% 1��su+Y�H���r����	�S�ػ�y,Ƚ���׊���z�]����XL���' ��1�Q*\�$p��B���BzƐ.��JE�ü.�߹�Y%�L:������cSe�Ԉ�DS+*e
!qd���p���������/*1���B�Y1�_"���N�Q���*ׅ�^�V�+�g�׾�ͤ�i���fw�e2d�:��K�*��Z�#�y�rr��^���<�̀�N��xU��G��%��X�$re�ł�U��0.A'�2��-[�G�d�;5�r�����Wtc\�'%�9��L�Uk��:��ؠgQ�C���VB��Ƨc�2;�y�餙�����I�Zں��3�VV1�S��(J`� �r�Tv$���ľ}�̿%�6���3"�4���C��>.<���֮��G���3K��"�C,Ԉ��V�7���#�S!�>q�?,k�}��x��/ײ
ˡ��,��bp��,��D�.��ܼ���{�X�+7nAYR]�(�\Q	$�r8��eIv��֋�d=}�؜�ϕ� #�c240<ň�e�Ӓ�V(�"N��-�SL9�0�m��/H��h2�yB a%[ �(O��h�)���y'n���صg/���(�xkG3F�F�z�2,[�����x���W�p=y�I�r�uX�q=y�I\s�U��L���xH6� �1�}�v	��C����iwhHyp��X7�/�Z_�r=dn�đ�X98R�E�,;���U��t�~�HT��e�E��,�-�#�ٗ#�z�q%y�g��������寢��[>GH�
NO��W�z�b��w���t�ZvY�W�V���\�@�E3�0g��/��a�#��B%��/,�Χ��ìd��:[P�̠)���}HO���`��(JE	@�y%��s&`;�?�����x�m�Q�k�������q)���q1��n���BaM�q�΍a��!��{ށ7��u�����ێ���Ajr�#���+�� ��_n�Z)�.�~Q�1�Tk���^�h{N��g�~�u @��c��(.��1���\A2�Y��]�~|�ڱ==�i�hW�G���i8ipmk����%6a���X����܁��N�797�7q
�3�� t_UK�e(z^ł�����2RV��"��)��M	C�0_��J�g`�V��8!�$��
�$�y�z�YXG)����T=�Ib<e1�3��AZ�>�үġX�8��u����+[��J�Z\�F�Y��!�Gfi��b��B1��kW`bhT�톗�$gyG���J	x'&Nk�kŚ��8Ǳ�ҋ163����VXL�sE�ZF��m��mp%|��O��@g�lIjB��ڮ������N�\�b[��$m��:k
�	�p����U+q|Pr����/�\�2=�����f���,BM�%��s�S5/�Y���z�VZ�6�Jc����)�⡠S���7Zί��*��K��b��`F��.�vA2��5ƞ+�h8�5��8�K��v�N�!��8�,���s\.��J�)1�,��������b\�Ĉ�*�$��`TȨ3,��4��Lx!S��\V�MT�}Ŋ"$9�\����dٍ�,?2�|�k_�^�t�6�}~?v<�mm}���"��\�lj�=����7����C����p�ո⚪\׬FJ˖�D�;
���.8�c\�⨘-�����>I٘ܰ��{F�A���/)i��9y_�I3�{PK_ڗ�����S�UzR%Vk�j�Of�p���C��+&{" �d��G5cb��[��.�۷���K�Oc��M葌���O��x߇>��.��8�������J$-����U���_}��74a���㲶8�l$�+6�1-���Ĥ�P��B��9q�l�Ь%�{�'5p�3�^�
�H�tZ�8������b�:E��K�ޅ�/Ə~��NW,_�����ڙԌ�/����Ú��۰V��+W-WB!rP�©�T�z�gI���{IEĂ�h��I,f/��}�����&�\F̨PX�b0�b���{��%�m��W]�\�I����r�>}Z_��<*�w����0���/��g��)�@v|V�KV�ȧ���(PHh��W�h>P���'�:�{��99��փ��1=�qq�3Si����)��AoM�Ĭ�Pɷ�h���)�#����z>��тz�g�4'��a����v�+�����y���J�E}���k��Zc}��o��Ί����`�,Uš�����m��CC3��}\am�86tE��m�nO�ƠD��F�B�SIk*�<��B��������_Z�"ۯaoԗ=sVyv�ء{���M�]a�ܗJ�S͍�i���!u�3��$3��|���.�Jhs��#ӵ"`E�Z-��)��5���D��Su,׮CZ"p�F���`4��Z��.��f�Cj�4��k"$M�����#�Z�Mjۻ:�1G���mزa��F)Ū�r8�5��~��$��N�-�T+�$�8-��	�	�1ٌ91�Qɶ9��D`Ȁb�dN+y�E�T��5U�&''���t*��r4�e�MSh�őBKs� ��T��=(����v�|-Z�s�(
� :��@Y�;����>���������O����&N���IFۯh�m�.ǯ��7���"ז���nTn�8� Q5%'f Ց�ݗJ�!e_�\bśɴ�T�M�{�.�����dωY��}�������e����c�'�r_����bÆ���6�o�����O)�륛6anv�]���,�� �p�0#Q�~�#8�J��̱e�ru�=����U�����q�������ơ�G1>9���N1���O=�S��ǻ�������mƢ�p����#ã��JI�`O����hB�ü8�F��_|Ri8�K�Z�0� �|�@F�d\�D9�� .9.�X����S�oP�����q�8���U^p��jA�ɘ�Ke�@�3�i4��1�y糮<�s���.��ֶNmk�-�m����fQ+���~��n����N����٣k�{���e�89^�\�a����Ɔ��'.�����٣N�s��8�GZ.�eX�T�qB��B���H^�xL�
�"z�$����x<����r�5����	ЪC�g_�ocR:g�i�Mu�J�dȝfU��l���o��֙�(��ޕ_pΩ�yO�%�o{�21Qd7U$�p��!�1D͒M��vq�MW��Ν�m�����O~����4���M�Z���+��Y�t	�J�C,��SVŮ���a���z����+�r�y�h���A{�>�+������2��{<��	!��c�=�A�ͣ?� W�ge�W�׎�~;тB�:fk��t�
��ٙ�"Ԓ�OkK��)Yzru5����Ŋ�f�³��^tIr�Q.q<i��ѻ�˺���Y�$�B�d��EW�2dK�-Ҁhk��-��o�%u1���d{ݘ�^.��eS�A{��$ja�^�z,D,�y�YW��%N,���SS�m�(��\eՠ�	�3�!!E]�zBᄒT����aպ8)�)���݋Ӓ�D䳑�<�Yq���ܿ��}���o�_>�i�R����+�r�z�!=tPu��,���%Y�hnI��e�N�� 9 ���Mnff\���"���}��OZ��y�`����{�Bfs�=K�;�w&~v����ԛ܀A�ө�w����}�#!��[^!νM�]ny�ex����>���7m�'?���DK�
�9����$�e�ő1$�\{�^,��^���Y�T�#-)'�n�(�e �:�Q�|�Z��Nu$��n��r���+�r��(�M8yzQK2��[����7�ds�d/i$�&H�bv@Y�R��4�h��ɉY��C	94���ߴ��Q٪	�M��TQB��8��;_8+#ǒ� �YA�|��`F��<����}����ӄ;����.��G��c>�QřԌN�p/-��Q�JNt�R�l� J���`�$�s&�E��}N�5�S��}W�N94=gM�M9��+�go߰��
U�%+���R��D,�A����;b�~yXec�j�:��)6 4O�&�3��X�@���I8E�Q	�L2��b O��]�q�񲗚D�E'�Q��=�kR��S(^ϞV�-��	�hk[�I�_�a��p�k���,���`;��o܆���r�h)�2̐�S1@EǐmK��}�v��{~=�=�7�u�c널��	hu�g���"�]ϔ�6f�>���������"���%���6+�Z5�}�� 7D�R.�UEX������Ipi�hy}�V�3���E�5Gt�cnf��	�7�t��˦��[��3,�`&_В���(²!5��;xrG�p(�����d�Pf_K5|]	L�ϫ��o~~���b���w �D�-�>)���f��|Ϥ~�!�(S�`D��x����-�T�~��g^���x����]{���T�=����Y�jT֩����:��d#<�������������?��Y:rkV�P��e�_�+�ܦ4���!0�m�ͮT�b�X"��[���&'��m^Ai<�	#�����g�n�ژ9���6_��QA�3��������Dj{�S
JI��kРs������PĤ�w���7�O=���o>�-_�|��:5��u�ݑ�4x����	M�~��!9��`h��d'���hE� !%go����K�y�2<��O�w�S�蒍�45���ݻ�W��$>��߸�[��Y-�<�����^oVZCK��hG53���� �`K�ւ���j�|�V�Nʽ�#75���e�F$`�%�;���Y���f+��)*#ג/��
W�E��m�z�|�����-E���ciP�7,g�%hr�Yz9mԠ�i���n��?����9�9ߓr��K(�C����	�
���x`���0Z�`nvZ��K�PG��8�\��/*���4ek��]����<�,�lNE��S-`��)U�Sp(i��Pπ����O�a��f;�?�h�ʂ�mŀq�JTU�W����K�8xA�o��o��9��������%�_�����������v�����R�H����^I��*}�7���!���C��޾}7��MML�yE�܇]#�[08˨;�N�"q<��vl���x��i<������Ϥt:�����*����m�?nK{�������ʎ�K$��w�����i�|{�B�S��A�P����
���,��Į�x�O^���G}��#j����l�S��qh�N������+�drbZ���d@ɖ���5��Zn�67��|֌!�W�l��-W���'��&Kh��y˖K���ߪaխ�n���xb�s����ܪ�i�>��☙Q�3�F��"�[�����;&�7Z�vm�Tǣ̔�sӳ�G��M��I�0�<�4���(vc>S��u��э��)%?��Q�����S_Ɵ}����?�=���/c�C��ݲqV�\�&Y�\v^Q����5�02�	�ֵ?&�1ʪ0�xi{(T�8#鰖�cJӘljQ�!DK[���<���2���������},��O�%k���תJw_�fl�&+k<�?}���>\rٕ:JD^�~�pJ�&&Q��lZ2^��>oQ��4�8ц�[��{���/`Ӻ͒�)�U�gf6���lzR��r+td�u����=J�/GK����F���8���>5�iɾ{��#��>%���c�$%x+ʽ���)��L�O�\c17���nL�oi6U
�]=�pcْ�h�@�ɱB��F�3J�k>�n�bx�­�p�3Bk�W|�|�3�����=vTR������4^u�e���k���*�c�,c�u@�_��ک�]W�]f�DqTMy
�`�u�P.�5rO�`�N�{9��}u�D�kz�D���\�٨��z�dU$V��@(H��JFu�&1p�5���3�􅈬�R�uU6�8l]��U�l��g*��w������=W�Q�]99�z����X���Z���{-��<ry{���@��,���ȉ���>��U��~��u��P���%?�����U�$������VL˰�u��J�� �&8mY{��S��?��/��oǤ$}�b;�T��.r�8̄��'rF��%m�U��Ϩ�
�Ln��=<�"턯,ɳ!.j6����N>-H�7-�"���ݥ�\�C�Ⱦ��!'K��`��҃��l���M���G�@���^/T2��i�\�Q��g&S�I��w���)�G�dXdڲf�yo�U���z��?~�� :�-G1��\5��sF��`����+VB2�2f��h�(-U�Ե��!�k#y^��=�X�1���O�*��<���8[��JZ֨�;I6�}7[u�]�!��d��"+y�K��ʥr�s��Dl��I1����O���V������������'pZ���ƸD�1�B�m�<>>���G��x_�Ȑ*)��3f�vtj��4#8���Y*�h\阫n`�QpP���4[�C�#�[3pT��a��숁&�����Ø�Ia|j	r:��ek�ů|�}+����P9��&&��ա���xDRְ/�r�B���wn�wa>���]�aT�����,��(�%(W����r<rHǫ�$Hb�{z:��c:�Bmv��~�[ߒ~-ړ��y�nlCScFF�%;mA��ױ�!�0�:�D�	S��39	�l	V�L"��Q�,��$�`�QP֒��<CMm- �.�w\��U�",f����9`�%���`	x$���y��>�<��0[��;��K-e��Q��w���?��u��䊛������%8���H@5�K.�L��S�.��3=��S@ܕW_������n�c�]���{2���ƶE8�Ր��HTB��؊���gO����%��1�/𱴜� �܂����
U3��`����D�ƂX���Nb8��U�����q��{��!ׯa��NqU������Ue�N=����O�Q!]�{�a���k���_�fN���J���S����]���bש�Q�[ډXSBG�X�PP[��9}�S�4T�Gr����eO���~Mt�a���g��/x��5���!�l�z�lڀ��59�˱��=���/�V���2�9Z� ���<;��.h�&{����)�����-���IdS���H��,g��>�
��Y����F��>,rs���/��'�=	2b�&UA{v�Qq�sXёD�d��۵��i��D�Tdx�(ɶ�oRæ���HM��";b`p;w����)�M�eP�����{����<���	|�����҈��9�<�c/.�չ�ƙ����o���*�i�j�Y�qj_;�j�N���\^���8��J��g�M���~o��j���?�elY�7��e����ߺ'R8�w��F�Z_���hlU��$�8R� �e��yT#�ꗕ|v1��Y��p�(��s��+�Z���Z(j�X��=5$����LZe���"��PS��B�̽�vɖn�x�x�;�${��ɑӸ�K_�l�A�i��F�����{��|T:r6�B;���>%Q�\�a�NO!/�fl�������j������1��;w��������>���yݿ'� ��ׄ�8Nf�v���t���*��[�+��1���/;>�Y>c�����`q�v%���?B�B7�C�떽�	_|���<���3Q��<�W�]��?y�QT�I��8�4������r����nĕ���dؗ*������q�_��~m��M�g�aEZ��C����7��7o�]�>�t1��m�;�}s9	f��cF����Y�����}i�|��{I�Z+��[�ǳl9?a2���'m��pIak@V���j� �#{h�ICJ9^�]̵]s/��]�sе�Q�����)�s9��8<�.ʞ:���z#�UA{��z��%�ɹA�/�T�@�Â�'~�\�썡����]��j'D�H4����� T|Y^9��$f9m� y�ڵ�J����'��V����89<�=��Ӫ�U�[�J#�}+���cVMG�s����aR����ܜV���7o�H	f~d���̦�+�$ �� V��*��Cwk���i�������6�!lD5W�s/���Ǫ�035+7�]"�>����o�&�y^@2�@<�7���2�?~���\�zn�6�89��ɍ���-�
rcΛ������)�iE[�:zF�
ƶ]���bj��rk�W�4`�=�bցZ,��x�-�fR���Z���9�i@4����%F����@��J�b�xa`��6����-�p�ś�j��ش�%ޢ����){�8��kDX��h��:I��!���,��s7��ٛ�x3��m�
�lAi]倒���n��a�u������ Wj�u^��^%�)98u�4���v9XOb�Ġ���|�F�Oҝ�ڑ^�?�����E,�z��E ��Yg�s%�Q~\qv�����d�m�l�lU��'�|J�Q�c���M�E���h�C�&%�
#Jv�\F23%a������%ٰ�3�w�W�{������R�T�j/�E���߳Z�O�q~��iy��LF���t5(�L6��_�Pc�r#�ø��'% �GN����)N�%Ӳ1�?������hr���VV�M����~��+��g�fb]ص�c�r��W*Bz�2������6-����|g���R�9��.>���r8���s>�W��T=�2�v��g�Y���nKq
����:Gn�Q���Fp�ԑ�$/���מ��;�ť{��$���Y	�EM�j��u�r�I��>��D�N�ș�.+mV�U�D< �S9�����0�p[׭U��n~%Mqe��ţ5.�?��YeW���1���}6��5���af�����%@�Z�����6�'rx�Z�����Cׇ�����8��%��e�/���Q��s(eRJ��bٔ��Dy�q��(6��Q,�敾�(l�>̈�C4��3���x�0f�3�6uh��JPq
�lAgI���F
�5e%K�K�
P4��	�xc�?=ji^O��/U6��ԟ/�olJ���V)�7����^�)}1Y
&��G]��5����(L������ރ��%Eos���>;�A������F$C/��$������x2���,�RǢLR���7?�:���&rq���?�Df���+���o�J 6>9��h̺׋cPA�̂΢F�	WҳZݩ8�=���$��R�kF����f}�ge�U˫컉3��Kq�-�a��U8rp/���;1;=����+תl�G?��ZU���՘d��|��{06�Qn�2�xX�L���b/ t����z�56�3z�"y���>H������z���3Aru�d��	,E�Ƽ~���;.�W(��̲�7�O6!"�2/�f����<?�՝���k���q�B���
�(Y!�AαCw�Q�=95��t��sGC�SZ����R��ھn3PRt�a��k A۬��H;1�hy�y��y���Tu�^�U����)�__6��z�5�x��Z�裶���� ����/vK8v��p7��F���ҸE���2�k��ү���9v́W��wAo�ίi��h�ӫ8��a�޽N���A�n*GF�\FC'FP�{>w�$rs3X'�U���7�۴ڂAGq0�	�tOLMI�T���`U�+��JWY�Q���HQt�:ђ/���e���AO�Ф+�C]�Ⴅ~U���! �t�S�Kv�l����� ��U�$���A����U%)n�R)ɞ$��X�\���Ĕ���B��/	�9�lAѶ�Wo��̜�SڑBl�It�w
Z�uܐ⊎����Tj��f.��x�c2e�ZZN�<�������A5Ʃ0�z�D�,����x�ƸWMo��r^@`�}R֐l�V�Aӿ��z ����|�YX��
5�d(�%�g�P��JP�5	!�Ү����+���
�ь��9�Z�Ca� /sd��YLP?���ݭ�:6eb����6���/�Ґh�-�U���ΥL��2,�˺E�lE˯<dV���({��3�p&�qj��:Fy���qt�6�1j���kW����s�Cxٵ��~(��[.��3���v�rX�`㦋��Շ'��G��`4��Fdd��q-�Qx��tݳ���g�'4ш���2�g��U�;�\�ʐ��tŽ�b��5؄��h0�꩞���A�9�Ԏ�*�'_UF�*�k�E��S��n��u+q���dP�6�e�:C�����ɺR3+�i	�Jy���n�2:t�GĨ���ՉT��M�Z�C�w�{�+!���OW+f[~���kdֺ�!��mѷ��1��<g����<� (b��Σ��:S����y���T^;KK�g�J�E�R�;�������[n�+�꿯�j,��������{�g>�:�2rU��H>f����:�[��*u�䐙=�t�\�4A�e0͒�1�*�m����q��Mb���8>8��7byS'FFFPv�b#He�b��*��삜2򁉜F
�"[�(E7��%Ay,n1K�Y[�zՎ$� >˥-�����e/��� �U3[�&t�Z�kF��M���(ʱ$S��;J%#���0cJ-�h"�{@�H��ؕ$KZ�e�w	�9w.OF��pU���O{���"Rs|&���	Ee��5�%�Y�%���W�!q��2豢yڔ��z��uY^vnim��l��[��WT�gy���F��F:���� F	M�U&c��=8��Xڷv*&*�a������P�Q�p~ޙ�q��@ROsgښ����$&f3���Zs��R�U�E־C' ����lF��cz���o�<zG�ZR�㜰ikؚ����d�S���Q#��P@�Fec�94� Gއ�
_�{�����V����"��2�f͢:��$�(j�&'�c�r�Hޱ�p�UW��˷!��K�>�e���nLNL�O��Oзq��B[�J8��*��đ�AC��\+;uz�o����_^S�{��U��/�� 8�}χZ�T�޼���{eҗ2���\�,��k/��s���9��
�4�#�hkƛ�WQy�+�A�=��k���oޅ�����?�y{≉1�t�����k�+�߂������1<>+{�x�bB��%;:��ߕ����5X�8)Hb�{��t����N�7l�2���R?k��rPշA�U^�O�cR��z�o��������,ZK_tI��R��������4�W��u{R�S5�;���֬���)4{J�����imiT��\9��(�Q"!�B�B����JnQ�/E�[�bW[/&��50��C�A���ک ��� ����W)�+74�+���r���f�e�`\O��Tc�܅��]���`�Q_
4��ԣ�( ���,<,�dt�'�y1�,��թ��cl�|�B�"�Y������:&�����ʆ��;�ԢFU�f��77�f�u,eE�zi��u�Q��( ��Ic]]r����%��=7������^��Y�2�ׯ�GD�d�U�!#�9�r�lF�'1�Z.�-p�wjV����嫔����[�����R(*hP'D[k\�t�0z���d���|�ߵk�]�Q����e,>G�Xֽ�k�O�]���$����σ��Ba	��(���r��}|��i �k^�D��������9t����EqD���xz�N�E�\s[SD��C>��?�T�+����~
�h�?��(��($H
�J��
�q�ed��X\/f}CX��X����Ƣj稶[��a�i�u9��S�OH��'i�:��S������ש+o�TyV>�6����z.�+��L�W_�j�p�:=L�:�sp3��]��D^�Qc�W��]K������d�	��������0�T	ڂG��9���ީ��҇]W�6�zֵ��zW�n2g�[��Dp�`Xh���cl�=;>�T*kub�]��t��q �[�r�����U[wSɱ���}	�n$��jX懋V�u��gV��9t����j*����W���}￴��Ul-�2�
z��=b �H��ULF ���k& ���hk�./ϗ�T�|{8�x"���Q��Z�K�e�G�4с<�$LV����ל'/>F^�\0d5�4���	Ș8�v�=�� �^���*J���F�s�9t�rjg�<^|s�����uBHH�H�dډ8��g���!5F� ��R�G�������8E�U�¬���#�VL����5�3@�@$�cY
��8��������5�s�^"|Qwen-�^<�>�m}V�$Bׇ�Z5d2����XV�a�{���K>�Mo�f�a`b$P]E�<�J%�PQ��ʎ���ӉD���yA2�)�d���IN�	p���J.j��Tͬ��Og�^(��9t�α9�)��:t�-Y�Ks��WzTy�H�Ho��̩�/*BY��9W�Y��W�(��+�����hu�e]X[��\������#�>6��{�����$���F�'�N��]{��b͝b����r�J���H�$�>�8�o�u�B�9�3��m�w���`�|Yi���<�U�X���@�����;u;�����<����浅�@�tAQ�{y߄Y�|�+�ȑ�kanR�8�����zD��㓣��jS����A�ٟ��>�S�M������7����;1:;���d�e445IvUP��zn_p�vFk���ώ��	 }��0G�g-�#~Z�f�_����xTm=y�� ����q���؋6ª�R��E�k׮���n*B�N���<%w˟�p�-����J/���|u�y���j�~�/5+\�V�����m�H�����W��1s&s�1�LMh%�ϥ�N8��i�'�l둿g�^P{U֪��F�WV��k�����B��f�\$�y�H뭇�Y^�B%����cZ�l���	�����C��>���rᖏ�v��z��6循npMΞji�
*5d�����XB6ǘ�Y��E��=�[�h�F�E�mnk�tFg��!72�D���"�M���U��^�I�D=x����~�do�D��dy^�R>Q�pk�z5֢.<��Ҷa������j�!�Tu���m%�imm㕩r��>����iH���qcsTDY�yw�H�(Hd����D���}�4���܌dU���*ɉ���PR���e/��q��UNSE9��g�5Պ�b �fݴ�Rg���6ص,�ր�\&��X,��*yq���ZG�1�&?m�g���)h�2ƛ}�`��}j��ݬD�i'������S���P�Q������!q^�^~%6l܈c�=�\�n������M�S CçĨti��2�U4�Q�Ǹ�cR���ln�B6����4�±��`�����z}^5^^ۃ<�ӓS5f,�[X̜h�BIs��������x�����Y,�[uc�D����UG�>4�Yx��g3��J��r�2'�e�Zlٺ�+z153�����O��K�������i=���61�4�6��n#�Te�;���u���.Җ֚��:|gX��ug*� ���+V����gI�D�d����V��hJ����N�p)�k`q���L�;�z*%'��ꉳq���i����a��G՜��՝�����-/3��Z�k�x��{^���Yz�EjD���ڴ��o����d-�Y\�k;9�R-q�|)����kpH�`،J�=;�����@ѫyj{�=hlhCS�	�ӳ��V �4�%̉�k5��{�|?�|!�1VF4y��j�����A����P������U�pT:�k@L�
��Iȴ�jk pA9t�]3��t�X����e��v��rr��w�1�������s��Q��W��7�9"��7Oz�%k���ٖ'�`pc�.V/S���V5�������*�Pn�n��La�e(�@ld<�,k�f�'���r""co��g��7��r��/�t�̌��w�w�}�!j�FQߙ:󣴟1��9U�`���
���|"r�M�������6��X̫�$lW3ߧ�z�������f��L�$�ᰮ�a,���=N��2�Y�����zYp�T*E�@��	1!��Up��lmI-bzAS��^����|}� ©�n&d*���4�n)��U��qSKGj?�!3�L1/�ǐo	�h�{v�["�f�i����t�xt�a` o�met}\U� �ɨ�����C�#�����`��d���E4�j����'&r��1�dO�m'�������ſ�)��3U�����LϤ���ͯk�ّ���oˏ��� �[]�����ŗ�ht��6	2��y�����d�9~���Z{���o ���:q���È ���P�D��{�w�4V��!��9 ��+Y����7�uB��8�Y$��WƜ���^�i[�HQ���)Re���x��[�F��zΪH���k������*s�Y�6Z�o���Q�JuEZ�5��t4�ڵU�kv��d��i_�g3�(��1��5�?��5U���:��Ϡ���'2��A�v�������!9��E�&L����:t_z�>��D�t�&`'�w#`�sP�����D�`�ʜ3�a	�g[?v���~D�(�Ͽ��&t
X��"�0�`����O� =��:��!�>4:��@j����ڀ���?e$d!�o�����!����)�1�ġ��j��|$Jv�pg�D@`�8fŊ�<��3d���EVˉ�wl>A���͠Kp 7�����p��5��k6v,��%�ME��H#Y���3D}�;ӏ��RZ��w��Rc�5athS��#��b�QH�]��([�mh�	�1��"4O�N!F��jj�2i�fggd��r ���v2cZo�s���:z�'I�M�H�׎z�C')�(D�z��Sג΄�+рDE�O'.����sl��5���@���{���i,AԀ6#�7z�s�{���d��Ӹ�}Aل5�;P�6��2�LT��Пy�F%=���ڥ�%�l̀:{\zs���ؙ��z"U�(\5X���F=	G�F�)3�r��^l���K�}��R���_���w��xᢼzmY�<Kv6��Uq����dw�*����k���f�q �x@�2
,��I1j����}���7,c`@����'��m{0�ɸ��|��kS�7`QB�岎��!8�����٠6E�>��>�OFұ���q�K �X���c��>���Vj�k�f�f����ٴ�_�x��g���(�:��81�\��?��?�������m=����ɩ3w������I,;&w����c��_;?b�hi����Y1}h��%Dv��$L$�W�Nf��{zM�� ����{���uG��  ��No}�]K�\j�m���r�ͦ�;�^ϔ�댷�ᢹ�+a�lL�)�2�9����;.*��У�|?��q��A�Q�	'^suFo�,+��(0��X:��S�
,)��#��	d	�ECs���~
�)C��T�tiI)�z	پ rf�uz�!�]�`�B�A�1>#��!0��7�Aw���4飃��������U9�K%�j�6S���Y_r&��y�jc��ǡ E��I/��|�!�bl�B�z���Lz��N� ��Gz�X:`t�L2�)�&RuM�8]���!. � �.�I1�g�kw�2�p��/Ms�IR��객�]���s��>�$��#T��Q��I��lm(M,,.IJ�ӄ �;w�%A��K��M*ҭ�u.6�f�AH�̀DcKhBR��1 �BQ����F��j�0����6.�?��X���̍:F���s�Bw2�|�LD�n��u�bT)�#��r�Шivz#3�Zυ�Mµ��0��A"|:Y��^mSȳ����t�;rL��7���T����%���NԸ�����'�}��M�K�(J��d��]q�b�rɚ��U�fD���A �\���f����H�03#���v��dD����Q?��bRTX�	���q��ǧQRc�A3p2�ڄKdA�#D³�(n�˵�]����I`�R ���_���ujʑV͕��)3r��5y��r��+���$�%���+��/M���L�ȓO=-՚��|��T��ړR{�y3P��'��w�?��d7^����۶DY������c̀�̣=�4�#�5bgJ����m_�k�� 2�~ ��	d��2�0�؞	fDn���_ ���ޏ�C�>��1֔ܴD�8�#�&(�������؟���C�>�����a����Āe�s<�+��l@��$i �a��D ��ed
���l`%�e�Ũ�@ȅi1���]PB�T��lk�K����}.,�X��:܋AB�i�}t9�}̀~c7!�]b�w��<�PQA,�Υ�/3S���v�Y��g��&��'z��m��::(]�[����G 0`AA�O�k� ���GȾe�b
B���PeUp�1f�b@�~$�<jLӿ���6gZ=pԴ�*'�ҁ���Y�ͧ{<+k�W�б�6j�� ylK5i��>��x�=�iD������������α��eggG��\c;=]&��é)��M�lfkmM�Kc��gȤ�0���#�<1-*3�yr!W���@p����؈�o�ރt�nF7!���|[��G�dO} i��бz2�8������u\��ƒ�$�	�L���#)a���fL�ԢUh���T����e��a�r�|���I#ǌd4�}�dژ���b�,k��\^ߑ˫ۦ�&W��=&�>�����}��D�ԜL�ΰ޿��FY�"BZ�\�i�ʩ���H'��\�r 3#!B���-��D� &Te�l�ꑂ'���ܨ?�W����i���o/W`�X�����yX	̚�:Mb���|�ԃYCօ���`��Ey�[��  ��IDAT_�{�]ff�U���ȩ;�ĉS�lt$�r��>�9��/eckO^�xE^|uE�_.]���O*�	kH:��U{�����5*��uB}��f� �f֌�u�쁨��>}�O��B-�]_D�)��QhH>#�� ��N]�5CKh�ۑ�:��9]�3 >�]1���2��������l^��f����l�3N�D{���Ε��ۯ��n�y���x)� 7�/9'��+꫘�O��~@��Z��a�'p@UV�ы�~�0��ɤ�	�#�  @�c������{*/�J"�FV��R�o3�E���]�\P2�?�0ُ}�񈀦�Y�Ө��rS���/V
+�a������KK�W��H}Cz`��ƻ�T4��t�Rܔ���?U�o�J��T��kSKߥ�&af�F�� i
�:�zkÎ:~�d0zO#�x�`HPHV��Μ�֫�w�����ԩ\:ͩ>�$�rMY�/K����U9s�y�WT�/q��U���)w�f#�Q7M2L��R�[�.`l�^��¼�+%���  	�^,A�$�F��/�ߛk˜5WGc�2�ٕ\�?���f_.�鉙S��+��e?���@R�!��Z�v�[�0��6����H�iv��4F�0h]	�����h�؉c��F=_N��!�IO7�^�G�R���ݜF<#*D\G���mY�"��K�(J�䌸��ݶ����s)����4���6[�5�FZ~w��������*5�1U��f�0����I+��j�a(*�x��s�L`��0`��_45ڮ)`�PH�_�XG����8Uۊe"!So��A�w�)w���3Qe�G��2&R�z� "���q�� ��l�x�|�IL��3��3Ǘ���F}O��t���]u�w:"���ٖ�+�?mn^���e����?���v�!ϿrQ��:G���;�p`��I7l��׾��)�؝������,
0��a�-��0�x�s��I�sP�-�P�A��e�{��<t�����W��� ����O���``#쨃�^^����%���9�M�*��Ӄ r��s~��5�d�P�5��G��zs�E���x�?q�L�Ƙ�a.aJ�=�p�A �W�L��2�9���Z�$W����I|f?��M�]L7�z�C�1�@1�����u�F�!@�ݵ���0B�N7JSȍ�a�
�ު�4
L��Y�3���︍���O<-�ʬn\Sb�Cb��D�|� �{��[� `�:�h2WMlh`h[�J�y�z}��W�{27[��'��8�g�;/�rFMcI�SI����s����$P��4�Ԁ��}H��:*_��/ʥ+k�wiU��_ֵ8�Q�'��{¾R�s��:� 
��1�\���*�X�N'c�<:���MD��Tf�FQ��J���,kׯ����F��AS�/�d����J��#-�z��O�V�$����Uˬ�Xޤ45R/OͲ��[\�K��O�|��T��<�:�Cy��D�����/���M��W��㟰n�'�JFJQ=�>���n�dsyN�C�H9\&����^T���>��;e��%����#��'�D�*�RqF��H;5IUX�nm��Ӫ`���0�p��U�F��J��v�q��"EB�$&Áa-X���Xv8`Ȭ����f��܈8���1�T��%��L&�X�(Kpԣ�3^�a��+mSX�1��^�6�5EJLi#�\�A
�;u��4�1IO�K��Ɠ/��\7�+�G��T��R*ecs���s3��KW)[Wk9v�G�+s2�P&������Y�{��n������(p���	,���t�� 
��K沒)��gӹ�cӲ��5���g�7�×�c]G�M*z�������)�A�k{�����=л��ˈ��@�݋R�ߍ#�9�>����t�}V6*�z��B��  V�:U�C�.�%��:�z�u�'Q6�1V�r̰�16q)���*L8��SD��	��}��}�w��j�s�]0�=s͆	Ή0���k��|V(��)�߄��bn��G���ѹ��!
��F�阜<qD~���ВHmOT:��Iefe2"9�>� y��q�ư��YW1Y9��<�愑L�p���NS��(n�e��}|����)[�"���?��+M���)�1�C�6�>�B�Dz���Q�t���\]�[��"���\�_���L����)9{򴜿pY������0�0m^� V�D؆1���z�i���63;E$3��j(.]��H���DN����h@#��'��uY�xA=���Kj��r��y��K�<��2bZ]b�ȴ��#���Y��el������ ��$��P=g�MSق#�,�F�zuX4�_.��<���|�Cr���i4��o�+W�-_��פ8�Q%j2H�wP�w�l%��L�c�\�5�8-i�>�ӧOJ]����N9}��V���G�W/^&_A*���@ߛ,���y���Kț����l�vX'�� ��O�-�N��w��^�/��Ir�&�UBf���9�;u�]3�i�a1Y�g���Z�Z1|�1� |?@g� 晡7������%8JD�u�)I3��A&�Ƅ*�aO��D�N3�2�:�����L[@�#d~������#�D#t2)i�]��,����TT�}���:�~*/�w��M��&R(M�^����rH�H�X'���Q,��K@�T��� � z<��o�� �Z�D�+���E� H:&�]>_�^���n*��#�-��[&!�VSz�@����tܹ�K"��s�[�����o��}������\�r]����H>+�uA웎��"����G
�'l!&��>��F�`�{���L�ˁ�ʥ!�á��k4�ч��4� ���� t�`���%X~$)V2e���΁��Q�@u�z�2��S�N��ȣ�r�)� ��;��Ħ��{�ClC���l>Y��fa��Q�m�����b�z}���ӷH0@M:1�0��K@\_���œR."�����G.\\6F�3^�ı��1�a���9A͖�)����C=6��ĵ���!�\�ㅚ��@DB@�(��JY���r�=��}K�"x�A��?���/���^�O`����Cd[��E��#�����C�ӳ���Ү���Ԣ|��Rɗ���p�5�a/0s���({fz"�h�@�{��˚���=�F�T�ht���{�\���iĸ+U��NU���mJL���JZF����^���vIv��נR�G�� �>[�a����Q.�k�mO~��d��5�-�Z�Ψ7�Sc��$E5���#��9
S��:�F��������������u4T&�'�,�VC��&4҅{�L�<�U�tE��j�3�1e��b,��`V.2�\߸.�uV�ſ�i)��@	8�����%��]�԰d$+�SѕT~�QU<����-�2�S��zҧQ�>��m��"i��+V۠�p��t^�Ty�"���5�{] ��	��o93,(7 +���� ��M����	���u�&j��i �G�@,-�#g�Ր�G���?&@qj����$���(��z�h�ܮ�]�,_�c'����*>r%C�䑤P��������ӯF�KpҠg��ǏOsx�\�QQ� _6�:!Em�DyK���쒲���0 �T�S��q'��L����$0����������*�8�$��������L6">Ɛ#%�UkS��b�T�[��'f��䩋�seS*������Tf�5��,�p��xN^%\Gd�\ut��;���~J��}o�������?��� ��@�Q�9��5�$������1�kcx|����,�>�4:�����4Em���8�4ԨI�3��� ��L*�"�%�_�^���3 !����w8��9�|��3����Sߏ9�� �:Ѓ~GfTנ<���2g���Pu��=}��zu�'RYëOG*a��Bb�hߋ��k2<n���������E̖@�: #�9@��T����j� ��
���0#��P��bY�����c���o9#��{�䷟Q�7����G�rʁs±�h9��8&�w�ߔ��FC�'�!-l�� �z=v?3���,k��v,5:���dґ�_�����j@E��IQ���ƕuG�� C��B�#�	#�Ȫ�ۤ�y��s��'���#��c/��NC7�#[��;�H<�	�=bz��q��O��� �E�/dM�y�!;�;�`RRBO�^�Ç�g��K����˨��ޓ[5Z���y�p�EY~��T�q�m�Aw�2S,I�Z��mHQ���d�h��"�So�6�kU�%�,����;^O>��{���c�Y��W�;�x?̳/��X�,/\ؒ��>_1@:8*�TR�\�.���ߗ�����׮ɋ/^��:�W��ĉ�����U�Ɔ,m@������:[ ��8��=�qL�3�cU/ȸ�F��IFث�Mu܊����W��KKFU��Ϫqo�@�snf^n={Z֮^b�R�S�ӏ�C��^�ҫT*�a�����?6t��L�ivը��~ ��m�\��Ccl]w�����5�+����&%-�gubԀf�xhı=(2U����4�u)�BnﮱV�[[���9u�L�$��wV���ls��C�"i�>[t`�z���/�%��3���A��|��G-5��H�9��7�NsW|�C*B��̤ԉl�!� �{}5$i��Y����Q���/A�&	,݄�0�\�B�=ᙀ��?n�y��85��E�%@wҹꈲN=�Q������46l}��8Ϋ��nw�l��lt�ah���eoĞz�@7E< .�L�:�)�|Nv6��Mw}X�/�`@No����dCY蘡F��F/�ue���]��HvJ�EΠ��rL,�[��t1�*�I�����D4�V�N֜�"��@7�����ZA_�޻�`H�i�t �iC�δ����@<*66C2�Y�h5����8i4PMKF�tS�0�c��F�����!2p:���l�')Y\� ��Y�B&��T�8������5���B6L��l�}�ؑu�����O7�"n*�^`Fi��8����h�B�5�VO?�a$�����¹�Da/_[���CݘԲ�,�s�I=بL�!Y�f!b�L\#�xxT�ِ��x�N���c�w�(>��:
��4���������_���F�]��Ԅ��`��v�d`	7@��[�������3_�p��}������)�J�Qc�Q{<���6�9��E�0�H�

��]�4T)��_H=������ʔF;9�h���n^�i]�C�G�*�em�L�
���q���~J��oPH��<u�8��0��د]�l;Ƭ�ƙz5k��8T1���r��	y��w�����r��a�N��U����ʵͺ\��;��L�c�i5zz��֣Oʺ:|��*�BI�mZ�ǎ�\�P�Z��H��dB:��`G���w�5����!#t2{i$�P����lUa��Fo|�C*;�A���Á*W=��E����(�����ǜf(荍)�����=UJ����1+�%�2����Q;�GTf��@?���f�{�o�B"��kO�S�hY8�euN�SY�8X*.��O�����m���$�41T���F�qC��ړ��
>���tc|c�*ɧU�' ��eo��U��p��;�H~Sҵ��E^OQy��@�����DjTL)�6"}P�]5�I���ڨC`XZ�D18#�>�Lt�S�jh4�?��O�ƺ���u��aG{#K������ WHgi@'�̚1Fl�4�E6���I0i.�e��=P�Wg�?������]]��K�	�LZ��H�Y�A4r��#�����O���	��=�!�$��d2�RJF�L)��A*����?��s�ַ�/���Ge��9Iʐ�GA�{%��^O�{D6�q�N"�Z,��k#u�F�0�ͽm���|V�"b�fGRj���=I��8x$A���' �X�ڤ�ƾD)	�Vh3��&���r&ɨ���ڍ��:�� ��F����UNB*`7R���%�3	�b�u���P&W��Dt7��L�@��4(��E���� Ȋk� sw�0;l�m��l����?3A,�4�A��O���ʠg����0R�;aZ#4�l��?Mi� �t6Z�<��E�tC'Ab����ܤἶ�����E*X��|U~�;�!T�9�6�EHy��t�{��EYѫd�'ƈugp��D��e���L����T����s�h�d8�.��p�vo:Bu��A��B�/���P�z��C��������d�y9��$Nҕ��e�K��Dpã왬�j�U�duS�Q�ט����7\J}�ݔ��o�uu��PJ�7�zoU&�s����NA��&��F}p:��F�������� ���Up���ɳiA�'��Vr��s$��u���Ҳ:tD._�,�;{r�{��ڡ���V]�Ԭ����,��=���z<�%������4W�Fƙ�tZ��)p4���V(�R�D؂@g����rE�����徻�cG��׾����]�tqJ"�ʅ��gt2.W.�"G/h�֗��Qgc[��6��ظ���c��q��h�*�4A�.-�˚+��l�nW�M�L�Ө���52���E�;�/_�6te��R��ǔ����%��3����9�Ω���f��Q���JN��Q��Ag�i}dvW/��Q�Ʊ�~V�uҐ�4�MN�::;K����s��][�M����^O�è�er�KPi�f^��q��fK���=0̉�^���Cƈ�k���Q�����H�,H\eiΔcd�����C�>N��E»f�:c��j����y][%��ᾓ���
)����N����цb�:f���m0H�R�=Q٘�v�4��^\*3+7�O��&i�m���P��Sg�#�j�ݺ��oR��3�� `��5Bv���ct��(�j>3���\���e0-b��G���b:2�c����,J#E���i���+�AS�e�����-�Xg��K1��*@?j@�9��k��Ә*�� �:�XNp�����&�ð$�l 2f�]�dR�P��?|�5�}
Gy����5�6?=E�D�U�9�e��Cul�>��s�25��!2
�I����=@B��z���VE��	I{ o��T�5�6D_a�@�F�怈�H�H"f�6��HX�i�{B��4f"��Ģ�!zd73WQe$l	B��k�ݝ0���y��I�?}*N��	,r ����^q���� 0�MH�e3)�.��r��
^�c� .2�ɘ�`�2"�Q�Pp��fy���-�z�#���h[q���iٮoɸ�
)�Jb�!ҟ�'�m�F	���"2XD�vO�XJYW�j{�/|Aצ���95��Ր_�tA.�?�5�����ʞ�;�d_y�%�z��<�8!G���!:�JiC3k�=����{�T����*��� ��G��긨�V�w��c%9��4��GO�:?�V���;����.OL�36��3Tb뒣	�
����(����1�hZ�ƌ��+��Ǟ���=����o�F#�E���?���͟�t�:{�O�X��D�_x�%���4�5��ˆF5-u�p}s3�fn�?R����ٔI/�q�S��$�z|8��Bh7!� x��k�12�=0d<��1��g��e��K{���X.�3�u%�
/P�5q�� �5����:��=#��hFߚzl�k���C#����&�6��F~�q[F����!	�F��$�/²Z�0�r"zM`8���M��i�8��E�N5{�ͱ�qË�b� �5B����M�� Rܨ��@�۵5�\M�6��Ų����~��Re�F{�A�����t鰅Q(���W)�
�g����ݖ��>a��%��e����ʩN�^�7�;����i�G]�ބ���Ef�+�^C\u�8�C7R��qF�|�����3��:�D���+�umOڤN�6f���$2،�*Sވ��ޙV�D�Ρ��wd�q�k&'�G�@G�c��)ؓ�1��<q:зcC�R�mʜ:���,�5vUvיS�kң�H�yG���N:5i�~X�o��1iM-,v�!J
���&���uLdu��E��Ĺ��6�to.����g�W�i׶���9=���?ڝ�^��	��Ub�\�1�I7䧄�i�L"���T�Rk�esk�(�Fz��6��Q���P�ҏ�E|H򁉙��볛�ΙG�'��@�j�UR#� Fx��3��b�4��B0��)��5�J΂� ��n��Pi�!)��|U�j�*Sj�䨮���[�1�-�ia�� �2��B\_S�)2�.�f�;�L8�`<0�˗���[�������:Ou9qdANh�9�dwg�Be��*6�5� 9�|�$����Cr��1���{.���fԛF����d����u;}9��7K�7��k{�pxI:���:�N�|ٸ��r67#͚n�n�5�N���.��V�}�.4�	�)9��	B��Q};���A"��[$��DF�^[S�%-���Ajd�ȫ��˺F�KǊO�K ��^M����et���,��d��v2jˡ�ò����:�b<�y�ߝh
*���MF�4�A;�O��M�<�J��@^�0![���^_>��l�_%��X��l��ft�]��Ⳬ��T:���AGf�z���h�X�urFj�rᤪS�R�If�c�Nn��YFv,`:���CV��dql��>
� ���њ�>���yL�{Ɲ ���s�qv$b�t@-�4�u'j̆*R'���%@�:V�ᥤ��&��#3,���̠d�1�*�����k�ҩ�խE 3��Q�>�\2��y�bu�P��	�K���6[R��������0�Q�RխVW�_"��G�
`:����J�����"����k�\0�-��:Z6N"Έ�sE�0�� H�� �K']������,#a�D�"J0t~�s����
q�q��? �42���l��ܒ��!7L�Î�e��M�Đ�s�o'���M�z<�[�:2!�0"�C��]�g�����F�q�x����U\��z�l՚�Y�gC�"pX��5�&��X�Ȏ�.���L�>��|���ʠ���޽�7l�D��c��"�\Iz�0@�8@`F���F�%ӳSf3,�N�{���#�W�����ג[N/��̂\��%���H�W��U�� ���)p]�tI�6�j�gę����m
I#�!�J#: �A�Y�.�b;a-���-U�Mɨ0g�	�PՋ�K�M�'�G�D\�����E �r���.�K2�!5�$�U��)^-=!��Hq"l�P���M�4wt|���'��>�Q*��::�RV.��F��t|������r����a*z���(Sv>4��-2J;v��loo�9��!qn�������g�=�y��r�Yyꩧdf��rO�.I[��j_���e�Tic�����`I$�/r�YZ�2qD� :ZO�
m��af܇��?�"fd(L������7P�H��:5�L�ཱུ�-U��]��EY(��O�0���+R�8�0�ıw�2�P�hb[�w�6���|D�R.�[�L�õi�T9g�R�^0����b�س�(_���>��:�萳��m�033c�~�RÈ�b0��8|?�;��YL�{�V�!��?6����?J�N����:��U�ߐ}�����|[*�69í>WC�"$l�~�=.��4��@/~.����X�p�l�CK\1_�)u��h\0�#�+SEF���7a���cT�#��8�]���%[����z@F˥J���e��(r�c�WW�G����2��Fgi�$�v�-X�,��) �!�{��Q:È�s�$�uc�X=� ��5�Nl>�[LE���q�x�}�M=�+2	h���R}9�O�M����2���(S�:�E25�>,��XH�ۤ�L�lq������3�u_��y��Ŧ�ù��h��IMԹ���0#=O�-2ߴ�DI̩��܁N�=]��r�2�b���5֩�U��V�ۏ�@�nݑ:��P}��:���6(��s���t�7 �����y��Q;�k��7�A��������#0��g������D]�RE�T���G	�K�!�V��H��P�qSW�>$?��Zff���?��<��_Gg���r�ߓ��U�&����n��8u��|�	�h3�
��v�����Q�����r��	�sr���a<��e��V�ɨm��Qk�RT�;��R頶竁tS�4�Y݈j�@�	��*�ZM�`.%�rVϭ�"nӷ=�\\���� �8>R��L$Έ��8�i_�r�6v�]]��'[Uy��G���ޠ�J�
�iD;� S�`���U����� �3�~�Q_����#[3����a����˓��}��4ꟕյm�M�Ta�F�^��N4�	b�!�����ē*#��Be��JDg@H�Q$H�3�26��ov(����4b�2���P�/�2��-��Q��DN����g)�V}O*Ŵ�չ����ײr�%*���U���Q2�I��Ge],1(��ޮ���<=��G�~��D�5�3sgt�j�cB=`4���5�f��j��H�88��B���w�M`S��`��<��ఝ�-kdh�]�9Y}�0:��8����c�S �q�=q���n0�����0���ؑ��Lk�D6P�H_����粥��j+vl�I�z,�TtM�հ��{��f^�c�5�q6�n�08�(	�����d84���aH�������I�Cnp��J:��	Q�B�-K�\����� �r<=D�d���r�l�} �h$�hĢ��^y��L�A0�P�j�LJe"��q�,7`�!�4��VW��/<7���"���m��&��:VW��a�KbGG���te�CaZ������!�ͽ���QQ�f�O�uU1��X�}�������-��	F�-�C���F]	�t֌�ǑmA�v�*w�y�r��۫�T��������{�vQ?Gf����5QK�X���E��'MV� ���ܝ��5������o:����1�!�5 5�J��T�!;�P��( ��=�qZk3���G��\�P�A¤�����SC�����5��G�G��4뛒�����i��T(:�\��G�I��6��X{o$��/p��U2H1t5���3�:�\.���i��ڄ��fnN�)����ьq1�*R�xA8a(r���lnk��Q�VK�cK�.��YcX�aWsʹ��I��c:��n�eq*�����9@�8�.n.�fe�-���e�ޕ�?��5�f�\����
��n��G1�1b����m����e���u�����g������F������k����`ڟ�Q��C4�]J���[�K-I��������M������j�/�o������[J\*?�(�Hȳ�;>SϠpȑd��%�
|䙩x�����v� Y5���Se���}ղ�xA.��@ ���|��mm��2ylooq��3 ����� ��3=�`��3-l"��g�ǟ�g�n���ڥ4Z�tڌ�&i���
��X�a�x��� �^8G�P���<�C,�Y?37�]�l
΋�u�����g���:ɤ�_!.�n_��
�@���X���=�j�PC߭��X琙ͭ��@8��`v~��G?9j�p���7�H���^���a?�9(�ZpU}]�<Z\5���ga`|�#]��0���p�8܇k��	��fB�
�+wZ�#*DmE�lc/�{��y��429	��F
	�%z�rD�榛��>K���?��{~�٠>���-��w��N9#W�]6�����{F]��#'O���-��rY� �-����`��<���y/8���:e&d�Q���:ww�ȿ��d�~�=�5.���%����͍��h&���U}&5}��1�>��5o��� a���ܳж�jRg��L1�z�G�{|eu=��t{��7QǢU����/�,2�yu�Ǿk����}O�g9_���T���@�b��*I��5�(�Em �lx�Yt�1ӎ����ް���3+~���̚��,9n*�n٩��h�p`�X0�~��Y� h&���;��Lpv<#�0��	���#�5�2Nޗ�����ʑ�q��Q�d���*�J!-�D�`((D�@@�Q;/I��
O�?��Bꎆ\�>�Q��@�-�O��oR�z����C�P'���.R9�μ��x��iX ��*���;����_{\6v�ҡY��2��8���v��I`���K/:0s��,LƆ��}�qß�	�[�y�μ](ȡ���E�&��C�P:�=y��o�ߔR1��7Z���f�p�s�ؤ�W_���h�����������R?w��l1��P* )Rt�z�<e�JܫU���0���M}Bn��#G�Q`X�)����axH��1,n��8�Q��m� R��aM8����=�Cߗݨ�筧O��e5����S=�OTq�e���5��*kT�bi��\��ı�4(�N1t�9�9�q�W�\�#"4�55�[ja\�T�<�z�`�
�ŕ�Kjb���F/$Y���:�a]��!53�L�Q�	�zG*o���.�����HA�6�h1��d�? Jx.ulU�݁i�ZWC�>��h�T�+�@��������`c���K]�)�#��p_�cʚO:tZ@�:*[���t1��r��8��tZ�7�zv���zL��X��]Ү{�:(C�v�׮�m�����h�K "�Z'���0�qk��k$�E3�v��x\d �N�jc@K��Q� �&���%fېuA���FQ�7�����糰���N�Y�t6'���.�I�E�N-uH����Ⱦ$��s�5�N�c����3]�Ç�Y&�"2;�Z]�7�%����5]g=��ܴZ���h�����,���߮� 8k���5IRum��1�w�	�E:�C?�#���O��~U�x��1��	��15=�{F��`�����6��#�5DK[�%Pץ�&h�@Yp��i	�>��ſ589��SM��K|r�F4��?��'���/���fB'c����39�} ���	A4D�9U�_}����s�_�ܯE�
p7\��o��x�!�qӲ�:����?�n����}(���Ezz,��>,�}Ǜ�P?/�?���q�(��7��9t�t�Uy�/ɝw�%W�^�ӧnQKH�z]f��u�^�.�|R���q�v�~�J�u���MĤ	]f3bQ�<v*(�O���
��R�$�1����~��_x�\��T��0%}�?�S��^�o?�|��F/F�2=#ǎ�y�H׮�<s�V����n3���f2�n�J�(�K/������~PN�>-�h����F)��ɕ��\�v%=��w[��g��N��44�f�)�uɜ�~�Р�F�:n6��N�L��;����2ش>�ǉA�2ˈ�߯�E4��aЋ	�$P�%5^���->@�OĴVv�]��nm� %�{���p= wB�YSk>1�F��eA�~�gWG&iR�95�9B�)kgKwԐ�W�� �=M��&�[`�`{z�q��m��Q>��� ���[Ά<A^��+eR��⍁�m$�2�r�ja<�GJ\e�P���v�0i��N�̍Y5��:)pPȰf�ЀiX�J�I}.��M ^E��r��!7��Y��IT5�� �h�,��D����A�A���U������ӹG;�ʐ��9���99E� ���hԢӁ����e��j��LN��d?2Y���:�we��am�./��l5�T�5��0;�@�H8a��ׅ=���^�����Y3s'�k�H�V^�d��9��5�0���5{{5f$2�4�:`��P(eI���Q�z������d�L	�p8�*��323�<>��f�M�?i�1LE�#�X ���N�I�,���`���+�sD1JA����.�-ctJ4�a�jdBI��$9 ��;x��
�t�Fҙ����U)}s�,Y�\d�}�n�N�b��_����!$�� ���z*"�1�h ��ه�=ֳ��S�T�z�Wu���(�4�IK���
h!G��1�����[������zC�U�8}ÙnR�&�k�O����pq�,ǖf�=��y�pj�k�R����q�̔�Ȼ��=���+�M���o��}�sr�Ē*ݘ	���FP�_�����X��L�aB� ����$D��A�Mc��R�B:	Q����z��h }���m�Ǐ�$Rqw�u��@��=��
�ԇ4J�|�U��1c=�����知a��{�N�P��f7�iuA��dD�0l�fx�Kz?�k�p�<��E�M����[���:	�ܜ��s���P���AJ=f���m�X� �n�$��}z� ޚ [b��U!W&�#1��4	,`��G����յuH�C�2AFQ�Qͦr�D��s?'8C��h�9��5}��y5��k�b6���"f�c3C���D����K4~0��0��=w����&չmOv�) e�,�����N3M?@�F4��7��^+�cp|.��BcC������ٖ-�B�sA�c�,,�˽��K'S��{N���M�a��y�󔣪�=ZC����7@�%P϶�
�Q�vz~Ȃ�'���kQ�8���P�s������/B���B�H�8q7Ž�){(9��ŶO������sDYJ�G�Cg�N�ƨ�/}�KWW�� +��������<��wp͑�
KXò�`�k�{���t�|;L�\^�����_���]_��ao��AC;*���㼯_��_������_5�?������-��)�x =�^p���3�����?���,�������9��j�k�L!��ZB�ŭ�{��_�U�nbtp�-�k��_�2y�mH������������=����_�E>��_�`X��:s���o�[:��wkh}�8�*�$8�2��h���	���̀9�3È=a��бÖ�	���ĶNN<>���U΢���(���g<L ��P���CZ���c�������������C�a���>71"4rr#�6�QOJ:��1HF��S�2U�b.fR��F�.�k�F-�_��ۈ<\�~�lg����������Q�q�qrc����
�F��Tt�#�aʣG�d4�Q�倎��kD���0�����
��FUʋq����F&� /1@�Q	��c�+���=�1�u$�[Egk?`�"��I5�d O|�1�_W^�rޑ���*��e���;4JLi@3��^|��,�9�6Rـ�s��ɀ�+)��7�7�FwB�ţ%�g�f
�`g���d3�'���r�5a��'j4܌d5�ed���<�_��6)Ș r�8[�@�i�u��Fk�"HgF��k�l�8}jnZv5
j5�8	��P7g��Q������*�Q[�3�ˉ[�ȓY	c����TV>�я��t�\s��ƵC�����M�� ���}�|�#�b�����<�-Y
���ׯSi�0��I�>�؍�c?��r��Y*�H��E:3�ޓ'Oʳ�?'���'Y."�$0�������x���~� e�D��|��!��7?�H*���^{����|�G>̔8iU���X�>�-6���ߒ�~�����`T
����G~������*|Ԯ	����S������yF|�ot5ڿ��{�~�'#������ŝ$��W/J��g�<5�t�0��ݔ���@���������=q�����V��ɂs�J�?�7��{$d����7��(1 �c��W�Np)>G���i�Rj���y�;�M�d�ei�1q2f4�'�=q�׋g����fˢ:��� �z�'�h��������$��њ�Б����̂q<p: �!`2#���	6����0��z�{���[�@�x��=����ŋl��}�^ ��@���ג�����������z ;���Ʋt�\_�8_������	Ifm8�G���s���I�?����X�Y\����~��2�w�)Cs�V[��^�i�g~�������9n|��m���@:L�Ro
ޑFᓡ
Z,#�L��P�j��΋%M]�ݩ��7�L�Ŷ.� ��ށV��9�W
T5=T'�yL�-
l��fS%�87K$���3����Ӈ�E��`���z�|�A4/R��I���f�T�jZ�̀R����w'$�(���ݮJ�í#��zkպ,,.��%]ɋ;lI��S���7e~n�(�+W����5��nP�ַ���+<#��V5���Rlb( D��� b :���^��c��Jt0� @�p��P)���FS��9�g�R�="�7�dF7/�?�����}�~���1�T&L���_���`|Rl����ڐ�rAΞ:��pU�/O2���شF��Z�<}��hZ���({��6:5NGõ���z���Uj=�]3O�ߩ|.>��qc( E���:=��;ԩz�Fr�T�QJ�)U����8+��b�a�ĺ����g|��7�E9���k��R�1���W�Ա�˒>{F�`N@��w�˒��r�':	�r��ο���v�iT��!  ��
�������[oa;�P��5L��xXt��NV���� z��ˊ�J"�Μ�z>zLn��f�]/�;ԕ�cMrU�'4*[<tX���(d��; �[����gh�i�e�dK�9&��r^="�d�����8����t�R�4?KlM܍4Vפ���"2,s�Â��#�B��rƌ��#��i�q�3��o��k��y�|Q���:s�,Uk����� � ����� �J[����#E�?�x�-d! �E����qg�gb@���jn��#z�al�Y�p�0����l��{�'�M��a��?bFpd>��͌�Xt���SOs��2�èHv?�I�uK�"�M<�����j����:��-�n�t�(\e4�	�c�D�Q�
O���������^���m�P�r�nd�oK���b�e�bm|ֹiS��$'L��`|$����56�!���ԉ�d3��h�P�2Q����>�l^�w?)]� ��rb@��眽��!�R`|�P�_���>���eTB:kvaQ�kF{�Q���{lk�OCY��B����%��j$k��ז�œ��[��'�3��I*��Ǧ��iL��d�am/��Uq� H>a�?�g�o���و�۰+go?.���A��e:4�gd]��u�i�S�?&�[��9/Z"*�P�0��*�0N!q6�ҡ5wr��U���Z7mm���?��]��b�yn�U�F������W��k�����owe��ɜ*�V�����j�Q`#"K���K)*SF ��}#2;���+w����_��*(�����?�����vi��Y�cL�Y�R��>�k�c�{|��}�� ��rE�f�p8	���?�Lc�*�,�l�(e�ݵ�e9z꘭��X.�4�QtW�.E �z&�m��wЪ���j=���������s�K�#��;r}}��Y�A��ޭ׸�P��ݪ��5�̭�Is|'�%��KE����D����wJ���(8��ňU����Q>��/~I�V֙���Ըv�=C��2�~��r��l��J"y��%��^�}��˷�z�P��'��-������'U��S�7p��%���wy��){7����>%�f=2L��Nx�o�/��_6��0[�'�&}�� @���AȔ�f8�a����G�����̅�]0�6FF��̨�?�N���������&�G�Gt��n��U*eb0���	�%�������E�z��2_��Wd�5
8���a�	Y�;2HX7\J/0Xp�J�ٟ�������=���ق��}���pHj�`�D�ȷ�|��D�����	�՟Q����[�`�I�{S�4� �����<��7u}3Q��(�"{WC�ɘg��q��q:�ĩ��:1p���|�ЄY��-�Y�8�훼0��k�����������&^�B�������������/+ŉn%��v&�ϸ�!�j�@�P�{l���*���ݪL�$���lRt�Jc<`��K/HVU0�GOJ�%�r�0�$����~f���4�LT��ɿ��o�铧�F�_��G�	ŉ�pN�mu}�-+�ȐBn��2;wX��Y�v��܋���W.�&t8�hL�~�6�d1�ꄄ�(����$�P����z��++�3<�Hţ�9R;U�p6��t��uU�C50�2�A�s���#w���M=y���'~�W���ˬA�-U�+�7�!�z�'{��G_�@a�j��{���E�y�ӯ�����R����SN�<-�䟓�U���M*R__�B���"=�ʥX3���YF�)���ئ�?Γ�	0��Զ�A�Fꨡ�������y��E���;�g^VE�i�� ��
�����7#H��U�<U�]Fd��@Zݎ�����s�Ү\~�<ǚ�9(��k��O|�Q.� -m0؋j�_y�U�ԁ{�L���ȓ�}�/��ǟd���H4�#��0S��W�sj�C�<�ښ�~����f�T�p��Q�1@j�
�9Ծ!�iK�5F����%������Kb��J�9a��r
"�.��3�(BKU��3*_QG0���T��I�lD5@����"��J�k�e�P�H�����6f��8'�<�Y��0����e�zC�����/�3H]�38�9��&f3�o�
�,% ��g�g�K��l��"�'yf�*�Ԑ��'�O�哧�~��A��7�It)�S�	��h�ر�E4��q�3&=���a��a���qH)m�t\O'n��ٍ`�	y��W��I��Ϊl\����j��g�l��%m�/�O2��2����Y�
���6ֺ�)�Y�K�U0��� 7�)&i"��Ἳ;5^C��^�Ͽ�����(8I��\h�I�����:	��3�@D��Vh%D�nq~F�\���u���rh(��I�m����9��Ҹ�6ז���m�	bwHW&PP�zcێ�0�@r��|�@�v���0�F�=�5���-��۶�&(U̫���ە�rN��~�|����<� H��6 �C^���_���G��F?4��;Ҩ�Ǜ43�QgFD�I��PC��F}ԥ� ��Ac�;��vӌ=���<?��Ϟ|�'�'�-����9��^x�ɘ*�&{'A^��%b��V�PG����<(�7F��5q���S��l %��pN��CGٗ�*�|*'�3�f�N�z��������u���G; 
�\����������t^gJD	�2���#Oy���ԟ��^P��a.0 �N��`8	� V��Z{��І��?�3-L�v�1�4������x�\����ԶdKk��dv��-u�@6�Uc�nVՀ%��e!s��$2i����̼g �����O��dL�~L������KЅ�6�L��2�a��NI��,c���cf���ˠ��������&ih����WT��_��Ǥ��i�?!G5�� �%�$�"R��N���6#7C���Sވhx�v�d3�0R^壯Nܵ+�dxa���Ɇ� N�f_�;"�V����g�����U�v�#��Yg^�4����U�qQ;�k2_Ʊ�j�TA�}�a�����Ȇ��l���p�/O������ҥ�dJ[�P�NcY%��!S��� 5�� ��Y��Q����D>�����ڈ?eӬ�>�2.�@����1KKBl�Z�1].cVHRc��^�Sgm�����D�)��14ا�6��T��yc�9�%���t/�:p`@��il�9C6�9f��d �?��Ǵqa$*�Fi�I�����f����H&� 9\3C�����7<�+��Ĺx,l}}�T��@ TRg�@7BC��"]��!�(A�+e~C�8o�h�;p(�0{8�pNFHo�J�3�}v�*�X�f�ÿ�=/t>��	�`W��� �[R{糐K�íΰ���8`�c�a`K1�8ktJ�Y�s��6����2�~��c
�`����1ʾ��8fBMpCKZܢ�C仝!�s�'\���i�[���r��;�c?��z���:��V=�}n&�\��|�]�4�	hi��X'���>�:4y��8Ɔ�
S��pp$��.�$8�g`� � �j�
����kv�4=C�����L1�;�~�w ߊ�i�$s�q
g_=S5=2{��d�s�|]�jvJ
S�2���q�Y���iF�P����2�	F��w<���cj'>#�V�C��z�c��p�[�� ;���d������o=ɾspB�
�S�t�o��/�z���7�ȓ	k<qeO�[�'P�`c�4��!#���Ndf6O� O���r���J�<%'�5��9�o���R�r�-&F�r�g�܋d�I\~��ga�H���:�pz�6�+���Կ���4!ԣ�}[ƿ��Y�x�\���u]t*���]S�^a�L��=o�W�ʎ|����Ԭ���N��)�/_��� %��g��R�Dh��,���`"f���<��3� �%ձ��|;��F~�1��)~C�D�.« ��:ց���6m賄�q�t�dF�=��l����ro�=��a��A�j�{�����(%����L��#)��$���\O�2���$7$c`����S�F�x��6��I�^�O�2�=�Fӆ%�Б	�ƴ*s�졣������!��UHv�N��K�Yc�~"�&��7�����uD:�eȀ�Qx��Ģ�F�x��{~�T����R�?�4�B�%�k.��729�ΨAt����Y�7e�Pf�^��[�ސ�'�#@���;�-�bn�2g�����Ӝ߳�}cӯ�vM�[ܰ�����j8�t9L�Diэ�\�!3!�K��T�����.����wP�h����	������=���^K^N3�`>���=,�>o��'����2ͣ8嫗���'��z�ݘ�
jTT�&3�c`�Zd�5�Y9}��,_�,/�{� �(D�q'F"D��Q*�>1H���$*1HL�v�jP�kj`�L�����S���4��Q�^��J_ag�mc�tR2jT��4{���[�la C^JSKz�,�LbB�Ú�k9����Y�>MTH�����qc�JQ���#7v\����)ֈ:=o�֥���H#�P���gtC��i�u���Zc���2��bq?!�Ǵ�a���0
�(d���jT�Iii��4�F���QK��Ug�lQ�
�U��iT�Tul�@�t����x#�c�i��eG��V��amc.oL�z�����Z�NJ.�t���F�a�d �ψ2���}V���?�
8-��~�i`��Ȑ��{�
?w��>H���!�M�� ���P��i;�2$<�[�ChhC*� �b�:ch��:�Aּ��<���Ӑ�iT8 pCcvp��kzh��χ�>�7��������,���ν_N���gz��l΋] ����	.Ra@0I����,J,�UU.�U.�M�d["��e�*Q$RiI�DZ`�b�yw�N�����r���9������%)���.���p�s��=�G��S[*tF�Y��c��ʔR�y�	By�� �cT�ϒ7�ŜUKP6q�lV!�P�W��3������Xā8���4c�������W��m�K�c`�?�wn>�Np������hus�{4bF�J��C�\)*΋��u�ytF�ė��qw��� �>��F���u	�>�:)��8�g�7�A�lU/c�;\K�n���N���Z�ց�@��1J��wU~�0rQi�t~n+�����;�l$��[Y����#G�h�"ǫ�*0ݿ�59P֍
��IO���;r��#ER2˲dy7Q�Y����Y�`��t����G��b�B�֕�����LD/��M���!v']Dp�[�ی��*�*պ*���$F��u�3��������c��Or���%U��9��.![����нls+gm=��G��.7�S h3X�{�X]W%^u��2(#�(�C�T�kR�/X<Z��X�r��t[C)�WlNZþ����{2�]#�I��n�Ė��7
�#������Pi�gn9�x`)�RuA�1|w�g����я}���_��^>i@���W�?櫧���9�c�ա��R��j��Z���ٹY> 8u�vvV�^o���:o����;TA=r����Fز�-ITpY}l��yFV��w�8( �Ekw'�NLM�B�܍ͭ��ͅ3:���䶦�r�;%^�r�L�P���/{�xڑʌB�"P��]Ӻ	3�<ϔa1�#xyN�;�?c�O^y�����PaZ}��=7�s��� ��a�`66�2e���S"`\ܞ���j�~�xh<�0����uY3�1���[�����{@Sa�.��O&�� ��P9�����9�#��N�9�Tf�O����a�<\ۉ/gˌ�B���=79�Q��*���L��v�ӵ9���t���p�3��7p�^�������x�}�&Ix6]�8�c�q�Q�x�᎑��4�9*5#9BS+����US�Q6x��j� ���g��(���	h�ؑ{�l�P跤zt�r�ss`>�1�T9��'Tb�[ �R���������h��.ZaZ őCt�1�%pX�2q��4|���co	�F[)�I�.Zmm٬Uԧ&���������5��$�����~O�nK�gU�N�k/�B��蚬�����C�Q��ZY9��d�@I�*N�mL�ȓQL�H�F��Ԭ���m[��"�5����a��;�sm��*�=`��옔��	ʰߕT�U��t�Ols���8f�b�S�ZE��4\�;0M��X=�]��"�]�:t̀*����q�q����;�|EY[O������_�Bq����O�	�؛�9�U ��PW��
�B��8�[olc���3���'��p
�t޹x���`^A:b�J򳆰Ǻ�W뭷N�GnP�������Y�\��O�^2�
�N4L2�҅CK�YC�z�kTp�pT�<�o��G��ч���'h�P����,m
�J��^�R�PL�nj��:�2T̼��X�q�c����s��$A$��O��� L��kYD������p��m������Dft����Y�+��M���}�QK*�)�a�]���7�R�ǐ;�!r���}���0�A%�B��3��lv/Np�&��J@N��0 0.ȥS3��#��p�� r�?�q���y�_�:OT�\�4��PH��L�(���d�����s����)v�e�F���EcO?��i+a9V�y�s!�G�On3�W4"M3�\��5� ���R_�f�.��ć�ұ���X9�����1�@$M�02z�4�l�B��Y��f2�ps�Ⰹf��}��Ȅ~5[����9�3�d�C��T���ԯ��Y�Z���rQ��K9kJ o
q�y^�d�sҘ���z�έ��KV�b��^����yb�ȵB�0Z�m0� ����s�e%o�{�3�
5�:������u��%�V���o� Kb�A� ��W��Dź���CD,�6oi���n�¬	'p>cܰrKU7��	�U���6*l��F���0�XT$1a|���u�z�]y�λdF=g�yG�Drpeż|
e�6Qv2TA�d�E/� ��ݼ����&F��-�22 !�\W�E�\��>��4�{u7v*���ܼ�?Q��m)��n�So�)��v�gb%��!̈́6������B�S��Ao�����R �W���2T��|=�r���4���}�|��CE��_���Oء��+C�o^#<O荙��c$lg�V�G)Y��J�j��`w9g���[���k�v��!� �e�Y('�=�#޵�`��� 1�Shlqp�(�T1��ypX�j6'�.��{�=�� `2�L%�+�['���c"�OO�J�x"��}��9��-n9�L�d�$?&�4 �~�l��i �\�ad4|f`�0F�A�a,�Ξ���l��j�QJ#�k�Y^����o	�+dd�+��z&2����S��?\R*ۜi���s�~���X	�U���=m���C��ӑl�7M�5�u�V�<���S���9�I�-�rɱy��mXA� �!��8��4<��p@!X��������}��<܉��[VE1[����Mi�V沽�+�KR��;P��JP>�F����Mڮ.0I�Uڒn?��ٲ]�(�>4W�
E�n�M1//V��OZN���@�.l�����r R5�b,�X��Q� g#��)6��0��[R��S��i.����h:��T�$S�/n���PR�F@��*f���}{��6 "-q���|�;��}@Μ�ի7Ore�V����@��Dv{�֌&1�{d9���\bP�bޥ.``��EO�Χ�g{=�F�}�7�dak
����PhY���lo�w!`2/��ߘ������C@|���@���s��UkgO�����Ha�=KRB���
�=Bc��
���U+x�]�U���~��<�� �*Cӌ@�� {/�T�=Z�b�;��������������n���5r
�U*��hHa���F�Ti���I#�c�8���[�悩|Xϰ;�e,�V����iD�y�C�G��c�i8��ErH�K�Jcġ��l�8�T�q��U�1c�I�ivq�5�\�����B�1b���xR��Ã����E�~/"�e��)҄�<i��o���yK�=+��g�M��ʵW��8�]�E���1̓�r�f��ޒAV�K(cb�pM9�3P�n��-�hS#M�d��KJ��Wp�&���ɨi6�O6����[�%�P���憵�n
���Mф����|t��`i�f���[J��^�5�*���E���~�Z����_�o}�9�o�'�B�J06��M	�T���6�,;CY��6 m�+�BE�%
���5�v����iY�."�� V� K&�3��h\�.H�P�V����ۤb�D��Ҍ(�0$r-o1�j�B�����P+?W�_�� "�~&֚N��m81ZF4��.ɛe���\k��|���%����&pvv��w��%KV�:@�U��D[��CVSG�`a�z!�ڱb ᘀ���P�o��v '�1cV�hDz}�lw�7���������7âh��~�ރ��ϭ�P�'�5�)�3����z���k��$̧� ����{���|���v�|�~�A(0#����|��P�Y�._��N������C*8*k^�DGd_�,��s��q�4P,��e��H�0"z��C�J'�]1�9�$Fih|�ahgTE�cݛ� ��g�gRc>�
�J��?b�?�C�����85\C@ ���O�E�x�߻5G�<�3L��\��`q��	�+�r�g�#�i(�A����G\Ȟ[��Y�C��
z���p��:�����;�gJ<����=+_b:yk^���R���|���/��ݡ�B���U�xD��z��p�Aɫ��v��,<$���oX�^� �+�@��\�a�	s�y���P -=��#�M.ދ�����-�N��� ��âX@P�ֹgǕ���C��}����~�{䙯}Y�?!�y�qyꩧL�,iݵ���Tv�.9z����7�wL ��@D����m��_�s���c�Xv�jm���wJz��� �Ͷݗu�t�̬�n��܌����ES��G��5�t��yp��YƑ8B���fk��d�y�3=��g��Gt� +D)O���~����|�:�mpcW��N�� 5Dd`D��u��뚈�w����żE������Ȣ�>����;힅ہ���8f�D���ʄ4��x ��>;�j����=�ה{ཙ�Jf�#�?�!wS�w�9��@�(U{�6�]�@C氻� �@��e��t*
[�A��F���#6��0�$.��N�i"�	��w��T�0>G�"�Q
V�������F�
	%s�'S�ی�s&�ѣ���}R��{�8ǌ�7o���u(�L�G��̇l_"��q��H�W,T�4��=�p�}�9�ug40��8�u*q\�?W�(hq�[+Xgx����;�F�h��u.z)0�¨�[�ճ���3�`6��cpsZ	z]�7�(f���0;��k��RV����TA�����>�%}ܛk�g��?;�o  T�?�LxV�Ap-堉���\3��]�S�kX� N
I�RN)*x㣡��?t����W7��X�IUeY�{�A���d��mt<������f>Ώ\h�Ov0w���vsG�����Wda�*��������r��[2����Vs��0����ӂ-km'̓8ld��[�ǲ	���� �&Ka((ݦs&56hM������������@ ������֚�� �۶���dU��ԛ�$�>]�{��c���@������m5FvUٗ�������W�V��ǎˍ[�r��u9����;w���N��e֚�]-yjd.qTr������(��uF3xg�IC)�Mk5�Ph��d��R7�a�k��Q��l�N߃�FV������ڻj�����6�m�����lU�i����Cr.]aJ�9�%���|�wo�/SH�q���G���#�N)X�<9�V�׼?W�u�?��'��w8�˨zP�P���<���~����w�E��8�,�>�01��<���	 �N�
� ������\po�E�	���p](|�%xTdP��,����8'��6�щ��<`,��k0C\���ü������sڲ��3r�q~4���Pa�>qb������91׸k޻��i���h�H�0J�T�A��z�����g���q�5�P��4�זq��K�8�ɢ�Ly�8t#Dke�)����zB�� �cd-\���آ� X��ݞ����`(�=�gs��tFF��G�Ĭj�S�����_����yN��?�?���z�����vu�i)�G���J$�9t����V��-9qlQ��O��|�c��/mȯ����&�-!��8��wPf���vv�26���4vE뛝s��7j}8q��\-�UZU���:X�i�w�\���=��TnAU�1B�T���?�uB=�}=l�T<+,zz;h`�����/1�5ꎔ ���1*�+ES�C]�͝-Y8� ��Hz�m��zu����47'���-j����X�,7��c�c�{�d�tZgm�۾����O�����9(D ��q�E'H%"DT�G>vȀ_ps���9q�83�|��L�D-��5Z����{�$v9�� � �!�H�f)?��L[(J�!�5��?�&�EWo#.�} �'V�DZS�T]�_2�*U}��[�1��U9�9�k�-JM0v�{B�a���8S����P@���}F!�ô�+�P0R�^7� ǰ��4u5 Sba�?!��+?�{�x�帲�A�B�x�|Di�S���%^ 
M7��N)��g>礢�ر\�af�O�d���
�q@��9s���F�C�`L]����<if6�|�GɉK�}�Y%� ��Ð�EԼa��xc�h���z��s{��'��C�O�<?C�0p~4�!����SX�ESPs�NN:�[{����.pp�q���Բ�"7kk�v�x.<g�&L|��cu��m���>���r��[�60��^��-��u
��N� ��.�)a������O>�OX�����n�g϶��T\�8��u�����j���o�OF�<xom1�POMq$���*�R��������_tN�}O/�׾}�|���g�|c�y�&qD&��X8LR�>�w�2,�aY�,��S`�P�Л�o�CA�:���M���i�ʖ�>��*ەE���c���;��W�^��zȟ�E�G#|Y��j�r�}[̓�Т�^+[�+/?'ǎ��<�$�����벸�b�Y�֬$ncmS����Zb�7;��^��|d#!�V6��4�L���Y��b�A���3G;����������l�f,�O������x�alũS�0�` �^��34Ux!L	�����G/s�}���q��l���`�|�rL�����fp�I�G�ƱS:%���a3��L)P���<��`o�,��>�0���q�c����Xf��0��8�,�m��8�?����@o�a;>�k�[μ~Nz����B�E�¦1P��*#x(w�Ue C���<0}n0�� ���s �9�m���PZxG���P�P�̈��Z���fB�Gv�Q~�ܹ���,���ϱ,�:��s㚸w(���_��!G���3�'Y8��-��~�8y�W�����7����!�'X��5D�;�5����:����b��i����;��p=��P��qO�ÿyLub�`|�H��`Sg��`��"?��˽��+/���ȉ[��ads��QV�8G�n:���@*��*��o�9�~/���������Auh.�?�4���ht����둞��_��E�V1X��Ȭ~EM�4]��b�yl � �^8�1q����/��/�^o⚞V^ 7ظ�SG�2�ŵ;t��1���f�z�Nnv� e���[�;OB�-��H+�<?w�,P,HԚ#���@�?���ޘQ��� �}�LmӪq��ѿ|�j�A
>{x���P�'����~V>�׏��s"�����m4����-�}�pO��J�lFB���(tyb���>�(lqKR�����a-KcN�����uLWF��	��7���6n,T>K�@�G[-�z��oe[L�z�YzpţQN�Tp�*NbW���ؿ�\��+DN��P0���0F�k�1�s�b�=�!v�	�pL��l�CO���1	�c��-��o��Ҁ���SB"Sen{%����\!���Z � (�>~����Q`R��>"C��ѻ�"�_�*uz���?GX���rȔ@���Bc��B�R(>�<czo�_�x1��<�-@��_C��BQ=�M���g�yƼ�#G~�c�=j=��!�g}}MN�8����
�ǵ����e+\s<�8��w�a
��9M�\��aJcE�?x��W��n�}�L�y00J0������q_0<@J�*�}�#z�"-�~��{,]��
�,�q��18���lnp�h�`��k�Q8#���[[���bۏ�.���0��B�xv�υ��y{��D���[��	��L�Ҩ�A��4���}��ὺ*{~��Y~���v�X/�K����:I�� �X{[)��u���6�$�����=ܛ�N]��lK5�˯�.���)��8l�诽yM.��ZRmx�M�X�����秈o�f�qS:Bp��d9L @��@�M�ρ�d U����2r���}U��<Kl�sR�Ù�vX�irt��Ю���z������f�"���!͑NPMe=�gTQ�g��4��r��G���dgS��"?�c?&���>��=2e�/��Q�o%=0`R����Y�����+�\eBjarDC��7T�h`�p�;�9Rнv-Ǟ�O9�C
��7G���*�l8`]��Q?]��;��	(([�P��,D坒(D��%)�dA�>r�[�N\��r)gdC���*��FL�=���ʈwX���-�\�e9��<�DT�T��IUB��y)���tzP���5��ztQ�IflP	C(�C��݌�?�c,��O@��y]zu�����E�9��M&S�K�rx���eA��s���oy|��;Y
Ȝ>�b��a��%�{E�u\������5�}�ԩ,�=�8:�1�̒,�AQ��x�3"�	���7�{��PB���H�~� (K��
�ک[#�)i�8���X��^/� hĂP�4מ��w�R܃���`'z��� � Q�0<�9���� F�<!����(��s��������?��Q.���+no�e��d[��w;�����C���ý����u��M��b�\�U:���0[��ˡ#7�z�	Fol��El�7*�:Q;����'O�K\q>�+$��a|��N\m���+{7���ߩ�%��r�:8Y�`.2F:,��z{�u;����ؚ��|v�kQ͋��4w���E$88�o�����S*�O��lWu�����x�	��\�u��LD�
a��LE���1�Jsa(�e5:�Wߨ�K:���֎\�rK;$׮�<�ͯI�ݑw�'g�]��X9�����SO���s\i�SXH=���xc��s^��X�"˓�5��j(L� (����|��0�Pbg@�k��A���&�S�E#���	�'�|���� �2����d$�!!��T�*K����A�w.�8��|b?ɤg��p�c�'����C���+}����|)�$��u��9i!�Ja�=�GZӦ�p����Ut��Bŉ�Ы��� 
b�m&]��$x �v��{�=*�Q(!O!	M��g�*̩��Ya�J�9|~�ÿ�(A��p^��6���&��!{�3\ׅЏ������{��<���J-da<@��zo��f��1%�׃�&�:T�L�@�`�A9#���5�0Xp?���9��1l̺�m�H	>��$F
Xj��F�9�3y2´"��@����z#���ӹ6����D�J�S��Ч)~Ɣ��8�Z�Z����]Ȁ���&�Ɖ���)Y�p�_~��W���!_[Ppc�T# N�O��H<���W{�g����+:��a~�:օb�����!sH�qѾ�N�W덖ln� �H$�L�LP�� �a��G2So�66��A|�걗Uymln���RU����q<JM�Խ��ڧF�w���¹��$*�Q7軾��x��u�9n���
�g�<�M,r��J�Pq q=ꍭ<���i�Q�w?���_�ƾ��O}��6B0��̚�D�5Ԑ#�0_j���iu'���-]�	��H�Z��ܼl:V�
�b8{ތ4w���0[�~ÿ��/��Q�������E�p�������iтh:��%��Djڰ�綄F�J.�;-su9q�1��@����U�X�R��J��e�������N���	�ܱ�7���Vo =�#c����\[�D;"4Fo���{m�|D�)�X�� ������9��J,�H)W�ܤ���8�Zy]:.ɸ�����A�N�|���X�ј�
v��!�'�da�5����`.ǚ�����/�6烂4���=� g�M�YWN���.HY�{���@h���@�y)�)T�`���:� 5��'���7D�:�3��P�x�����Of
�!y*&�a3�
�P7�axx>��]� �c�� �%���ֵ�s@1cLpN�ډ���G��
�@T;R�0.��cn�7S�^g ��J�����W��Q�a�0₨ ���2ŹP
fs�N�38?0�qm*E�j���[[n��c�ݳ<ӭ�O3M�~I�J/����p6#F$������\q������1���Tr�9hܒp�=��������t��-WMPs�{��.�)��c�]��{>��m{rsv�5b���׽?Z���Գ��-�͎�dT�Ɋ��3�6��ą�?XI�.������4�P�*`K������
g�;�G�YG���H�-&P\Z�`�E ��U��P+¶h R,�2F��
_xL�(���1��u^r�#L�P���<x�1w�>���C���]y�7������~�R��dv~A.^9��T�g�R�3�v�)���A�J��(?˗�3�MA�-)3��@���Fȱ�@vϙ��m���_��k#Y�l���7��3T�\�����Ai�z��\�\��j��Y(��oK=W����zYn� Y�qQ�����w>�	y�#���Vs[~�w?'��:%۷n�f:�םU�搷(�˫0�n��"Sެ	�vw`hx���BU�˱,����Ǿk\~b@�mݬ��WChF������ł~�Ց\�j�����2T��?v!ʙFA�n���������O���>yJ���z��|���X���5I�ĕ��3t�Ci[����S����5`z���s�q������Uì���3k�<r�k�f�a��1��Y�P
�#�����wxd,�J����ʨFY-3��8&��>U+ރD�Jr�R�B��0)>��ҤT6C���c#˱x�=2�1]*�v �p�9�O���������f��M�/�} 7�^�P��N�����8|�4�m{�ӵ.FX������Ҳ�����בw�XBq�Z�͢N�E�=L@᠒Jφ���U�m�~��A�T�
XK�\�a��{������}ꤔ�M��k�eX��!�677t.]�3�;�)��E�#��PQ �B�R�5bp�&)9���n����EY�Y��8��O�Fbp���S�H @�s�0���=b<07�+x�� 0����8a�u��T��ft��2�t/�kU����F:vϸwC�#򥟝�[�s���w�5o�z9�����J�,"�����3�����y�t���.ȭ��K7"��
������Y���8���`�149f/1��#c}�|;�-�2����B���T녪5�(%�*�r[#;L�мd�n �� e�����j^a~���ӆ�Ycqa;�љU�C�N��2��W���l�zRUO���5+;+���vS7��*Т���{U��RQ�h��t��<�K��lmA����5i�Pn�!
�Z����hMQ��w���*� D�K�������ȑ'$��I�C��,J�[1�]8���Q.A;��S�yR����cD��C�p�<��o�cw��~��g�+���K�T�H��;��ݔr<��:,s�tO�vJ�َ<,�~�jƗșSg�Z��ֆT�M�b��B�rtE?s����R��~�ow�f(@hl��ei��f+��~���'�e�!�FKξ��������P罷�b=�W�|xإr"K�L|;�$� H��}NBvy����!�X��4�I�v����2�����^a.<<�Ax��� P�����Q�%]ɇ��#�r;�q/�s,��5B�6�9�X���k�0>��;=QWr�7ń��=x�[}�ֆ��=��H/�1?)k�G���n��'��µ��gX;NB8X.������x	(|(y6�q���"�<�l`������`9ڬ� �9�qm\�5�*x��x��%0��%7���8"/nߥ�~�H���Ü<���-�v¸w<�&8�Q�� c`qK6&>�A '�$�	�3a%~�����(����k�H ���/���&7�G�['��\��s	l>�w<n+��t��!�V�����7�� �C�P�yS����S+5�e��[F4&�v�^ɫ��z��#t�!z;-�r�C��@��� !<��@�Ò-UjE�0)�|U���	�J9L,�$Dk���{#]ܥ��&i�7��FIQYo�4#��2��^z�R�(�3�U-�<���B]�#P~6�<#kP&3+�Jb}��)�T��'���ڱUd��N�k�S��}�*��N�-�Įo17NQ��F�"��{�����PV/�E[*z�G�[�����Ͻ$s���)_Xt5�s��/��/��O�+��+'�WO�K����CG{��R�\='�hK��Ը�(_��l�U�]�������W_3��ٙ9}��\�|���jE.��"��:�^�C]��|��?,���ʗ�&�n\�JA7���#O�W^�󡑂Ͻu�a��GH�-�X�`��?�V�#�!���za�V�+n!I��;-L�</D	bx��J�`b}4� ���`ió�}/�%�	�T�̻���4���o���T88����(�#�����y�}߰�˗�y�� *�Ne��sϙB�w�o�8"���;�{��M�<��9��8�昳�\sl�@٪n����=�p,lm/|���O9`<`�Y�]�C���c��6����Y0?,A�Ƈ�f[O�-qJ���G�+d�M��%�|F�ٰd2̧��;����L&=�>K�9�#<��C�0bD����u��g��p�v�E>��k����}|ڌ�ng�g��E��3S�%����+�6S��?:+9rn�Q c��%u�N�{�q��y�4U"%X�i?[P��x�[�˰3���X	P�q��K��T��lB$'�䡸��q�Z����j�Ή�>�8��"�� �yN��E�����=��q�\� �ȩ��R[��+�8�,p�G�I�>z����<�a�ό���tw<B�yx�Y��ԧ3Ҭ[�g-��/�ܘ�͜N=���Y!��s���-�B��/���X�H�|��_lȻ�W��U����K/�n�#�ϼe�õ���e�\���5y��2_�ͿK>���M��� gwwK��g?#���R)��Va��z�*�Nˌ���e|��{���[���?��S��ٯ��|��U���y�)��
D��!W�V{C��<(��rA6���Lf+%Y��QocM~�s�#�+w�l�.���`�d�z���E�Fm��3#�ݜ)���3��&�O�y�$�t&�:c�G���!��[��VF\�n�`h�J� (zI:ahz}aI�! �3�F��Bz`8�'i
�6�eq��9.%��V_(�0��A֠#�:k|�4^G����	��@q��C��E �)�|�û��Y�5ur�\�����9��p=*c�f.�d4�?x�\���#�,5Vp\�k(�`!� �;tA��J�� "�&�`x>�~�����1\�WF+0�0�����x� 7Ǚʝ��S�ao����՞��l�;Ӎf++���gO�W��w<�W��V
y����ܯЍS,uݳ#���Sʒ*�qU�UKE�5ѐyȲ�%�<}SVo\�s�_�:$x��B<_�S�.ݞ�x�h^��lF����QЍ6X�ʜ9�XH󼁴����v�� �Q�[��V���*�C��Z�m�	L|���ts�n� u�Fz�q߱�a��q�X��{����F�jZx���q?����M�ۈhu�+�d�O��U>�"����r�0�P�mU~[�n�ڢ�Özl35�g�^[�K�ސ+���\�,���$�^y��r�p�n4��W�d;�輹Pܨז���n����o���3:�ݶ�r�Kr\�<�FT�Bة��ޒxؓ3o�,U�O>���6j�օ���\��
�A�s�@�i_�n]�͵jT<,C�~I����	�v�L�h�ڷh	�89_�'��q:�#��<��4Ԉg]�ʡ�y�U�237kq����
^��V�".�D�9Kt�?�w�-�(+yzy�d5�a��f�;��2��F��P-�.�&�~&6!���5l����)؉���ʱ�3@�1�L�}h�w���s�nq> �!��ozy7�'�2i�yH	K���R�@�#l�R7�h~���=(��9��V07��{�2'e0�|�(������\���N>�X��cT&4��P7��#��2��b�(K�²3�	�`�I�K{�S��F���>?��`�lp���V,T�D�2CE���	S��/@�vT�i�ׇ��{;oW�����Y��s� �������P����-�N�����[�]z݁Y�?��-���\�zQ�nݸ,��  �36�b���Yt�Z1&�))��H��؎�J�)h��� �����X:(�s�+�޾iHd ��;-U�=�Dq�B�q�*�ʌT�6V�o����r�En�Y�N�/�b��#؆�F�z�ǔ���V��v��lV��5j���%Q�掣+���>�y�U)�{��uCjey�}wɟ=󜜻�-qy޸`��#im��h'�g��4���Pc��Ӕ��M�Ƴ�q��[�_ԍ��E+آ�+� }��&,�Y���7en~Q��1�ml6��'�����bc��ߔ�뷿 ��cV��}������;^�>qDν���UIG˻z@����dk��ߦ��ob�BWƒ3�0�j$=���8v�r����c�R^c͐�sޑ�a�����Y�L�H.vFYu������&� "�J���5�$��N�|L{�3L�9��$#Cά)'g:���P*"���#u2�IZWd	�k��P&4F�~^#�(C���2���[�}XoMo�Fr٤��gIÉ\�$���ǵ	\A�TXd@cdF`��`��@, �*a� �����du��i��lq|�Ks�$E�Lq�8�0"I���Oc�� �lRCC1�Cb`������p0Hc�T�0���s�cx/���Vo���?�-�dh�ܩĜOW���o+�n��t*�ޮ��7���%U�瓦@M݀����|�&�ޔ/����+WA�
f~�.Uzj��˱��g/��䵳'-_;Q�>I=���ʎz��LT!SU� ُ/y����(�?��_�~�՘�f�G1���7wv����=�PO��Ң;~�*�eK/,��}�? �jCN�9/gu����T9�n��TUcA�S�s*P!|^����G�@>�a��Ȑ�dJ�a�0����V�oMS"c�C�8�a��ސ�9�mG��u�U��FF��w��ϜOԓo�e�PY�[�r㷤�ݖ�{  u���/�s�o~]���k7��g[5E��|H�U��+Wo�=�?,�����zT~�7G����W$�9_���UdW�w�J�� ۫7e��KC�[�}��7���	�ݸ&�jɌ��-��C�G��>�d�:�;d=C.c8�{��Z4��hJ[��	Bh��|B�z�,g3���6}�B��f�/�.�:��J�N�o�Y�([ ����t(;��SW����wqn*p�s�ܫ��(8Yn5���������K!���z�%|�c���&O�鼸��,Ã2t���,���,r�S!�k9 ���|z+h�I�O4uH(4;���U�2
a%z�6��ĉ,�{�7��u��.	q�Jcf&��k���C���I��$�g�=����\t��$�|�����s�_��G�W�Ϛ���-����Ψ-��k��-6��o����cv���W�NF�Z)esǨ63� ��$e�g�chD��o�����s聞��:U�ƾ��;r%2��$x�>�v�w�g��H��B�P���:k��zU-�ֶ)�beƔ�-�ԕ����aꗨ��Ku���2R~��,X�`�9���HonV�}����p�u
)l:Dn=u�uU����qy�{�����x��������*�'��J�нƬa)HgT��_yK����V����Jn��r1�ص�E�o'�]X8�9��4�R�C3�$
hB�f�2�2CE�Q�B����X��183l^5���nȍ�˲�v�Üܼv^f�E�?7�7e�,���̜�Q-֭�\R���¢���؝G���>�J�bU
���@�2�o\ݍ��^�g���_��ߗ��/����l���EF�]��m���;�~}��gU����@�nʫ�}U��^ԡ�n��5���*��ˋzщ^O=Q5�rŜ�w���E8 �Q�a�kr$�����Wz��l�OC��P��B!E+�������f'8E�g%	���mf���XW�=HeO��!e*y�.���0,�?=I晙K��$ʙ9g���d�Z'�����䅿�Yx��s$!��}�f?$����2�I��p_4&a`��d8�<tݰe+_�
�Q�Z��il���7�m�A�|Ή���%[��H��(A������s��k��!kV�L;�����F����z���i�P�����GX�{��gԁ
��4��G�)�Q�n�W5�[:���q4ʙSV*���Y�Y���Q����(��>�)t�|"˻�6r�Ϡ8��QFf\�"���m@ "�#�}��Nef阾�o��Mŕ��#Uȅ�
�z�C��4*r��q�i��PE>�6o��$Z��whiF�pna#<S�r)l�������=w�m��?��~�eW=�?��M�bx�!��9��˦��,#��lK�Y�۷.������rBڽ�*\�y5GPo^yj����+w�9Ƽ&�3h� ^{G�M�;S�«[�BhY^.Fmr�B}���hBR�p;hk�nޒ�lxpI=�vO����,�����o]�g�1�@������PWs}M~�~V�~�a���95�����a���������t�=I�/�lon�����Ɗzo��Õ�����m9zσr��w��J=W��Z�QT�d�%�����w�r��*�����U#�GV��WT7�Ofuy��e��ɸ��<�ם��9����T7�5�|O���fJ�!a�1JÐ^T��7z�,o
��aH�p�<Y�暌3E�s�{�F%C��A\�
K�.�5�NƜ4C���Bd;`����(�_4"p/�<�}�*(v�s�>���)�Z�g�wH{ �E����8{��y��G|��r�֢hjQy�
������-�Yf�b2�/��!�j��_/f�k�>��ԂGa��C�r���w!o�wd>u��I��C�2!��^�X��Bι��1�x�$�|fR钿���N	x�a�rU��e��¹�cj�F #_�шv������c�.?��O�o��祧�V[�5G�i)����(sIi�ı�c����F�؏���;\[�诰z�#��w1�����\����w��H��A�3�B��ZYz�1�P�P��d�
��w��x��\��Y]D�}ƞ���	\|��y8z�in���{�<�R!��E��~�ΎYY̺7=���g,U;-�9X�������ɋ��P]�D�o��oC�A�SχO��E�)I�X͹[���=�����SĮ��^�SťV/jr��gk*�c/�✑Q�����Ū�]u��rIVot�ˆ�P��_�@f���ާ�����K>�eks(���u�ּ~��������6�T�^���F������,�KS)�����tc����U�������93��� b}}��F(_ɍ��<��ou��,�jE֛h�qY�.W�j���q�F}0����#��\�!���R���S�G/�0�eT8!���8�ƅ b3������( �n�]�Bg�{p�'=�=�O]��N��#u�Q�4b��0eh�B�}�z��G�2z���`�u�_e�Ө��&��ŀ<��ؓ@��P~TP�qN�qF<��h�1tM�_�X�B4�" ����*ݞ�a��{�T�8���[���|;˹j����ѐ�sCP�I����R�K�g�b�1!�!��C�xs\�� ��i���z�',�.�0��脧�)�7�>��,����\����~��?�ӿ��h�.��o�w�F ��_����qxd��}o�v
=�┃�����^��(�C@���;�C�f,.A�JM��T67n�H'�v+���U��������ֲ�PQ�kgkU:M���y���%�?�L����¢-m�x@y_4.h�'��s�I.�rM�嗌�5�F�����:w鴼q�E[0��K?u��z����LE�������!t��E��y$�弃�s�ȕ�1O��G<˲�9�9����~�1r�CKW �@���$UA�oɡ�G��5U2zs�z�n�uH+�ci����4�uRd��@�w�e��-�y�Qi�Ʋ��1>te��%@�8ju�>��qO�"9���'� ����s��r}��A�����{Y&)��͞g���5�52���u�J�%C���Q*Cy��T*��1�eC��n5}_ꢌ����N���ԙN2�!M^o���\��FڥŃ�D�U�w�/8q>D�X�O?_�җ2-���Q"�q`����T 8��2�W�����ei\��x."���y��Ԏ�Α���
=W(w\�$.�<�v�C��Y���9��'Lb�Nr8XE�MC
�C��2�%f���4�6�/����\6ž�k��h'����ںZZ�?9~L^{�5���u�<��B@ex�S#�X(Lc8葇8&�L��rsP�`���a���c4*��1~�1�M�1���A���C?�C�`�������=���W���a���0�F!��kS�\�7����/�hW(s���7b�N��M���J̽�=��m�;W�?�C�*���gJ,�&��&���֖�j��w�RT+]��@��Z�)%�':�h(jC��*h';��$Z�n�by�	c�>&�$��b_�ܐ#w�b9g�o�0CG���3�|�	V(�o?�m�+�-���p��"k�kr�����ڞ2��N�+���j)�w���HOEAǴ��÷�T[�<��Dà/9��֪��@#��F7�N[=���أ}��n_��m)G95�&�ᶥWؔ�k��u�����S�&꥿���R��r���@�벺yM�db^�����v;�5�q�q��K��3H� aM�n�3�+�-5��%�
&���To��M�zl}��!�Ո�q��Q�А���aS�xjT ��5k_�ƤӖ�Cõ�E��7�hw�y�P��z�!��y�2%*�J^%�M�S����}��z���aiy����AO�A���������X��i<�#%d��,�:J��4c6=z"�CeAÂ����A���`��!���C��ׁBv�<��t����|���'���4�G�ǔ��13���A�!bB�o\��g�0崼�����~�03�*LaP��7wW�E~��G�5�����#d�c~�&Aq��9e%�a�u�;#��Ѿ)h.�Ƨ��ڴ���p���m������P%�yX��hd2u���5��y��͐�Ї>$�>����i�r��5�7�'�}���=Pk���V
=1-gu�����ֶc���9��O��G�K�� D?T��"��]��+�٧?)������'�����	|�y������,��Y.���!�+?�ą���`�[h���j���*4p�b]�l�u�����ѿ}2�r����N��JoN7���^G���W^�e�ؗV�KG�(�����QV�/Z	��`�R���_#�٧e-Y�=%�������3R��i.��,Yt���mZ.s(et�������kMYX:.�Ɯ��r�t��D����%��s#Y����p[;M�!D����y����{�%��ܬ�n�ʟ�ٗ�ܑ9�@G�=|�Ʒ����y�"��5�t��fTyW԰ʸ��5-)�R��JT*Ky�������!�$�����>%�K�
����>+'/\1%d8�&4o�G>�s�SG�R����z�y����^,�Ǻ>��c��|�~���(�_�N�R`�7�P�X�mP�dB�h
A��S��?�@%��!�ar*i��8��@G�OEF��%X�.�6s�O������ ������}�*���^����N'p���c�29<'�	��yK�bFTB�IE������t\�x�0���|�*��G*�p���4�m��0�p@�p}��CT7�����5]��~�QR[w	$z��̈a�c@�#�猵�{>"�Oh��}� 1��_�{b�` a}��:~�m����D4zèAt�'�W0��.���U�a����=�����>%�,���Q0:���<X{Nٕi�@��v
=M㼁��Req���k��s�q���o��DU-�r��!����uy����t�&�����{�Jd-��y�\�faW���*�M�!�]��$˫1\D!�r[�$����3��ɓ���=n��z�yBPPϿ��Y��v�����K�<'�.����bY�IN7;��,��U/B�D4H|�Y{l�igu@���e�(wZE|8x(�ή�]^�`��s���� ������d��a�:55:6%-�$U��ݑ�#G����*PG���	tEg@�ʹ*j4=�����8���qƣ�ys ��V�'04b(9Dc�`��O,�{>I�<#[��Y�
j�K���C����ɓ�'��_�Y5F�8q�J�H�@}A��.F���۸�FLo�/�A_=x�:s�f�
׌�f��Y}3���#�����P���(t�{�#��8�g�����2��\�����d<s�T��Ԩl�p��R1�:�4�b���(�k�C3S�P	���
���4 >��6"��]�J�cE�6�!�.s����c�0P�f2a�X*L�)Y�BC
������T���S�M�#0L�0�l�p�ib�0�A%GE�9cI!=��`��j�����a�y?2�ke��4<x�ҩ�H��1�c���z�xF�G�)����%vP��l��'S�HH�Cb�#)��~��3aF^���Խ�(��8p�i�wR�!�?���i��z�cI�|D��T걤Q�K;��NIEƄ�W�Vf:�j���-k1
�	��&p�@)�eU>;}�S����u"�L��W�/�@�����&����9rx�� .�ZTk�&��,�Ϝ�J�&���ߒ�9���H���tP���+�+���?`B!Q�N]�yF�R*�j���8�{j;�� ̛��7nN�+q<|������Y��xS�f�� �aGC�X�e��
�B�d����U��ڐ箜�F4�ӯ�*��3�.���#2б,�Rm뇋�_.!D=�c��ʧ~�c�<W���/�"�p��llޔ��9}�����lC��*�R%U+��Q����J5��)�|�'+�|蘔�٪p�����!����B��ݦ�G:�U4����+r���~����kWl�;q�lo�µ5�&rg{˺�A��$�):0K=��ɖ�5�:� ��3�mn���is+'RC�LelPLP��hO��gzCc����d(��DH
�� ���$#����zC��!�~��4 <jz����r5���<�#�D0���s�<9P��!���;�6�>�m�è@�� #Q��O��i���FWX�@ϓs��kY�g.��@��c �}X.����Ȩ���4�8��*d��y\a��r�����{`�k�F���uF]�+ehdq�p�3Lð���߬�`؞�<�ǚ��d2���ݨ|���0�>pm���^}�+f$�|�>����ڟʴ����V
�i!S�0t��^��K���s�q佼�Y�� <b�{$�����ò�ޔ���/�͛�J�����ݲ\_ݒ5
͝��wU���V��B5A>�Y�Q�y .1��{ �(��ԪG�3`)6��j�����X}��/���4Ԟw�=�z�iн�x���k��d��w�X��B����.�G�ʅ��Rj,JO��ܵj�r���;z�9�d6�X҈�v?2�`
��%>�c���\X�q�X�u:NQ/�uc��VP��TÅK���LY^y����~Tʺ^�5�f�?�qy��3r��We�R�
f���-�6����iE~�COIww"o�|S���dyiA���+RH��ܲ�|�!6�{�:~i�3��5�Pdiy�,| p,4��V~�1nv ݗ+�2;��q��t��R���_�/����G�ӱ_��_M�<��zS.]X����{Nnn5%_�ˏ��G��o��%���䭓��3�U���c�n�wy���&�w*2�Co�lMᾱ�����>?�a�V���}�|'�A���8~���9ư&��bH�����5���d2��H�,�\���J�X����I�A$6=?z���e�r��W(i|
<9Koy��!�yn�9���V��`�V�76i�ܱ���AC�V�1�5�ѱi����R[��=蘻u�8o�3v���-����R1��k�)��/;�Qo�D묘fф�k��@�K�V(;�;Y4�L~{㍨�����z,W�X9�Ů݋3�J�H�1	>�9k����sQ�$DXE��*w<�(0�h2b��+;��t�N���}z/�s�뜿|-34.��n+:���ྡྷ$��:}�Do��m��(�N�B2J"�؀P�b�r^�L\Ո�!�Z�H�T�:��v��><��b�93;�3U�8g]�_����Ηͻϡ�]�7.T���2�p@���{ݖ�S���GV2�h 3��R�UU��f��? UG�Otc��I�{��%�ڒ���,��U��,�ɭ�X6o������ؖ�����z�'`gkH<(ʰ�Jsԑ�Cw�9Q&56�WS�]����2��H�:�xb}���Nlñ���������QRS���w�z�đw�f���f@��+����7�ȓ��r�.y��9���_~�_��������37ըiɂ*�B�(�����Jg(2��w{K�'�F�(��=�\cIn^ZU�eF���:����T�����|�'>!7nm���W�ݏ=)�.\��j�i�L��e9r�N�LH�gG�Ks�,�8ƻ��ſ+_���B����ܐ��ȏ���}��q*KwGǪ�X��R�ycF��@䓟����?>i�R�b��z	u�-���U�_�z�<�K�����K���ڪ=S������/:�q2[ב�D6h�J�:,;�WCjXE�7ڮm�#
��k0�u��ǁ�%���ʒ��ng��ַS��I� ?TI��g�L�
cC�a�p甏�Ϲ���\�A�EGEb�� �(����,*S*%�e c���$�����u����+z�T�@a��Q
��أ����`�]�p�>�qA����XNw}�ke��Փ�j��SO=�N�-}�U{n�Ռ7Nы,�(�R��9Y�`N�����S��L�ݱ��)��aGH��gǚ�gd�"�Ô�"i�팕|Z��B�"�R�8�5gg���ow0�rf��Y�0:���[��_}P6�½����4Fi��h$~�1����aDíO�/cӽ�:2ā�R���"�Vu�:�o�q{)�<$$^�xzQ����na��r�9�_���ueF*�`�/-�ZS��#WG�?ri�j�i{�¥V��L,���Q:��s��Uf���,�����lB���S����=E��«�"�`~An���P!�W��N����Gx��5Z�/�ح>c=�.ؚ*�@u���C�H:� &����(]3� ywz��Ã�?b[`x���~����4Q#*��6vk9X�^��B�V�[����Iʹ�����s?�I)��3k��/���J��ll놕�zFGe��:������7���]�^M��}K֯_U8���«�;�U����e�5������wk�
\����YTT��fB����/�'�W_}M^x��|��/HefQ�������9����O����_�e����Ͽ�]�;r�<������3��������qD�ܸ!�g�ٳW������/�"���)tx�Ǐ�Ȩ�6��,̡zE�-�j��hGe��]�{�G�5D�%+��4�yrT��sS��`m;�F"��IS���瞖,V�Ҳ�M27J�6��C>q��\Y��C�WLϔyNzS��{����;��x}F�X
Eb*~����=*e^3�0� HC$?��HnX&�g�k�Ջte�����Ò:�o��P��ر���K3�"��7RCx&(B����ds#ҭ�D�J�팛$�aą���q�ݦD��\4��!�4��3��R3�r8�ZJ�zpsN}��'A����V��G��,�!S�e����f�#���ĚV����{��m�Ї�=I�x:��V4]l�cچ�u�P0���H�
[��`R��a�B��!x,���-��dai��ES��(����hB�W%]�E=Ra�Eg0,��ղ�	O,/oV,�$���H=�~Z��W�T�5�ׅ\�]�!B_XX��Ջ+�ݞq�����Z�}����2+�us"_����{���g��gO<>ò}��pƌS�bﹺ|����Qj���ac㠆��\I<q�sz�q��p�4Cbnv�ʺ��y,/�䍓g�s����?�����z\V����U��_����w�'��}TΨw���s�籾Ց_��o�bY�G�}��������YYTo~aaN"�`.ݸ�J��Y���5�^�-����h���#wHO���"Wol���u�+�����~�V�Z�����؃�ʋo������<����8(���[��3�uc[������^|E�:/��Y����ߐ��&O�}��d�Q�ϏeN7�Ճj���m�Ns͔��S��~��2*�p�����6�I�H��܄B&$
��Z��F=���*�(�6^#�&���v�Fa8�S �/�����gX&GϞaV~��	4��2g T���� �iHX3E�c톀+������g隠 �OE��?@�|����$�CF	��p�q��ѻ��jQ;O�K� ������O]�t�����7D$q>v���/����9~(r��	Z�A���N&C_^Ȟ#T���yB�5�k8�a�?����זK��2����/���D�c�p�X��@H�Ź��0�0?�ޭ�S2�j�N.v{�=���S�o?�t�W�J�O�O&��/��,�~��� ��ys����rQn� ���N�zŨ3F�>��<�ć:��k2b����[��eZ��mȱ}��<,Rx����峒td�º_��(����_����
�JUnm^�J��JX�8a�5t�`�ZX�Oݸ�q��f_�I�<�4Q�W��:�BQ�;r(���;�U���/ب~��[⊤�pu��9"�SOx���Q��Br.L�(as(���	���t�-���:V\6/���U����|I�����|�ߒo�y�]O��k��ȏ˱{��j@��\۔^sG��|�����릟��j�U��U������EN���k�T��+W�����&2<}I�7��*�r����}�.����m�X,>l5�(7;x����ɋrqu]v�H\P�=I�2��ʫ'O��ѣ�������▼�k�%G/�xؑře�����ֆE��AGV�g�{�g�����!�s�3����:C�,�
k��-�>|��S�-��8C�Q�!���)���a�R&���(��qPq���=��Q!g|h��`�*`
�0���h��L�z�q�cZ�%y��{"Ush�г�ӆ|N^�
s�}X]@�W6�V�� Ri3=A*_$��ox߷t}2�l�1������)�*y�i�А��*��܅8�5�q�wh�G�Ǘs�REIf|p��>�|�D�+�n��a8�f��@!��k��aF�؍C�_cS+[W���7�������GEn+����l�"2�Á��=s�����Q#�[Χ*\��w=*���W��5��׾�@e�� ���0O]>�U�W0�&
�[kb^i�y�����Ps[jZ�>z��{���hh	����8�]��*e����-����*�+���z���h����̡��t�SW0HP��h�g�������Tu
6.6�z�9�k�AI�%X�����K1������Pq�\�z�=z�~{�G_�x�V1��.��¢�^�^\:���<�ݗM�� �_8 ����v�/s�Ey����zk����(�e��%��HTg�׬?��\M�r �Wd��Br�!7�GqK�˥Ʀ����4��Q"K�N��K�1�R����f%��޼���iI��A�i����,��#�S9��몜rx�yJ3K��ܕ�g�y��1]�}}����[�h�0 QŇ?�!������w��^x�¢��ԛ�R x�FT(N�_����r�̽��'
ܐ����;����"zI.G�τ&iLI C!Ǽ+	z��wo�[Z�����?�9�ܹ�Tݚ�J�b�
�`��-hFE��	��V�M�ml�ډ0(("*(��EQ5Q㭺ù��y���߻���o�ϩ���t�q��>���7��]�r��
�Xk^��s��n%��ސg1�]�E��If��8,G�#��`������ñ(�-ޫ{�>�xt�J-]��u6 AIU���PP|ifl���ƜG
�](t����7y̑&�c^}\��re�k�8N����3/b�`�5���$766�q̕g1���M����e�iyh��a��q���7pp�04=���;�{ѐ����r"_� ��ge����:f��}?��ף]�E4��5U�kW����=N�a9ƸG�X�r���h�k�ic�nm.�ɓ����C��
�����c�=.k�]�x#�o�(\�؅Ҳ8���@��	���/8t�
J�D�}��T��k��#Ʊ�abQ ���{�1�Jf(�]�XUa��ϼG���'��V���|�o�,}�����R�0"ʽT�IM��� ��VER�@�j  ��OLp�g�
߬�@$�!�yzы/�LP��-0>e�X�ঀFVOyر�h�8����$�9��r� �յ�9pP�̳7��g���.��G��ӏJ���jX��9���'ͱi���j�|��lH��~<�x|ĺ�A��(�s\�P�C����M�djfRM��ue���z7=(f�D��xB&'fU���8�d��4�ŋ�eciK�W�g8���ʅs�lӊ�<\�/�D}\�׷%�bx�4�u�S���w<!�����������ʓO��gr��r��i�UG��� @����]I=��Ɓ^�0wZUz8��)�(;gQQ[�u*����p���"6ç���q�^�{�N.�^�߫�����xn���¸��=?�����"A�?�{�.C|l<�o��0^����W�\�߯[TfD�olQ쯎�^d�rs�s��A��H�y��.L1`��B����K� |�<��q�p/��E�^����tD1R��XY�s���M����2H��؉�:/�.��ދk�g��^�Yd(t���#`��aJv}���Cu�{��G����<̟�h�����@�#N��]ѓ��������7!Q�����%�ӓSrp?�r����G�����\h""K[:���;�1�q �p³Fa���i��&,I6)��/]L��>!Gx
kvT�ɱ�l�-���3��c�O��������yTz�z���^vg@�elb��+ڄ�\F�Z�|��J�;���C��}U��ǣ�l�J(9�+9�(L�]K�d���$
�X��0�������,�����a�٭��g���O�v�� TGȣ^y�Pq]Ω�LUI�O����sv�	晫���'�й�H�(�ŭet���Ͷ,,�Qe:-s����gXLm�l�̯�d���Wy7�������� ����W�`�齏��RmD���`aK�������F	����� ��X���MVIT�PXYl����@�&��;�����jԓ�W�K��o��j��ڑ� l�75tC.���ρڥ"�<�r̞t/c��n x�ׁ@ED��z]���.�����u?�{�8��T�p+��?33������J�W��¸��?���"�X��;��Q�E�����>o����d��9o�" aqϴ�GDre�
���M1��>!��cRF������w�M�T�~N�=`��F��.d��"�{��n�C1�쯹'�a{�@�X����r��c;�;���X������o��^��eyn�9z�s�<�O�R�5�<#{>p��0�K�����v����B�P��ڣ�a�ۅ-�'q����%L��3�`�q�F�۔oet2�ΰh{���_�/�m��m�裏���E���,�5M��םl&vtl��B]aJ�U��9���0m1�T� ���Ar�v�n��Zƀڗ>J��LWorm�'���[�����ٔ����X�6 �G�Z6�O5� �%CC�e	ƴA[�V7��IJI�ʦ3 �@�8�QR
�-n.����ĉ�l��0e��xB�N!EbM�wL��Qg��ڐ��s���C*[���r*�t����k�(m�ducU�Ty.m��2o��D]�k\�ԓ>sw�{�,=�>x�tt�-��ޜ��B�}L(��v����*��C�,YiNα
@D��"���P�"G|B���⒜b]���?++�.JoM�$����o�B�T�>� 5ָ.�]��+�s�/��̄�P��A���^:/��{��N����6+P3?�u2�5� ���ҋ��yу�lA���5����b�����8/:zA(:�w �{�`���)=��u�N+�ݿ�
��Mε��ߍW
Eo܍�̈)(�b��"0�=�"j�,� �����@/���c�,�N���pC��������}�*���Jw��F�3�qSDi���(���{�G.k��}m����b�`o���'��+F��)W�������`νϼ���9�u�mu�i���������G�2���jw��{��n'{�"�����h���#�����ƙ2��g��?GZ��G����4Ԋ�d�6!k�-vA+��-exS2<>�>{]0���Ui�u��r�m_�@��6���i	eV�iI�	�<g�ڨ�9�B�y�)��*\���&�B�q)(�;�C,
$@��Ӭ�F�P���O�t����8�`��P&J���k�H-�F�f�g�{�Rc�ʅ�d�����7�e���,a����aA����p ``B&�Ee�����#�	���6_��a jF��X���C���&�0��,V�����@�/������r���W����NcJ6{��(Y��G��;t@���YS}fἴ��-HU����!g�^ 5� �+�����I,,�.�B��(xL	=�R�$}�����`���O���/�^���[����j$���CM8(d����>� �/�U�=G��#YYG_�2�/��8���Й�:pX��1��dr�<��W%��r`Q�[��+�Pq��ȱ3?m��b(�o�Q88����l�v�֫�y^�B�Cp�n�ő�k[9?��*��t��AbV5�(lQ�����Ѭ��C̑\�x����y���m�[�Z#�Y3N,�õ��� 7`��U�j熘�w��C�<��6�r`b_�u��*���7�B\�={�B�灡���^��Qo���N�륈��1t/�Ah�p���g�QTv�!��9�/_�C ��U$�
k��t1҂��r��2�&�ÍO�5_��R�w���� qO���8o���{)7b�5.�G������p���M%��,Å%34T���.�2�ȥ+f�t�v�A�C���
Rl#]8�{�'�~��&)�j7Di_AU�f�k��Rң�� �`��wV�nx�X��,)��+McW$�?N��~wD#z�Q,�� o� 6"@!m	VVBE�#Jl*b���@^�J��g �	b�j��U��٨�Z��z4T�@/m�k����}������₴[���oy������E^�����{ Qg$Z��L���'V�O�V�N�{g��(���4�L8�B�M��7����e�@b��O���u� �/��\S��r�5ϕ���4�21>��ū�g�C�NZ:�Kg�ek��,/m���<�י�������9���:�_B����z&f�����I�j��ͩB`�t����ȁ�t.����k^U�E��aW֗�n8!o���j ��~��djr�����N��ܼ��*�ğ|RT�<QnJk�z�B-�z�k[k2����Ǥ��+�URe��\�s�����'�k�k���ԃ �Ɂ��U���׻�y�N/��V�.���)6�`�m�_�u��=�^0 8Ax9�禍�<ʔ �����i��A�)��V#�S�1�z��+Q�������Nh!��TWnΊ�J�ñE���:����y],�J�4C�=k�����C�P�<O7P�lxd��al�6��ͯ�s���ϽiJ1/�!�"=��{ӗ"[��1�Ɓ�x<U��������{9���'<4_��`�|��n�Pn����(\8�����O���XG�����{0�p~�o�)Ϯ2R��|��:��S����d�y�P����ޅi󫋗&ݝF<�G�*��6�.��SRR!ߌ��TxE!��S�|`�z�m�y��G���S����z�VWnw*8(v��%i?�s!��R�w%��z)�A�_(v�cr����7z(u�w]QO0V/��R� �uy�5iT����ũ?"�*�`C=�~{M�-�nV�V��c= �Ճ2��k��i��/�#��mOQ;ohL-��:��3�p|��9/B�_Q���z�Bc5��6��I&�jT��jD�*ֱ��D&k��OU�;���d{g�h��6�<��Wdv���K=U�ωZI�*<�y�Y��6�Y7�t�]��0'��i��0i[� �Yt�J������C�fM?V5U���Z���M�p�9<)��U�WDV�wdr-VՋ��䑇� o���sea�aU�+2=yP���IWZk�szB�C,�뗘kGh>f���Z�%]�b\�k��uB�{��=L/CBn	A�@���N��%BPHŲ�e^&�Q�$S�.���Á�A@ȹ����������k��DU˼!z�(Mr#�S¹h���π�J��kg�&|��c�Y�Ӻu�FCz�xV{~C�Ë����<���F�ZX�^�0S�n� �ޯ+$W|S�+�#�K�\	S�+N�o�VGY����V��?:�|D5�w)Z_?9��v<����!��J)M%3� p��[��=|�%p�����8rE��ׁ{��ׄE�������>�G:���jr��#/����YL�!�W!89�2"w��r
���aF"� L�B]}��E��
��Z�x<�m-�@��#M	��%����u:���?3Q.�j�R�T%	���Q�q28w�R4��Q4��|���t�F3�Ի��X<5Y�&/m,GC�\��U�Ywvz���u���!j�ި
W�GVo<���9d��hJ�#�1�q �@��
=�#�R�1��(qT�2��øo�����+U�T7 ��WRz���\IZ1`�TT��7'7<�.�{��`mrEFy��96�H�Zb�j����j�ڇr�ퟗ�3�Y��ݗ�3K�Q-�!���իF8(*U��G�T���=��C^ �	K�҇�9���
�-�A7b�ϡ���5=oc��~�rJ� ֗���d�L�
���*ן������{�=���[H7|�.۫r��URkJC���am~jFV�6�a
v<��A���§	�#q����B�`2p���UWC����!}��C�riAf&�����*��|�M�ikc�FۄzzK��X۾��³?���ԫ�m�@�R�֎�\�H����>�
G�����)�kH{ԫ�LA����A��M��u=����4xY��Zv�e�޷:�B�8/~�X(�Z]�p���e���.����k�V��wՀw�[�=�<��w�(���7����zq��1~0@ �9h�d]�C�˯pnS@ә+����u�^��d{nߍ#�`���3�ge�1������pI�sB�9���źq&ż�߃Gf�)r0�+{��\zD�H��qnx`�<�eda�{/��Q����=uRLx䢘)����Ϗ�A�?�3��g:���"WX?�p;k#��	V���:ZT�W�B��r�E�NG�OI�M���M���v[����F}�k��U�cC���(�!K�iX�!3"G��{U��I�7w��=;��������^{_���	������u�m�H'1�Te���0`"ƨ��z�.*�垪݈�-�S��4 #��؈���%/w��A 0�5\�z���B/ð�&� ��(�Z�k��������䃍��cd�`y��xF�l]�Z�Ѝ<h�x!B�ҡl//�+�?�禛,6�|�J2�B�)J�XG_&n /e�m2p]�cB����i@�y0�H5�����Vé��}�)���Ŏя��\��}Ӫ�k������7JMixb[�r痾�M���6��XE��Z�u�t�1i��i��҅���c�!N�c8��yoaU��R'�Yuv<���Ғ�zI�XI�̏�sĲ��IIW��%��g����}��_��!c��EJ����@i8�[�Miw!��r��IV$DC�����YC�!r�H=���4�M&)"]H���B�������IM%�D8"�j�Ig��܏zxm]�h�[�f�A�Bh;Ry>��=��M��^�<Ȕ���)4�=(nx:�����y�{9���zワR؍�r2%5�ʾ,u`���9(|g=s�W���{���U�{v�;~��"�vp י!p�V�x�<ރ�Dۼ\���6�����ZW�n�I~<��J�z�[x�ָV�vo��O���E,����#U��ѡ����%�Q{�`[�*eB�7g�s� ~zY�q��gQ�b#W�n(a<��k��uo����SO'���e�t#�=sD��\^�� R�z$�s���8O�PY�	��b_u?/@�n(���)LJ�p�LC���U���[j3T��OSٚ.��3g�Ձy����[t�N�O�t(�����	q^-U���(}ťKKw������?��?�[]����Ss��	�����W�C��X�:Yu�4T#i��2��*�u������H�^�d'^2���,4!a&6b]2�>]h{Z
)hz�Qb 	�,��^m�'�HWC�g9G��#�ߓp��X���]+��zA���a䩤�dGKѐ".1�r�6H�ԛ}(��Z���u����HgsGJjL��N5�~(x�X��Л�q>�R�q�Sy������ok�[�f�<0V#��f�9�Ǻ.qUN�*p{U�-��6dnfRZ���W%�0��G�?'���Y���3i*����?=5!��y�>vJ�<|@�^Z��ￃu���iY:N�g��-�� i��[�1FX��HF�6ij�S2���7ƽ���4)�@���A#������:hzwV�Wɥᖼ�%/��z�	�z��G(0���[��7U�[]1���'���m�GFG��˟;�_VT9=�ȣj��JmlJ�z�j�5*`�Q�F cC!�
ͅ���<#�IF�NCVP^W$��k�7�\�"�o�uϩoomgF�^� ��|���-\��������s
8ɽݩu�B�Χ�@:7N����w5 $���Q�l[�}���V8��Vίn!�Q��\ā�'&ǲ6��u�u7�U��=j�s�
И��,�����Ȁcn�`�9AMƳhE���xs�kY�+<΍s�SW�.��y�Y#O�x�q��q�:p��u�` <��üW¾�������t��wߝ�݈s��tT�ü���� s�2��u�T���W��:�Ѡ،,(tth[Z�d5�u]�*��#��eFZJZoɉ>���_Z��>������_�{4Ln�=�
5.���n�`�o&<��y4���G_���!U�zS��NdS�r��ÜHtD"%�
�a!|��+����Y���:IJ�4�i��j�B#�q�Gi�Qc���P�q�$�{�}�&rZG�3�nVw��߱q�[�;��#*�N{�!w����þ��Cg1TX���R��[���� ����F�w��R�^_�ז��,�}��Ժ���>�4X�T���T��t���ڐ�Ld^���A sj�%��"gTU�vB=�I՟�** \T���lo^T���ϮC���ϼ���|��a��p�y^t[8w�B1e{�1I��d��C2=��ų��,��lS�THo��xק�9�ip�Q���2+b��g��l�r��?A=ÀJ0�!�,˄�_(RPĪ�]��9:7.[k�277+o}�-r��Q9~�J6��h2�2=3�e211%�.���������[�ron(k�[rq�9r%����!�87\uL��Ve����G��ʠ�#�a�%�媅�Ϝ}B/-gJ�ޏz~'O��uU�~����k����V�44N��R^���0q7� ��C�@�"8�
4�	lĆn_�� 8�i8d���~����<�n!����:3
B����%�Kz�G8��n��f���E��p��e�-��gtĵ�bO�:%�~��3T�<��4*�Ν�9����|�7�\}��y�ZyW���0��=��#w�q�.e�
��`�ܯ+:XKS`~p_�җ8��T���qg�����$�43d�����T����x���z�[�"ǎ���D3��$���7~�7�q���Ǐ����v��޴C�G=��W~�W8��v�^4�;��N�+G�܍F��w�ō����}��t��C���gʻ���P���������o{��2P�K�{�G�GY�D��ds5R���|�����h��q�
����i�%zj����4y�;sK��N�����Ǆ�{�-��xpt:����B�&U�����U �T�O0��o���ty���Y���7S�VJ̳�'B~xo\p��N6L�3�6d-vh���Ήӛ�n�FQ�R����м�l>P��V��Y)5Բ�B����]���q����e��U�5��[;%�U��4����Vx�)�|+�K��L%:VP�%���u�Y�o}��X삦�� �4���Th%4�c�:��{ý��a3�� �:��>OW�Y���©]U���m�𞞗�N=[N�����~��*9�����1�ssR�����
����B�:y���r���IU��ɱ�4'З{Y&j����c2b�[��<eZ��rI���}Z�C���5u���1FF�2�uz\��ι����U��+��]o�#G��SW���՘���6ט_{�K_�Ȋ�wZr��S2P��z:g�8M����nW�`^ϋ�8��e�t��2UW�G�X�O{��J�M���>�9�S�s������0���j���6���iS �[�%���ۼ�~�^(-��Q���~�_H_P�E��^��ڔC� 0�2����=T��;poJ���Y����h�A��D�����y��Gآ�.�eV^Q	�ȏ�����y����,�E��w����3��Ͼ򕯔_��_`TG��۽,���#r���`��G#k������-�"�z׏�x�g^�{����L蓟���uǝvu��(��o�E^��W˦�Ihr��tNa��u��:f�z�����Q��LB.����7��^���s��t-S�Q�����W�bu��v�<����^Fc���wޢ��O�� �����ȃ>ȲF���<5V��=�y��n"�l��nߺ�sn�����?0"�몯f8
�$��\}�ƚ��-2)|?qk:� o������Uم���zֳ���~Y^]a�
�x`�g8��xu�5��b�� �Ĕ�g�<R+��_�W�(�e21`���t�Z�y���QKߟ�+�8��	%j#���	���O>C��#�����ۈ�(If#͛�<�pҮot�6
��^������ظ|�Q�8����:Ґ�-���Ӟ���ek�4:1"��*��9E!O���6�*��N©�*6Tϫ�YN�csk$α�F8=����z���j!���f3ĩ[�"��Pxb��NX���!��ў1�W��M39�*���P�H)X�C0 �AISd�2^��A}nP,G��z5c��-#g<
y|D$Z�yZ�BIv���^�B��'�cc�.֐�A3T	 �%=�P�5l�Ko���$�>S�h�M
��s�r�+_.�z����
�F3x-�,�鵟'N�`�g����&Ir`xm��X�)���o���P����R�}2�
,x���.��1ѕ��;��:�m���Κ����C��-���?J����GU����u_YZkK�t7dL���_�y�k��<��U��9z&EJ��ّ��5�WC�P�zpsS*<��^�^������gے�G�ȹ��R�����u�2M�616��&�^s�xn�/3j�P����,y��@�������3��N^������"���A����?�C�}6�pF3�>�k��L#g�+�&�p���Զ�~�]��V�u���I_y��.n�vt�N�gU�9V!��IȔ��5���FҸ���7Vj�4���Ս��@��g��<���{�P~���\3�+�{�W���˪ ��j�Pq�pj��ӏ��xϽ$g�����D־�ϫ��bcx�0�����1zx��a��!�JI��P��>����� ���^���Pc�d��%���;��0�`�yn���fy��Sǭ�y�8��i����3� ~:Ҝ)-��#�)��{����&�:O��t8�#pD�׿���屇fo�^ې�ztf7�7�LtO�ļ��C���|�>$��s�#md�� �BE��ڪ�[䵘�1XYYf��\�z�������ю>�T�ų��r��~��HV[�UU�� �¡���կ1
٬�)#G}D&��ن� ���K�O��b�l��x���u��Y��%����%����?q�����K�ݡ^�y�c�yC�<qF��rq�T0D����s=�A��O�B_^^�8�p!�V���L�[��<�$�9;@K/:;��.��k:�FN�GO8�t@��6@qq�3��CƱ{0�A��/#6�ӂ'pFz��=GN����A�����
X��aA6Y��
���=��`�ݢ���x�B#�о��`S��Jk{��;�a��4�'th�Ȑ���		`��B�5�S�Z� �`V��G��˺=a�����C5U�c�)��U v��+�7�Bn��7��Uy�?is��oxQ���J �q=�pI}�1y�G���(G�?���Ի���Y��c98=.g�<���+�21���6-U�o����_zL��Ⱦ�}�+��7T)_���7�^����HE�W��"�'��=�9�=��I5(vZJ�!��_�,���P�m��1��l�Ѕ'	/!�;�S��)+����WO��0q��	���?o�*������i9��9��W��n�l�`��_��,'���Jv�1��*���^��y��'D����J	�n|��-�>���˙b8�}�{��>�O��	���b�$P"�E.�����w�}�#�o��dm}�Q/����@	�L�z(~�_��2������{��#e�g$Ld�������<�������� �����˿�G?Cz�� 	�s�Y������������@=��(�\Tcl]=S������8�?���( �4�J��{�-����ϝs����ٳ�����۾�C�W
��0�ʋ�z�+:���1][˗t��70�ʈ���4,�P
�?� ",Lp!�BD:���[��H��Q�Ȱ4�Ȁ�@�#����jo=5�;��&&'�v��и��#�<���W]�3`5�%(Ws�*��"�p{�f�4���c���ӏ?ɵ��v�� ��Qʇt��z3@|Z�����׾�55(O�<�Ci�>�F����3��b��7f��uLi��t\��$Wʘ5����!F���U�:��5���~Zz�Ӊ;�N�6�+�����ʇK��K�%&�N�w�3��Q+ge��!�R��Bd�x�y�(������f��w,@,����Sn�uԂ+%v{�߯��%��C<���BOn}��:G�~��[^1׽FI1����1MC��4c�����P��D��}�&V` Eu�Ȣ��kE^xn�!����,���TX�~�Z_���|���I���k��� �JQ�_#�~��u�1(&o� ��J�VO��z���(���OS���m������,���p/,���Ӳ��#�k#ٷ��Jz�
���p�nV����NU��\ghxnnB.�;'��������T��$�u���;4<��a����H���{ks���@<I@)#��	�
9E�����~�>����(v|~jr��SW��>�W,���I]�S*�,�ܖ�3D��jk�ʽb5֘K����hy��?���(ez�q�hRD��nxA34^�'qiqI�����YU�[�I��2�8z��3�� �uc�D��J�x�a�9��w�#� �;���7^�w\g>�L9�V�x}emM�\����9��mD�h�Z)��yuDF��J�7�At�¥�\CŒ) aP����W���Zj���!��M�4m��qx��2�c���Q���!k�11�E�N?y6�W�Zߐ�y��s]6[;F��Փ�5C�7��iI/����� �HS�K�z��(:�!���X���Z�������uY\^�_#� �p�M�ΝCO���� p��6YKo�i9���Z.�U�71?PZ*�Ѿ�e�%���L�� '�!a\`ȌP92й�9C��x��I�(`�"�x^b �f� Պ�L�@b��u�P��V(�Ú�}l���.x@���I4���!����V;����R*��0�յ O}[�aM�`}��P��� �Cj��ԅ�-i���Q1�<$BJN��F����B��Ӫ�+�F�1�H@M�����rlPTR�u��#Z7������шE�dG��i�j�73�\\�w����|:ʕ������w�CuKe�݅��!B��\AI��������a���~��s{.GO?q���:�S ��j��НP�����n��a�A}`M��o
=��ɷ�Û����r�����꜏�GU��(G^�a/	�5�f��f�.��7���Ex�bEX��'ev� Ü��M��n��2=�_F�W�?�Ct���㏝�����lI7�yZ�/~����{����7�HP67T᩻�h�h���\l}�e��z��rP��@Hri�����p�����j�C�0$B�-���)�����4��SW��z��KK�D�{�����h�&��[Y��AB�G#B�y6���1d�B�4� T��	�״�11<�e��LF�(6�a��{Mh[�]G�XL�����]W��"24�����Π��>"���c4������A(�9���a�uU��NYT��|�����*)��,��v����ň.\=��a2������[ɓ92(j�T���t~z��.��T=���q��y�>���gg�aX���w@f	���y�� ��=z�P����0�2��j��#a����h!49����|�#1�Sv-4C%��J��`�AHK5sC��vw%;1ah��z�;-�ܢ%%��gc*o0 ���@� a�.�y��+�����B���P�'*��n��]đ�%�z>�Lƹ1^����6I W+�
{J�N��=�B�}���)���_�$�s�a�GzRQ����i���#i�-���4$ ~��yхQ?�vN�{@��I��9�\7�U
^��^���|#�k��<��*�d ,��$��?�]�#�]�4
�b����R�&0_���΍�<��B����ޅ�u�39b/Fv_Gq�U����k9�K(A����8�F�;���xB�߁T�U	%`�H���y��z;*���W��n��dY�^hG�..���������[�.^�ݴӬ=/��Nӧ>G>��CJ����PW~n&����,D:�{���7�T��b��J�D�kSR/˺z4���+r��U�����ΜWoeBΟR��O�?&���������Vy��S�(U	I)x�)�H�*%�,ꂔ�x��V��#�3�g��0��)4�л�zիdrb���Kz�������h�$1�~�1
�����
�Z#��Ԝ!�'f�����7�U: i�)�K�Dhu��W�(R���Paưg1�<qTz�W��� u�U2�Xfi <�a�$�ı@ G����34������[��^
�-~#�*"ނ������F9'�$�̥*�/^*�k# ����B��w�<��ܐn��OC>��a��(�S��X�2��0��V��[b,ߛ��F�fJQ`�[��賣�R�l�S��U��u�ٿ���:�g�/�^h04\"K^B�oct��ֺ3,����B�#�q�հJC���N;��ԋs�*���}�TM���W׹��[�ю��4P�"R1Ji�C^�`��s6�WT�bS��˫������A�{C���!��en� �G���ٮas�Yj�;�׎� �>V�x�D�6?Ñ�aAnc߂��$*cB٣9c w��
kvR�����GHSV٭Jg��<���(SK�+�$�>`��|�Z.�sp&�fu����]��M�����J�!�<�<
5��,$E��
��U^N1>f��-��jXq�"�=����`�4����F3�`���Xk��.%ði\ѧ��w�\��5W̱�S���o�ߤ/�r⛢�a��n/�lpd�d9I �M��-`��p�``�u��E�ޒ�*��*�Q%�3D�no�HK��_�*y�[�,c*�W�V�ء�l,��Jlfj��noڠ�������{&W��mԪ�H���Pm\�.ɝ��-'�<"O�='#��z��L�g~xnL.^\�����w˱+�b�9��}�j��m�x�<��A���!��������Ol���>�U@S.�ݾ����2/6��½�c�ޓ1�u��馛�ڧ��/�'���m��vNkY�T�O���x�u<C�'x	��P��򏥒�YW�W�v��@ �r1�(�����	J3���ݯ.���yN_S$6*��IOK��� �0+���f��	Ld�����P���� <��)V� %�6�cǹ����^,��R�V��6���-=}>���|�����[F���0�a�X�_��|q��4�x6�!r�� ���Dx��y��+�!�
��4rt�s�q�$p� �x1T�n������ቹ٬֛8���r���(Wq�ץ�Q-�R?��'��0��N�00ּ9Ͼ�s�N����]���#(��ZT�ĭq�0���-.��� �aprP��)�[�3I��aP�!d�a��d��L�AX��#�����e_�X6����$��8���x}W�"ރa�(��Ç�`�b��[�`1"4Äi�f}Lr${�l�x;j�C�N+k�� z��ޭ�)�i8T��,1F){��%;'��w����>����B����[��a	Xd������Un�R��G��G�ye(�7�	@��Wٸ�������\��"�z
}�/��� u�%}�OfB��}讖0
��ـv1�爍�%�u�C�u�CMz����5a����A�H��j���ͯ�Y���oW�!e^9zw#l:;=�0��G�Xz�W�cY|�(v6={�N��6;3�B�*~��ǟx���y�	�x��J2?Ӕ��z���ޯ�k{S�f�c���>����zy�5Wɹ�ge��	ݐUY�tI�*��N:�(��7q ���D*��"Ж�.w�B��9�����2L�us�����t�}_�������BS�^�ߕ�<�c��[�8�ÉI�Q�� �F�B��	z�`Cԁ�̵�� V�
���W~0ʞ���	�C����zn��FV{l)/���s���3�Ye��zmL=u�"d�O�$���
qD���Zb��s�F�a֬�T��8��{#g_;Ŕ;&���)S�'���+���Ag�'�M�-ˑ�f����d����p��S:*kF��٩���b�� �\z�pp�;��{pP��|82)�3����~���F`W�V��c�c�{��Դ6���0���ؤ�X��<{�N6>t:"��4��e�`9|�k^�u���|^���IY$4�o����ە,�&�jF�ʩ������ʾR6}�|�am�gʲ>�1��;$<o���y`t��������u.�z�x�b�n��eH�����1��Ėi����T�@�����0s��j(TqV��?"��@ǡ� �7\����[V-s�f�؄Iu���&K���m;��MN?M
=���!f@a����F���	�{���@�kD�
ҁhN���w��m�{\���S߭`���F��+���LRŐ�������p��\X=k�Je^�����ƚ���T����ѕL1����W
$:D�Xݺ�]����<���|Cx4)�q5Y[�^Gn��j��x�4�%��'������衣�(���ϝ�W,��gv����t^=P�3g���Ǐ�[C~��cW���M��XUa�kO��u�D֗/���j	����]/���W��]N���v�Cp}��k��գN����6�5��r�d�B�G����GH�@q/-�X��H�.����3��0 m�y���	5bΐ���L�H%�m�����[�]~�gV��'>.���2e d���2TÚ������LF�b��@�����`J�6��O�>��͖��5!qjZ�����Qk}M�W�meu��7<cA,�n��Y_�����	b�2E���dc���7qJ|�� �!h<B)���Y�e(Q(�}���ב��)�*��Be�4U�XI��6vA�B�Ye:�B�"=%Mʐ���J��"	wP��{îa0\��S�{����Rh|��F��]�2䫆	�ph �Nh'���<���؋������{6��!��[P��.��H������գDmD�  ��IDAT�e�(�7�X�Ȉ�b���V��A�j��w�����{)��*[��$2*�z;{44Y�[.�o{W_�z.���F�q$AZ���>�0ti���^�ӓR��W]��`m�K�8�:F�ށl�z�O�p�E�O�} cAW�^���*�D��2ə�4�;RR͉q�o�e]dl�p@cF��f�g|bJ���z�K֤>u`�zZ�(���t�Y�Bbi:B�ّ�@3z�~��Y+<ω8 /��P�i�!ȎRx}����~�����5/2�C3�#؛�v#ď��`�ʻ.��ċ�q�"�������E�����һ���S
o�� @����4z���]zވ���myZ��4 �z�V�U�+I�*����o�^��hr㱫U��|C�b��"՚u*(f��s�P6r�7刐0}��Rh0�!Rh,O��8���e�x˼P��ēg�!�4�p����2;D�t۝��pI8�5��G��?~�[)P6�79�%d��,c����<�J����?��4�k��V�>BF*0[!��eY�M���u�ygC����_���P���Q��l��Q���+u���krc}�!�Z���1�j���<=����F~���*+ˋ���!�%l�T_Z7���КΚbB;~�b�x���0o�~펟՚5�`�M������rͅ�Y�W��-q�Qq�<��r7�"�F�ᠪ%RU� +�_ (n ��y#��x�h�2#��V u/bJ{kkC�:y���G^�X��7-7�����c�W��E��lR�s����������?# �mm뚏"k֢�E��ʧb�
@��ir��,L��:�#��6�����^O��C���bր?�����)�d�0�+U���P|B%IC�b)6`���� �[��G7�m��Y�R6YKi�ȝEt$�K�[[[␾LF��B�� յ;|_F;�<uH'"��(ň�-#'Dc�(��1�"d�����2���U)+�� �,�Q����}���5�	ekXǵ��%����84�ĦБ�	�،�G�* 5�*��鍤\�/���ld#�y6��W�D�����eg\c!��'yz��$Cb���ʛi�~��`��]9��~��W�^��*�w}Ə(�vAI�{C���fJ`7Y�^O��:��u�o{�`�|���qN����z����Ŏ�H-��UQ"�;
��S����rxC+��b�֒&*6;a/�u�vU!w���ݕ[^��r�s����e.��-7<����$� �촹Xz�!� �E��Çs�ͨP�L>�� �M�Oe�y����i>3�F14E9y�z\gX�c�w�%���Srõ��ӟ��Ǟ�f#�y�ur�5�S9�5�����kD7���2�_I��h�އz��r������Eb �}�7}���Mo�"��9>��q ?���*~���8����f%����Uqą������4Aw(��P%��3�.ʁ���W�ec��P6X�>c��$+��r�6�,70'��IF��r�8T�D.l�{-�4:�(b(�$���~@5��ރi�PO��$����|�$h�����)/D�kM"�=�?6>-�(��.�h)���>H�Z���ȡC2�lp�n��:����`�����ߒ����i[��֠"�X ��Ѝ��� 1A�����}�=,�^�>4��ABS�c�Q�0	�b�xL�k���"�V"���g�.��4T�����=�i��`i��Ȟ-��#�B&��,[j��H��P�q&�����k�y&B���;*��pfK�#���3�)�~�I32�H(��q��l�B�������ϜJ���vq6F�E���8ʝL2�\wzB�-(��YIq�4A��4ס�ES|	�@��a�.�OIz�˼��� ����Ss�r����}~�k�M�撁�lbM�=�H�=r�[�\Eao�<W�ç$�Õ���9q������
ݍ�R�u�e�P�È!)(�`y~��+��R�٘݁sṉĳ���y���:MU8��}ߧBN����~�7���},z��!D��^��.r���/��\���.Ꭱ`	U�i�a'0�w�r�)w����?��mZ�gΞg���+d{g��\;��w���r��(+�l�ǻ�q�am����9�veM�12��К#��jy�z�`���.�z����9h:i*TN8����%�e����<p�(E����s���\��bww����a>����}�}���'y�n����˪>��~��L�k���s��
�l@T��e���4~Cz*����H�4I Ñ����ӀOI虐�R��J#(�4(p��(�q�3?�P�6j�:�Li�1���(�Q/��d�%xa(����f�es+ԭ7dqiE�=&���^���j@�ҔMu4j��P�$һ��4�,�7G/1�w����N�M>�P�*�V��c�u�J������fQ�����r%����O�"�u�s%T�6Fyԓ��ؔ8���"*IG���D�n�W\��w�8�s)�3�a׶獃�`��֬6.��8���F�hWf��e�Do6Y�3lo���6'���Ӳ��0>5��vDG �s���ڧZ�_$�)v��!���@`qz)�1��V]Y;H��H(�G�8��¤�yE컬���W��{=�����y�^�܉j�x�����:���Сx؟82PH�	j*ۯ��pˆQ ��a�d�����	{��dB�'�C�@r����W�Ln��Y�p�����u[��#��B�x �pP�Ǐ�=����n�ǎ�-pPC�M�b��n��An�V4Ta�Ըb5�cr���~�G_���0�}�~�d�k�ʴr���Ry�7���ƾ�@q[�yr����̠8�����������>�;JJp-4w@c�sx�>����O�u�nǹQ�����c�Q�5�r6pX#��|�%35�G6��u�X������S�6�J?!��;�A~�[�(�c��*�B��E��IlL$V�Vn��o�[S"��r�w�v��p�Æ����� b���3��4�l^��Q�%��,~�2 �-��`���/[k�j�u�y/x�<��rם�˱�7J���wS����5��]h��)��vO�8>�a$+j =��?���=®���E�O�β1˵�����vL/r�Ǽa�蔳ȇ�!���"N���-���e��ę7�]�˗ot<UY�UP�YOuD½}��_��3*��!�_�ΗGy�]ϖy�������^+�WK�nCd׍�BT�h�܉+*���tk`��e��H�b<����.Zp>��8��9��T���������Ңk[-�������iS��L�6����kSZ�޺O������26;"n n��z��Z�4��*��Y�{��[�Q��sߛ'/���nn���)���:��׈���g3�=��d]����n ���F$�(�Y���`S����3dg��a��`@��߶�e4�H���B�x 
�t(�H��9N���]��I��Sʳ��.z�~��U��(k�����g�������R�!�3V!���<��<|�^���5��;2� s�s3�R��df�&�}�?�J�Bu;;���ú�@���U2e�uua���q �~�u�ˋ�����(S9��ƽBa�gZ��!U�h0����X�x?Ix2>�͌����\sJ���/����ij�k�u=2/��K���5Ը����VO�}�y��>��J�u��{����!C�ۺt�w�y����h`����4��k�$�X�_NY���o^z����I�����<L�|�MZ��AS)�	P�K�9.Ͽ����	�zdZN?qVZ;�����n��km|f�����V�7����e��������qAc�D#q�S�]�[� ��N�q�C����09�4(S�G4BT���)q>Eٴ+��
�_pE���`�]����}�|9���GN�b��aS&Oq���8��}�9H"�f�A/|�����z��<�T$�
9x���p��Z�D��`��ϙqG�?e�T��w�[}�#����bцy@t�iQ�@�(̴{�y�bNca��!���5(�"���;6�{��yv���9��%T�g�W�� ���H��ʽ��	�aw?�*u��-�������+t�/u����F��,|]���I��Ld}B�� �9.bx��xd��6�"�g���#�:��z(��3��?�w������1�@�e]�^��h�C]j o��c���޾�����ۣ����	p �C-9�=5ݔ�͋�� :W�ap��$^�v�<�ֆѭ�����W��w�����k?}�4;ݡ���7�͝z����RqlUžѬ�����~��	*D00��4'���>���!��Y)�,z�[�Q\�� [)��9X��^GD�6`��SI�y|��LB~;�U~�\�Ey��cI3-R����n�޼��0({���}l�?Q4v��F�� �?����xS*�I���A>��}3r�_"Ǯ�R���̻�_��������(�z�UדLLaS�3���c������e�B�(��f� ��<�+��/#ʢ�D�ॖ\&d"��3�F�{B��"{.7^~A��;*�QR��£�]��E�o�W��3�8!�޿�=Yڅ.��q�^���a��X3��M�C��O��e�)�k	����n�M�P���S�x�4OEѨ�!���+u2&�dC�T�6�R8��Es��x�r�Y�s����մet!,(�P��X
Y�\�|	k�iYW��@M���9��fD�n�|!�@�<�d� �.8����e�w�������w9�n'2\ 濈��k���,��B9�}�cEN���{�P�Hc�a���ވ�\�����O����r�"'Q��(�i������"ؠ���0��Xz�!�|��(��E��ɼ�	y��_N��*�W�@�#���9�� #[�L�b`(ָ6��������w�T��̲{X�{��5�#�9�V�-�@Ͳ��JP�����tQ��{�+G����7ȍ7>��͇CT�w*��c#(
���������O�����	y�k_ˆ!@�����4)�w�����%����`h8Y~������ �0Q>7=џHI \�0<�z e�K[	�S5��{�B����X{�Ϟ ���l��Y�yn��Ƭ�_/w�}G.��v��詊�=3���J>��s!-��X�H`hD�y]��/|Y�&�)�:���v뒜?�(��~����-U����;��Ӂ�l����K����| ��ĕB�w���a���xg�l@\��K�s��<Ȭh��@w4���7m��R��~9�}��\�o��X�w�Ã�/����c5�)SD�"ɰ;f)[��/����W�d?��B�%�]�/���QpJ0w%ȡQbys�����V���7�n��'a̔��*3*
kr�gyg�-��n�e��v-_�-4Oa�Nh���`o�Xwo��e�ݓl�i8�C�G��¥B>w�Q��0e�+Eo�b}7�����7eem�̃ۍ�ϯsy_��Qw��v��bw�b�����^;X���}���ɮ���8��p�z�F�W�X#�P:��/烂p��2.��y��2=��X3��2��s��-|��s_SeyT=�ɩq_��
{ߣ�>�Mw�'���}��l%�#��FIr��X����r�7�|���o�;��z��z�$���Y�nD�L	"�bx˸&>��g���Ggc{(������r���=*�ᨯF������_}���w��򒗼��=�=�Ǿ��>������9y�|�`?�o�������я~�D1�V���~�_��#��S�4lpO���`�J��3J<�'>�'�T�+� "k�����*k�Ƕ}U�z �*����
�^�>SR��j�#�D�Qm�ni����G�U˽G�z�k���_o_fGe���\��|lj�n Y���ky	e�3R��O*V�>��Qw�H�7�e�oeU���V�����e��(�+�����:�	]�\vI��ՠ�O1�g����nY����R��*o�I�?_u���)��
/��J&3�@���*��\�B���h��]�O�.J%w��\�J`cp�.�Сt�f��Ġ�q�q�Q���^�iH=�ЖX%Uxd{j��S�dN%Ajq�|DN �f��B�)K	�u]c�,��	I����&AG>��y�;/Y�0�ճ��	%�C]�U]��Z�yB��"8O+(��W��z(nȜ�{s>�^F�:�',#�� ��"�ۥ�C���Q�c�nh�p�n<(��Q3��s��F�cSH~}���{cA(W3JA�g�õ��Hp���>�|Ǳ8�P,�ݍ�8h��
��몴�P��QOu��] ��� �kie��v�l��7R���}V�M�T)ص�2����ޖ�����z[��UC	��}�������̍CA	ó�½�λ����#��?����Ǩ����w��k�&�_-{}�ٟ}�m8ݓǜ�m)�	�:�����=(���Sr�W�g������h9�ȵ'�-�@���ɴO@��*5�\ߔw��;پ��~�b�;���,���?&�S����9z�q������o&�U������ߗ�}����T�gnf�z.5KI�S��1_�+��3��U$X����!��3f�!M���BN@�^�E�.M{����
�)��Q��8��U�4�C�hSY�eF"���څ��Mz,�@�uV�G%y����*�j졼���Hs���}�R��'h��
[���#W2Ú�JvE+R��ݠK�ˊ�"u�a���rv�N�Xc��r�X�����'Ǥ3PȎ:V�k�15EY�M|�c��7�5�]���<�ʁU�قj������#D�X(YE�@L��.���7�4,�ɑ����ی�Kt�-轌z�O��?�(VF)5��dO���2��:�;�)�r'��1�v�ݘKB�c����kX�����ب��8�F��ӁT֨<���^����\��vo��\��H?�"\���reJe�S�Ӌ*�6/-I�f�dyeI׻H[�W9�i��ñ��9C�`�J�5��++�?j�)''��eK�Ą�Wڌ��@���Fq�F�~�R�A�&�vUJ�j��gc8�IT�U��~oT�\?��&ɾ����P�S��OlRL>{���D�: ��<i	a��+��C�ޓ�jN�⹒�ao��"���v[�~mϱ{I���~׶�Z9S��p�������.�r�-��ލ�������Yω�B��^7 �����{����l��pIZ�G6��'�n_�*x��������&�8,�o����nB�冒�A�
��<�z����_�b����]�Ї>$���F^����>0F%�wQx����N?��G>���|�w7&��a�ܴ����)�*l���Cz������z�!c�ld=��lH�t�#�с�������9>�яQq����-z�W�|�����|�S�����|F��;��	�����{��^�N�0��ϟ�q��z����0�iD�����E���Z&����.Ԯ������l<��(�@�
2�A|�����3�K�.	�RB��^i�����>�šo(k����G���0��>���g��F�d�(������*bX������s���; ˽ 	��q
��~d�K��G�wm#�~bP(x�iI�_�o�jv����v��CУ_��u`� t��Q���*
�Z[�X��������6�����8���S�h��(�d��uw�i�(����'��ۺ����Ao%��m��2��=�O<ř�Q[^;5��P:%y*��^Өi$�7�qԐlԍl���UP���j �x�}A&�I�}: �s���Aw��}sD~��=je�/�3���/���M:,pd _�D�C��>Ay�Td�>��4����x9b$�ɽ�I��Ȝ�X��<�Уr�����)��kRN#�9;��`�1�v���Z�vzb���x�|ffz����Kj�V�7w�ll���]�o�\=L�����\ks�� �[����ؘ����z�%���z�üS��"׹{�,ي+��ny�ݺ;a��K;tK˕{b�s�F��I��!u��;���ƽF&��8�B��C�c��fy���Q\��@S�{���2n�?�0� ����i�l�&0��+������KuZ�i�������~�{�����z:RE�$_����y��S>��O�W�W>��RI����3r��a5(V�~��~�x���W����;��c����촜;{�
��Pk+�2��.6U��T|�2*_�0�$���٬�,J%K�ӆ�p������?�c?�h����|�\��T�(/��1V���ɟ��P~E�:˼z����>���ϰ��NV��.s���I %���u�q9������4�@3_���Rn�V�������r��ޣhd���k���؉`��g����2BC��Uٻz�́�@c)�v.z�~�!�o?f%uR������Ha���w�ʰq,�0{�F�(	��p~0w��H̐gʦ���>�l�c��Q�\�S[�j�
��$M�O0�,	�G���L����<��c�\�u��#�R��]oRb��2�vފ�TøX+����t� Z��EN�:)�X���uxH�4�/�[!řq����iX�ev���*$W���0c�9�<�^�G�����j���`7?bC"�i�L��cU� H��A����ẂR���5W[ۛr�ú��yO��Q0$@�����򦨍U0Oe"v3��yk�?43jxھ5����۷_&&cYZ@{���\{ݼ|�ß������מ�-.]hWdt���q��#�����/}��k�;����o������qG���;w�}���{��Z��r['�f'&.��13�������(��iQ�%��˅���]�����'&�=碇^��Ñ����*x���<-c�2��Z��E�=�~΂���O���n@���s��EN�/U* H5�u������6�֞8x�q���|&�f�@OP.��PP��ox;��^�~za�5<���Oʖ�FȜ��:>�=���ൾ��7�Y�zD�C(�����!��۽D��q���/�u��a�	�(���y�t�a1���h�^�r�w���������/�����#��Zq'3�\�y~��~��1��@�zǹ[;]iN6e��y
8�3�����uzdt��\ϻ@b6)<U0���*�dh�����ߜ�f�N�~�*�I�P�P�h�^";R�����D�(A$����T����S�oKQ�^������/����$�w�WfFg�5�Q�Qؗc�m��1W�O�쵚�z�� ��Z�l]�f��{��p��ַ��c�Q��7��|P�ۭ�	���K2��%�mF��<��̙�Ja�����e)���t� V�w�����-F����(��#����R��s?���ر+dg��2L�MI�\h��d+)��uH��6d^�L+b��!\�?̝F�
�������@c��y����*�Qf��pRU���;�l���^D���5���Q�h�=&1{�������bP�Q�" R���������<瞙�+���������.�;s��s�9o{���gzei?����9ە�1���6
!S�H{�*J��??�ǂ�K�JyޖFS�� ���NSYΖ�8��3��+�86��fH?ׅ2�ɤ����CW�c����m�������HpUS}˿��g��'_|��+�9����"�;��<9||m��o���}��E-:3���^P���$uN�
DY^ �u�c��}Y�~p+U��/ho/��~Yv-k̭wEs�����w�w���(��!�p�(˘��h"w�`G�Y��G�Nj�)3��fd�2N*���uE ����m`�C�{�&��FY'��w�����!R���T�ÏZTl2Dz2%�c�D(Ny�o��q�s���<v0҄X��H2!8V^�_]�1<��5��{�aF5odT�ޅ�	"l���z*�G������T����wS�nG�.�m���{n` `lpM��JX�������5��e��qb��Y�ދ�K�1���������7ȥ�^�{�ܹs�Y�׀��Ȓ%K䡇b�B+���I�2e�L�i"��!���=�l�6��_w���ׯXg;y죑�3'�Ζ]7�	f:��Y��`�,(j����P���]3FS<k��	�����{�P��n�B5E#��!"��F��'�r�o;��t�}��'���Y�9� �;A��cG��=d����>󬥩ى�M�1K�;pP�o�~�6��E�l���oz<S�nAL��9R���mj뵴8ڊv�H�w�;e[]=�Щk�q�\�C�k���f�;�)[���!� G	�__� ~��d"C�j �x�ײqs-�YkK#�+Y��8�B4ȹA���3[���4F�!h�#
�c��F�9�d¼OǼG�� Z<�R�����UU�|��Gs�1Pz�u���J�t�A��׏�)S����&�OoZ4M��JrW��� '����(ZH�����3Y�|G��-��kʩ<Oܟ�@�>��dWR*��ƭ��p-(.�`gOwlu2�x��Î����n���c�z�r噵/ϝ��3�������D����x�� Ȍ��C�5]�X�(b���j��6��56�w���0w}�]�vG�'����- c�)��t�M�Z���5��m�ܦg݀���]{9N�@�1�}������2�P����GT�f���q��v����¸�6�H�F|����HY!-�I'žǜύ~�M��p������f
�kuc|�ĝ�����M�>�)y���/�����B�5j�o��PGG�,j�Օ9��m�i6����?��R3�q,M�+�Ʒ�sMO��T��^y��7Ec`�D) Q�'�|B����?��Y<gd"�M�F@��ŋY*@K�	���W^�E���='q�8��#�h��#�N����!B"��Uv�d��Sk�|g�ĺ���RD���7u�!ӝ�����P,E�A2�m��� 7j��5��KRgC�	���A�<PY4�$��q��{��7ѺΚ4B=�|$nk�gJ�q��e���k �w���JP��@�9�ȴ���5e#k�?0�-�M,����WL��y�L�	^[VV.����<�=oX�LEe��Y�Z�ӆ4;6�`D����7p0��6q��6иϛ��9F��5kW����׀�`w".Qt/��`)�aԌ��I�`���A����p!҂{͆��)q��Q�����P�ZL ׏�d�Rо@��c�O�������R�(k2�-�"�3j�E����`;nIۍM�f��C�5�0���Ca�N���$j�V�Ђ7�É�y��R+�ejT��(���eD��@�N5Ȑf`�3@��x�΍b>{&�6�QL�3�}yذa�H���>�D ���ֱm�s���[������O<��wf���F�8N>���O?ݴ�����y_��d�%���u�<8��t�=;(B�(��1��I��:������n�5l�����
��{M��#ye�}���m��5��,1��,���ޤB�9�\*�Re��~��|C���Ddz��}}T�q�y���eAn�<wT����(�d��^��!�X��g���8��E��L#�H���jY�WN�z���ܘ����b!�~�~�Ǻd�ҥ�4��~���=w�M�8��������� ��_|QN:�DF�˖-sdQ���Fԋ��~��G�:r4;Q5^���<�ߛ�}�����c���]����Q�&Q�<�q@�8j����]C��g�#���~����/�����6dp�p\�o �Ps���dժU�h� َ:0�V��f���q<(�!�ȹݷ�Օrwpj���1�N�ּ�k��P�͝�3S���46������|Gۙ�凙6*��[��۝H2\��(�*�s?ѝ&���ȃ�L-V����h���f��#��b$ww��dSD%FN�=p"�>�0)�u � �W�I_x�yn��<�"����~ �<E���'�p�:���p8$'q�444�A �PTL@��}���A��Oj��l�u�K3_�ٳ�e�6��dO���H3ݞN���WJ�Ф�7��(p ��.��!&�z���aJ��'�K�l2:X�����g�����T�G�geK��d�d��BǍ�(�u�.�8>��]B�Z�d�I{�Qꬾ��:5:�]r�����s��M��X�:���9s��*5��jTO?�4R@/^���G��Eg����-�=;�R��t��I9�Ѓeo5�H�?�χ�����^{�i?=����D�S�^��HA	�#�����Aiy�\r�E�~���_KH��w�t�+*��K.�A���K/�"o��&��(#���JIqAGsS�7�M����_��;��_�g/��^~b鷛jҾ�O��2i�O���P� ��ߔiI�Q���N���es�I_YR7`Τ�3��tw��w�@ݠ9���8lZ�����2s/�\�o�m�â$y>ooD��=��֟��P�u��I��v��;;���[�[2��B��`<��4N�]����О&Z7�"씩��:��q4�K7J�y0ض�m�V~h�FB4�.d+6#Բ��׿ʸqc�SN��"˃:�F�e�ugx�V\7P� �-_��c:|�p֜�7���ΐ�7��5Z]qL�θQ{��Q�Fo�qp|N� )�C9�����ϟ1���0�scs�9�x�n(Gq��k���Q�	'����t�Mt ��{����g߽پ��h��J���jK/6��g��<+>���Wۢ�Xu�,�ii4���&�ʴ����#�a���t����	
2��%Fˆ��:�2���x����f
IZ� �G�IF��#��g����2��@Yq֏���L
>k�`����u�g�,yA3v��}�����d9�bB#t<���Gn��^u00kr���ԩS�=��b�
:�(�`�G�q�Yg�/� �Ǎ�;�C`Q��\��o+߬^��}�F}�=v�_��W�O#���63V$��,��|	����"�͛ku�Hn���s!� �y�9:.`�k�FNx������6o��V� L���
| �e<:>�@�`�i�CA��=�\I����Za*# �uBD��>�c��~�I?��;D>xo����J��C�u�<��R��� �̣s���j�J'#듩g�Ό˪��y�M�60����ڥK��S�#I�{�[v�u5���n{�*>�w9��g2�q�ͷ�Q^�v��1�gRT\.��9K�f}���(��(����7��Z�y����X/'�x��=���%˖r͏9�����-(�q��D��ee����y+��yY���O?�햿?�p�֦�k�;F�BE� p}���'���M�-��Bp�EYpؖ�n<��^F�n�8,2آ���ꋜ��M�ߘ����%T�Yd^
zt�h^7
�$$� 5�Q6oGT��,��i"�|h[�l��M㽈H-> 瀗�סvĥ�'��6�i��稬*g�mkS�zK��VP'�F��/���`���L����'@�ZUD����a���d+R���[��\y�U�v�j�0�����4_EE�n�7�{G�Q-�:�Y�����{Na�<|����,!Rq0�@���x�!��o4\�ͪ��n�SD�UUe\�o���V�{�1�8�AX3���F�6�G}�}� ġ, ����gn�����>�ʊ~L���KxVpl���r5�8�7߬���Ngr�E��>�p�V�,i��aN�n8��ύD��&p��5F�1hw9F�q��+���߫� ����&F���.�'��a����jX�4j=)� L1Kd~c(~#&����c�ñ`fy�:n��u9���lX�zj��P�A��R}�����GR���R���(��`�����Jy�Ǹ.>�h`G��L��?��ر�%Eq� ������Snh�&��yMft|�J��t�by���%����ك��/Ȧ�[�QXX�(�-��u�ḷ����W�������:��ӎ�7�(>R��v3���9\\JU3� ��)UԜG��}E,>�Gp���][l	++�S�1�6�?�Rџ��g����ߤ�"�`��~���''q���dʞ��)?>Y�}g�|�Q9z�̟'�j���:�{����GT������g�^x�))�}N�{�Nξr�o~-������0^�y�)��OO#aU[s��{�Y���,�������0��q�9�H�C:գF׵��|�������䕗_���"Y��r�4eO�����䣏e��N�'�z�m�Ao�	��dbۄq�ޟ:���/GqP��_.��a��}t<�<A�_/=�`�]�i��3��;��}�(�w
�,e�����A7��>�y�p;n�������He�t�pG{6K`k�6�����;Z�)n����38ȫ�ˣD�sݶ�uI��)Oc�}����`�3�u���D6l�) j�����Ė�!���>��V<h�.��*��¢���2%�T4�@��8�?jԹ�6�����˘j��.8x��^{-#pm�n�>v�x�����1A{��
���3�#D�0�����u[d�����`�lOlMM�l�:��s��j�8"0���Qܩ����9��&M�Dc���������yٌ�<�����s`C����#�WFT��=�}��NI�<��`^!��t�1�H^�C��3�����io���q�<�X�\6o�N�bFf��E���:��ϗ0,i�!{�x�(cy�A1�sPS�L�I��4q�qyĽ92N �����۴��n���SF��hƤ�A����F!�}>T�#�9D�܏X�c���_H�l�(R�S��[^y�5)�(��O����D�
�Q���������5n��y����ϡV���ur�I'��aͺE
A� �q3��m�y�|+4��y��Y$7�w߽e�K��;>P��Ka��M��r��_�Ҕ@CG��2�!��1R��1�Р��s��z8IԽ���~�QN��?K��B����C�`i��Ur���bu|�Z�lC�X�l	�H���gvذ!t0�x��d������d�ɓ���JiE)3r�z4j8/!k��*�*������s=��#Ҫc8t�H�z�2>#�'���+4@�Z�Mj�FN���(���:l���\�g^p��/#��@��Jć}[�+0��D�'�eʔ=ֿ�����:�=���;��fk[}swv�e�7���#P��<4�a�J[���/���u&M>B��;�n{�=ӞekP�g�û���w\�K�;w_��,ؾ`w��ll��Ѱ���d�:�헵�u֦�t�ub��`V�S�wv�lK`~6���"7�� �[<�d~���?�,2����hJm���o�J�~ՒUG��Ġ�a�,��'� �`2D�0hwݕ���_~5ǐgk �!��ܮ�O������e�FW0��^ >��]�δ�i�׹`�B��f,S����_r=#��>�\��{:_}����H�����6m�H�xL_��˶���
޿r��n� �x�4�����eox?.:az80\x1�]�3Y�4�!P�n$]B�.(�A�0}���KƩ�2AM6�I� ��Hv3�2�E��r6h�LѱX6o![�R����S��t*j�ޤ���ӛ&��,F�H����Ey��,��jQ#sY�D��սN ��o3�:/��JwW:�h
�SҭNlee�\z��dR1�`+|��j�r�����W�x��5��P�T�����������u^D�$I*)�����:)(,!Cc��L
����SN�7gϒ�3^������f3�|��iU�_��`�ԑ%���AM{�]<��Sq��F&�������(Xe.�ZC��s���S���en������;�wu��t�p�2�$�>:���  �߲I~��.���uk���=<��c2{�O���U߮f��7b�h�m�It�}��d�g����4��G�W��M2N���j���m-<�`�ڜ<e�a�+��m �N:D�v�=F>��3�w��|hЁ�2�����R��{oh�H��H*���o�s�=W���ղb�jihjֹ�d;�#���n �e�Sb�_>Ə��ђU��m�5�ն�����e�K~'zu���!9�4K������6Rw��w���ջ��F��~���]���on��܎�=_����^�m��=�0&8�2f�3ȯ�< @� ��t�_B$������V eI#�� Zu'�h=�|yH�"��p²m�:2b�t�4X4y�nR��~�D
�^�9<6AD�@�"rE䉯��Wҹ�<<w��i�
��~�? ��x�hma�s�p��fC��ŏ��	�Ø3R.5��Yǹ���G���_�\��>�1c���re[� �[(�3ܘ��;�<�C��#�F�������d���D50�o0��i���Z����΢�~#L���dL�:�gY���>8r襵] ��:�=Y#B�v�|S���x���De�F3ǟ|#D� A�`�?�T���y^����<ב2���]x�&�'�5�m։��+�;��ϫ��=F2�s��9/�e�="���� ]lUB{��ԣS1�b:�~��ߩ#i�|18^%�5o�6`k|Ai�q�jD_P\"�׬%6��O~r�̜��,[�B�ԍ�9���wߕ�|z  ��d�a2j�N�֬���k����/��Z��[	!���7Z�`H�lR㺷5T>�;D�=��0�he)n� �cF�g��b�א�Ę��L�6<Y�h�@2�k.��G��Q2��o�喪�<)/�bMz��`�kkm��!�d�ر�TH�!K$�g�l�:����I��Z��-��-�>��K/����{���YM�]*����I���&�Ю�hE�Ԫ�~�a�H\�C*�����m�q;�B*�r��p�`�v�m���[��،�e�{u���k�d�ٳ6ok�:u�{t��(k����-�r�����O>)S��SV�����J*�y�a"�;]ـ'�+���-�壨�<�?������Զ��g����l&���w����Ţ�-W�=�;�a{��^��m  ���a{=ݹk��Ht���)b��B��_�g<���]
�����10�V�ގ���|�~�9�c������X���!�<'��=*��я9�.v�;P{G��x@u�<����XWs#��;rϑr�E�4� �F�FF�/R�4Pj a��h��D
Q�'`��(��e�z�0F��N�����@E;_���?�����S�;린Nߋq�
h�ɑ	YD:Ə�s�����N�/^�{�{p�_����`<�T��@���'�X��c�6\v��Ӕ�
�����#e���L)j�ꔅ<�S&��0Q�C?�F��7�e���fS�e�z�Pg���� ��m[�_�*�醋3(�A����P��3��<����e�!iqk��z�Q�K;�#.3��ݢ'��I�ߙ�j�65\��A�5"�3�<m�o�h�DAuN*);k��l5���'�l�s��r�Yg��~w#Y��~�u�ɲ�v�,X�D�U ���7ˑ��� 3u��y���PuF7ޓa����g������+5:}��b,"��p��pcMG���:���~wgB
u����d�\�٣�ڴ�9�D'fO;,~0� <f�A��f��	1N�7'}k!~���:�yO������üGA<o�4�C��wd���v�qG�ĉ��rx�:�'�gV郏?��{�+Gq��3^�Y2i�޲r����'�ʚ�d��˄]v��3gJ��T2-�:6q)��O~3�:���2A��ig�%>��t�ar�ԓ䡇���C��ig�%���X^z�Y�Ӯr��˟�i_�Q>��Ǝ�X�!��_Sb�D�K��C���IGo��A-*��7Ȍ���/�?���3[u/Ž�1�=e�����������	�_�����9��/�c�^�G>��]�eF�i��6R�a�]�#`��"��uTr���$�(�]˷��{}����m���͊�X��;%������n?��o�u|G�5�u�->�� !�p��0�Hkz4�J�t��Y�g?�"q��vl�|Μ9��.;�>�x�R2<�������k�a��#����!���u��aL����N�4��~o��Z�c4�������` W�g?�C�G]h{���t�4f �[�Q.ڕ�O�}?��q�����e��8/6�~��Y� �[n��-!RsK���1�/�pD>���\��&�dc���hQ�]���<�@��u}��~^�g��st��� ��ѧ��7�|:F��.�r���ҋ���� y�!ioh��+�FmP��ńk�>3����7uZJSfM�7m벮��m�3�����'��>,��2�)�kЉ쇣�3�p @j�,-�����۪��F���@$H��X&�'����䱧�P��Vv�i�<�ȳ�ƛ�į�q^��Q��&uJd��gdU��#�;~�<�䳼���5̺@F�=��#G��A���C2���Ǟ1������dOt��p������
�hi"W�E$~a9���XL�L�0,QP�+��A}|т��P'�f������gV�4�d�@F�bU+Y��O� �B �s	����
����E3���o�5W_&{N):@2t�P>j�\z��D����l9���[5��n�Cv�8Z^|�m�􋅲�Y��"�^p��W�>p� ��?2}�<H�j���_�s(g�;U��?�����䅗^��3����Y��s�a��b�p�\Tc�k�չ]��ٖ�9�G���D��\t��RRX�iv�eWȵӮ��/Δr
���ѕqh���J3��w��9����N���L8n>�42$b��0b�~l�s6E���%����82+l����?wj��Y�KI����i}�z����o����ǗE.�,�;�&����5�M��>x7m���Fȍ��5���9C�`X��T���̳a}m/����H�R���)�oo!�um��p�M��avg-
�V�δ� :�"-� "CD:H7��O�rcD��r�� b���Ĥ����4�����Qȳ�/2�f����m:�F��{�_h��^;z���5�[��1ئ�o����
������q�k����1+$c�(E�8K�sG�M�[:R(u�e�Z 1�c����2g�t6F�+��<�ׁ��js ���L7�l*ìC�^�9����%��	P��w��}��ܸ^���,�d�N��4;ڰz�H���������A����p�����϶7�ko�Hک��6覮����a�S	�Y�4�����kE�'�����l�5�|��'e���щ�����E((���z�*����e��5�ڈ<��S�XZ&��w���$��Q.����K�:�⺤��J�X�X���6Ss����)�g�,G�6��~^�e�2��Q�I�BEM9A��	s���$��cM�5Z�~����-~3��<6�k�:Ĵ5z@�N���>�6i��5ۑ�ɚ׿��9Rӯ��s��w���T���V:y��U���r�]������5�s1j�F�	�3Y���5k��,[�u;j�8٢s��76���:��OV#����3^�%O����̮���2�gSՙ+���|T,�n��o���S�d��I �ο��-R�b ,eղas�:t>=~g���O�W��5At��յ��F���=%�:lm�_<��M��Tw$�����eAP�= ��z(�X�3j��������L�s*�
Ez���9�Ծ��}��F��k�!�iM{n��|JߠqI�M��T����M%	>
�/�C��jg�̆M�P�R�>c�#ܔ�� M�_n�k�=ش��A��r�iKJ�1,)*aj�9Dψ��Vg���t��
_FE�n�0���k7��{�v��G��������nFJE��c��ދ�������;묟˼O?c�������mns����ugk`4PR�:�t�|[���ϕ`,� �	-&��f�ѩpZ� �Av��#�#�<BN8�x�ݼQJ��dS����g�L��!�����aÆ���w:��y� i��p��c Pph ��V �ׇ��}��_�{�}�\`⬧��]��Q��v&��Doih&�ϳ���c�r�r9��C��	V�u�n�~ wZ[�e$GS�F_1@Y/�����w}^Ņ�8G������p fL�!_H|�����R/k�X�Q���l�T'!m�V�R��A!�>�gӽN��R�2����8�h���9�]'�!F��;ׇΝ"�`��D��J�U�,�ڢ�
)W����Cb])))��0*1���-�d��+�N�}(��k��ӅT��`kS�dѽ���[�}�E}Eң����l��:�k���j�rk�nS��QL�Ԕ&�C݅����6SR,��ǽu��-&��(�Ad��g q�0�>�bg����4��=�a�T�(�XW��uO�gL�I����f�\�L�XKII�0��MZb�rϟ��6A��U�W��hW<�k�;��?�E�:�!]���|���7��{~��_ym�<��'���+-.Rܦ�q�<���'�V����ț��ҁ�=�N�X?���ʇ���';��{�P�u����(=�c:���	i4�ч���s?�bu���ZL�0� �2l�,]�B-�Z��0f@6�ޮ봰 ꋵ��[���H��ǶƦ�Tw���,�����]#�p2����⒩���6�8w&��uc�}�U��QJ2)S�)9C�Hf^����q.�_[Ͽ���G���&h����t�������|Q��RE��gb��&k^f(����@���w��$�s��F0@%�y嶼3�/`6�iT<9� j�	����&����g�KӒ%���1�:O:�M��s:N�X"������@��F�=���w��r�M7Ё@��A$�׼��V��2n�ŵ���GMu���	�ȵ���\v��2�� ~_n@r1�[EH��@$D+��.FUW^uk�Ӯ���E-���Cf�H�d��kzG��.���zW]�O>��C�喛Hn��3O��7L�U�|+a5J%e�l�����QMU�J�v%���V�^bl2Pm�*�� �R[{��M ����&�Yj7����"{O�K��e�����
J	7��������!�hK�p���V��'k�]��fWAXо�̛�@Juc� J���*����`�C�"��x�����:з�}"�*7>�7����[n���֩�+�Ts��'K�*\L:�GBVB��$�Z']�M�����Wrcg�6T(]��!77�m��6�Y�4�lXK�H��*�FL�ާΪ��y}N@��HR����Ji�Z�N���U�q��UT�k���a�:,@:��y��������AC���4�ެsy�n��<�F�&T����DJ*�u!�Lu.�H���W�]*]:;!���ް���F�^uN�:�A�B���a�aR�7�]g���+L��'e�����`�c*ݫߓ	f�,��$=�i���_"q��H���`(̮	��?�$�0C�3�,K�d�@:����HޓH�$��9ZQN	��U���<Bb���tJ��\��T�h����)�p��aXub�0�*�d�<a�:�%���C#��v��{}i��_#�f���q��o���9t�@��G�eL�qay��}ku��	S�����,J���i�9ZQg�OHAG�*I�}����z�Q�0��uL�d����ߟ����ҁ�>�x����/��W����x<U$���B7���j[ScT��gړB��pn�N�g{�ړS����Fޗ��}�5����4}���!nɥ��!���>�Xʛk/�.2<dl�ԩsn��=����Ms���I���r�3�w�fS3�[�g"S�5��A?��b�ͩk��0��0L�mm7�<X��K
"�,{s��3�=�4iw���M���k�q�T���n��~�pc�Q�b��v���/��?��n�~8��x7����6����Q�*��csGE���)źm�V�s�8V|��4a������g͈��!�ȫ�����7\�|���<Ƕz�U@d�g��*��6��u�xQLڔJԘ��q��򫯘�?��|o�,]Pg9� �H��E�e�77.�<�j��zG��c�<k�3��NP�u�޻P�XDiPv"S�I�2`F;���d���������<��}Wu�tc��hT�1��T6�tc���w��d�}'��]���E_O�ܸY�@f�Ջ��w��9��sM�w�m�^�~3i�����cB��$�@��2k��e����ܡ�m�9ɔ�lА���~�}�Ο�[��ya,��pO�I'4�nVgF�+�!�Ǎ3)��8|${�A~��c��e�.�����tT���1���t��x�P�z�"u(p:�������ac�n}o�f˲���aj�8��^��?`���7$\Ee%zݭRVZ��^�*թqد��.R47�k��^bS��-�i�|�T�q/�}�C0%� `PhFHB�#e1e �hPn� �G\I�|�u��d��<��b5����螨΅W�2��Uj�;���s��SZZ&�j��!/ "�'�_�$�jТ-,e@��
�6��S��3�W���vqY)� ��fu�%m�N#�{ZZ?#Z��K���BRX�D�!C{iHK�w���Á����$�@��7�j~�˕�N�c��/.�|ؚ�������=Ǟ��H��v�A�����ꐈ��ir˛�1I�^ui���l����K��?o伮׺��v~�?�S���~xm���0�J\�59IB�׸m=���a�n��칿�qX�T˰�@.u]\���L�� T����C�5��Ajq�34b���$�F�t!�魠0*w�u��0��;�s;�H�b�������;��3�z���Q{���Y��Ѯ���vҸ��5ꨙ�v�T���j���b��㏍�;i(I0��O V4��x�ٌO
�Y��|?7D^y�5fUn��zy�ɧ��{�,3_|Y*�cǵcOu�["4���E�PpD�5۷P6�J�05jta��cwb���$������@jӶV���a�s�ϑ��Q�+Ug�w{��t�I$6��8f�8:[����UG ��N?�
��!��zo�9_�]A�!�´i���:嫯1�P6���Lz~5� 2N����y+�c�;T.<�XHx�?~N���5iڰM1!*�:'�A��\�2If�Y�ȕ��P�z��ws�� ��S�<��:�h�J���J�0v�P,�W�ʇ�&O<7C/>���1��*kI���5``�x��hO:�x�y®,u���aj�L9	z̾ӣ�Z�4�q�lH[T���vҫ�������1����d1�z:w7��͋��,�������9�ੜn�2RH�wBd$���F�muL]CڴA8X�CZZ�!�^*R��a ������	�3j�S�ެwO���� ��Ҡ#��28=��(/����t��B���%���5y(���`D␡��za^0t&�y�D'�3�[}}�-����'��\�p&���֘^O��tk��6����2] ԣc◵�7K�S��qTG�M�YF�"ץ�lS����h������0&�r4�d:hpˁ!��::e-�-?z�ٗ����_�7�\]��[�Е����1�t9y�D���C'v:���&��HFr��֘�������pw�ǭ���澵w����Àz~�h������fzޥ����{���]
�9-�m���?�k�[ ����k�"���l��a#l����9f��\��^�"���?��N��),�҈����r�6u��h`�R�5@1lr�u��hc��P����͵�L��������U� 5	(P�"a�ڍ�6|��	�d�(�5]��Ef��fs�@7�
�ՓO>E��+��R.��9考����&�#2����B�"�XOeE5��[cc)x���d Ep��1�e�^�e��q�W��g��>��B⢍S�7�i!�id5���KiE%3 ���������F�|���2d��+�(�l@���;t�(!u�T�~@e�!�ٺy���ګ��D�6��U'�U~�!8d�� E�Fp|�t�AX]
#A�k�z�M��Ň���	r�1����NU��Y��[���H�˩��]��dK;<h���s|ǘ�����r����6ȴ0���H@��f;��̘����n��w�]�=�T�G��ᇟF���'���1���H�:��=v���ote��FαO�"G}��t��u��!Q�� �	�5"RE$��u�H���
��%���1K���k���2��1G���1\L���5cbk<���D�$�Hd�]���}��F<l�^c�����ioC�3�C�<x�re���DB�AJ2K�:�@L�L���FH��z�NzW[�lٴ�%=p෴4IY)�Y����Y7Q�?��)�>�0J�,�~
���tQ���,i��>Z̐� �$)0{��802�E�Υ��'���V�GeĞ�d�׫���Fj��K@�=����x�m�eYS��ծ����M�:C݉�^A�+���Ay���ɵG�����w�|z�j����B����������+Wm8^<	�:e�̘�K���2�q���ԫ�,#�=_� ��q^�<,D)Ӄ�uX�
[_c�נ������美������w~ z�<��� �Au6r��m��~�}����}���/ڟ+M��)��a���� Q�-g�-	�ϴ��G���c�9�BD�g�CR��G#���"����p@|��������������mT�B*�]�cC�F<�NA�q�[P$ q[�n��R�`Q�Q9��{�t��5�)O3�O�('�"�u�@�8H�F?�a��nnj�̫*kx�/�-��n���h����(e	n���Υ!nkk!��"ؓ�$� asJ�����r�A�y �}�ݹ��(��;ٔ��\�!#2��P�B6��.��.���w��/��-����)'
���=gӋ�zO(�f��q�P:0��q��GcY�;n�Ӧ�&�￿�p�-��ϔ3�<C��R5r���E���K�j�tᒐD}Q��dIz�t�w��_)�v���o,7��������6�媒R�[��7��-��ʃQ�
 b�$�h�,e02~�^�$v�ʫ.�%�i4X$����:2~�yP��a��)����C g}��K�?�X))ʥ�\M���a���QƏ-/3�+d�T����,RԨ!g3I�+tޡ.��x$`R�pH�pH ��x�L�8I���[x�[���3L6�m���o:��ĵ��ɡ��X~�����I�zD�uj��|�̚��t��*,*��z�>G07���})��ك4���|�,'�L�oдa���m���Yٸz�v��RӯB�����>�ꈩ�k�fLV�]/ ��3����t�Z(���65���dۖ�g�+�����lm����%7l��A�H�۝0��X�h0"�Muk����S�d��ǝ"G}�\x��v�*�OejWBL��Q�¥:�e�ҙ��+��d��2f�p9�ܳ���:�P^������u�*�����3�����{W����w_}������X�fMɿ�|9��O��U]K׮�ҪP{k���L6&���e�����"m>���F�g2�����s����v�(}�����������j��k����=�\�8l����@��{��v_��c��3Ϧ��ÞF�cJ�F�V_�ԥ	�x7��"�H��L};ө���2�E��؈.�XG;�)lL 4j���U������.�D�;�By��Y2��9�l�R��.��(j����k{��݃j�;����pz��"�� ��a�� x{q�슏(Z���Q9��tD�Y� �qM�̍z}7�!��ҫ��s�f��W�.��Ņ�t�W4�(!j_�l	j�� �ъ��c�J�����{
<�S{��L�8X���p�(�ذi#�۪��1���l��:x�˼�>�xD˫�B���tvh���>��,���h ʂ�p�1G2}�`8��Y!���"�q�o��#O��kx�ϫQV�;A�fW,#���3�^#�쿛v��5�9g�+K�Y#��rn�i���9� ��v�5�s�ؾD��s�H�kHsg�D^ � y��]�s�B$"�sL�e�\IL_(��W��4��pB�	Ή��J}n�673�2����ޓ�cF�#�!kV��x���q��˥K��h�fT��2"�x8F
htuL��9k��[(O�g�r�6��a۳Y��9�~FJ��Y�;���FN?���/._~�\>�;[~��h�&]~ٹ2r����0ՎdT�

#�
���..��ɍu�a�B�CJ"�j�#�SC�D���m��e�Ʀ�r����GM��r�a��]w�)�-���y{�IGKcK\V�� y;�X]]���e���i�r^_?�Wj�[�.F�)�1�'ʽ��Y�*�󌬵ٳ�d�fҤCt�g���P�t�v�1ҿ�P]��IsG�:7_��M[uN�\��/����QDo��qc巿�J�;�h9��c孷>�/-��O<Q.��t����e͚-:��R�Rw�[���}��<�l�[~��K��v��ɞ< ���_���+s��r��omj�#�/*�����g��Qv̤5������A���^s�5~�W�;�w��4��kͷ�	���ðf��݌l�3⽍��k��w�ϻ��~_��\�?��F@O�F�a��F�5��S�n�so�7�N��1w4�}�S�N�r�"��׸2�l���ς����y�� �ٿ,�O/�c-�qx� m�P�]�n�w�������#�:R�9�x5�ˤ��AV�:�bAd�i:Q=7�����R���|K�	�z�2��UTVр(��m�t
�ԓL1� SZq�ڲ
�)��
m�p(J��HKo@D���v�-����+�����r{�9Y���Amk��	�S� <��=R�h}A]�[���;8�;:�R� 90�Ct�l�H3��z�Nv����o�>ZW�U��֛�innQ�grΙ�#2j�XA���wfK�:��j�'z2N�\�@xi\|>��Q�ɾz��S�~=�ۿf�,ђJwf3F9��RP�xtw�1t�~�P����4�E��ݦ}H����s��j.�dy'5:@i�M4�#��Ȗ�"���з65��S�gҝ,��b(h�+�{��G��W_!=�VÈV�0��,6tш����Qg�X��'*��~��{��?��'��C��g,5��jK��]Ft����3�:�7G��O��1#�u��� �7��Z��Qr����b��@ƴ��5J@!�)g������E�\�Z�Z.��|��������E#�29b�q�/�g_�.67HiY��sԔ6Ժg= ,��v]�]M�wD ��O$Z�שQ���!)�,q8)^p ���d9��)r�Mw���o�]w�!o���\w��e�̗��-++�a�Z'���}�ↆ������ٳ�˯{���\>��_�9�+KV����}�ϡ�x��:;[��.�w��3�0㒯VPuؠf��kl����O��^?���e�ރV5�XKcF�d���c���/̖k�����9��=���/���H0��X')��԰�t��ٳ��_������K&Oܭe�qU}���MM��Vm,_�aS�?�|�����in�(�(L$��ޖ�gXb��`�a�Ű��tu�L�h�u7�o쮏��h����}d2���������c��1��qX�5��G�����@��{�3c���s�ϸ�� 2��r��֐GA��z�Z"sq�!�8#}����X��I����e�Dп�lX�Vs�����bil�~�ÌADq�[�Q���3�i��d?������2J�"�wL����* }��4�θ�������_�!��`/+��ȕ�kd��huK�9���}�(���m�m�ۍ�)��W��Z3ރ�s��e�[���u-_�F|[�K���8dN:�D����P�ՀD�YR )X���M�p:���+Vɶ���=�Q�$]2����EJ[7)�q ؁`�ҥˤV?ϲM�k̀�,�P@-����F�����5�>�赵��$���755t���h�����i���|9���X"��L�LB��^{��E�T�L���H� k ����nv7�n�L������rן�ū։'\�g����{���j�T)g��3)��j��d��E푔Fd�F�E�R��$H@�L�{�	z�!��t�b	�K��N�? -mq��+ق���\l�p�BDpW�HA�_�O�.�&�bl��$3��9_��HJ�[j�jpÑBӹ�y��)�tO���Fq�KUE��B��w���Y- %0�4�~_n�2����à���sM�F7��02�m�<`��w���Tb�TW���l�ߢ�S#����Ր0ayD���=��C�C�2S����Liy3��3ձ\�i�i����1��t�}����n���y���=Ŀ��O�(�ܤ��[@���;���OZ���ҿ��<������w��R��nkj�A#�ȓ�=!�xx'��cwH7��󪩮��ƭ�裏�W�?��n�A����y�5r�QǨ���y�9⏖KW: ���i�*Z�ٰy�<t�Zu�u� �M��fpS�^��q;����ֹ�֥���
y��.]�q���\1��z�Wݵx���+�+���L�����?<�Ӗm{5��jk�E�w$2��h��t��� ���s_�ǌO*ѕ�=�%��ٙ�z���9�)�HUj��0^0r�h�����X�j�[�����E����~x֛/�e��n6j8����|���>��5�}�#�~����~�V�|��i�ʈ&��NQ�V�\����*P�F�Cp����_)K��3�^���.�;�%ػ�fXX\&��z����<����0����"U�'R��W��W�n�7W�i�y�GK�+�xܻ�ѝaz��~�&9j%G�I0��E��Tk�6�Ö- ����: �d+(5[4�ӓ�S� x1:
d��'���v���!����V�C;B��gyeګ���2�Ϻ�/Y�T�"0=��x���nrؑ��m�a�`D�g���,⽁��X�f*Y�9� �b�1c�R�%�r5@p>[�Ht\+uch��<gf�2��/ם`vd����8M���ܰU�<X�PO���,��Q��|��ZO*!��r�-������|"�x�r�ŗ�7�N����Ԡs0צ�&2����LR�|�R֮Z!�^r����ʲ�d�{���S��H�}6�E��Tw�B7:0��V�ㄝv��v��-#l��_S%(��k�.8�A�}Q��T���"Z�� ľ���ǰP�<���`؆�!�«���yQx�P�B�܂�L�G$�U�aLן=��b�Zt�RY1��՛���Ȭ�rF�)�$#F�o��I`I���i��/�C?��W,�$�\x��Z�H��m��X�5��LO9�Y�.���&���Q�@�cLKK
�ԟ�z���b]�1�z�)(��ԉ���}�����n`�ұ����d�	;�:"+�/����u��A��{�I[�r�CO��v��j���l���m�>��jy��g�e�9������ff�P��frX�2^a5��@@:�E�4���ά����urۭ7��g^�ʹK6l�L@`�Cv%#�.�R#�?d耷ضq��3k��Gȯ~�k�,+��?��Oiu��t^�=L���"�;�{�� �^�Ok����	�w¦m�D]��v��e1q�=V��.E��|ePD=ި`	]�ttI \�9ոU׵:*_�\�Au6���&�j���Q��0�*g�`��l}��������wk�ܿ�����:��6�>G�k��Cirw��cw]�ޟ�����������o��\�i1-��H�z�����9����n��k 1Hq�)L�=�/����Q���7N�и-�|�X��wyeY���i��g�̙\��]v�E^�m�4i�L��������'��<5V�<XI]۪�b�[0X�|��_z�7o!��&5v�h4��g�;�- ~It4�a��ZN�h���l�?k��z�Fy��eب1r�	'�W5�MuuR���Qb����u$�m���=F������`�;5*7\�I:�p0��O��13v�,_�D���IjlF3�Ƹxv�OFm���=�`��:"��fPk6�S'=?j�1���n�s.:_V�q���"�@Ɠ�����KJE)B��'�s����a����Oe��2�W��O�g�ȿ^�7����f�e��1c��0��^T���xT^|�i9����0u�N:�9�cd櫟�SjP�a�u�3����w=��^�=�\�tm�SN:R���o�w�}��#Ͼ(EU��K B//�t@�#�PX,�J"���򯿔�;TN>�h��_�I��!�AY0��;��K���d��!��k��=`�=e�I�3õ�NQ���ҁ�[P��~�>��A 2`��Zͦp�2=Z��� �.@N�"��T������n�C���Jy���ү�I�+&;M#�B�fS��z�=�Y�O�Iz�%)����)�<:D#����i�r�nX���j5|�h���W�|�Vc��98f �F���se�.��k��C��v�,�?_&W\�K�펛�gg+C�up��Yc�a� ۮ�.Y0�ίn	�-l���dcL��{��C��,JWV��Rz�.�LY1�1�`���f�\z��r�yg���XZڌ2��:!iC��G�N2/�\\P(o�����_���lfA�lPǤ�4 �=�tj����7�z� i��J4\�2;R~��Չ���J����x��u�1Y��C7�R�e-��8dcR�uJP=��߳��$��š8������� #hR������0R��D�>���o}�������ݨz{���o�a��{#��� �o}��a�k���'_G����c(p�}�o��IH�|�U�#��3M�0��7qP���j��:b�pL���:�h������@�7��9���5�H7��Θ��lި�V>21 ���xD,H�o�ۦ�y��mk��'�#������2߲�N<�H�<��kD�f�f.8�%1ѷ;�a��+��3��.=OH��"���}�5k����Ԯ�,d��uD�(����n����g4�@�1B7�V)/���F�v���$���}�eF5-�q9INfœ �f�~P�쁄"�@�+ꘁ�c�7��85b-e9cӦZ�F�q�r��u�RV^)uu����Dm8��4���n:�� #���5���ۘ2 ��O�<["��]ό_�w(��$�I����ݲM�|�q����R�v���Ug�2���D&�YR�vkT�y�U?)�g�%;��R�*uV�@��c?�7(�@���Q}^���@��X�ke�rӭw�;���ͽH�K*īs-�����G ��ϛ!���A��_�*�w&���^�Z|�aR�z�%k�^7X� ϊuFF�1cx��/5U��nͷ����W�_@4y���Ys?a�'�\��Aڒ�y��6뇻�G�|��ȴl7��d��\$��{�K(;�~�m��̱2j�u����V���_,���^�+ģJvR�4�O'ۤP�7�S~���Qd���nm�3-:����A��C/�C�{�:����ȴko�/睨�OJr�:����r�M��ܖ`v1֩ν:���Jt'�xA��l2���dN��f����Qޘ6[�RZݟ�BQ�A�gt�ĖJ��Ȱa���kW/��2BAyZ�u���jt<$����
�~"�3j<�6m�K/�X����Q#FJKs��q�z��x@�\�D6�3�1Q
�#�5ƳDu�} P̽��7錋�$�te���#U��h������}S��*� <�2d�����aЁ����.�eI�'�o�=��-7<s������ީ��������}{G��5��pk���XT�14?|^Y�����n=t�盱�������ҭ�,qTF���!�[��$��3�y�������j�D��LZZ�L� ��l� ��j�I�c3F��q��(84j�Q���?�L���c�c�$7n���F1��O�I2�N�Y�
K�B���t�SO�י��l�)�8��`F�����s�ˆ)�^赇L���"��D�d��H�������/(�5j�l�n5d9@�|˔�7X���_#?��k���f>r��!��cM @翮ydY
�N� �<3��VVQ��v�hQ���X�f�����8OjD��}���\����CEҦ�<L	WC����#��8QG�#9��_�Pl^���1U,��!� =����|�ei'I
�dwF�v߃�y�:��tzH~r�2k���駟q�� �IN���_ʔ���)g��c9����X6l����>#�|��4�w�s�P�C7�}q�u�N�����r�����!N��]w�CN8�ly�/��s�K���1�,��>���Q,�_$<�9p���O��Gy��{��Q��	[��*�}])Y��e�F6L��_^y��y����5��D;EŐ��U�%�HTRh�J9�9I��MZ�
���tւ��/83>�ҝ�ĳI�:�[�#���#֮��ߛ#�6���Pv�4Y.��26j���JmC�4�Ʃ���RZ֩��^p��TU����6�j'L�(SϾPv�m����d�ڍRPV�`)�Ư�(��cz�"�jo!a���j���Ŵ��Ev�yg~��իu,
��;N�C��[�F��f�$:h���L�n����R}MF�/�/�����{��u�8�nP~B�-���G}F�8�julq̘�U��
p̏� z�Q��1O}��֭�2|@��v.����!�g�M�]�N��s�=�~Tf���TT&�	�/�[�k3�W�P!�cy�	C�ut4��� �%��P���1��:O��xGAг03\�wH���� ��)N��;��Zk$=J<�ԋ�q�Ɯ��u�^Qzv�in��n6��=�62��{��Aw;�����`Q� _ذQ��렸�< ��R��"�p�Hio����e�﹧'��%NF�l`�Z����X�(��̀�6a$�/�4�C�ש*AM����d巌~�w#z���&:n�>iU���{U�.�j'�����^cbt�=,1`J���F5ZN��D"e�*�&�����!�&�3��$"�mP#R��
Ԙ����y_J@Ƕ���=���x��ESC�F�U���W��L7G�\2!)���������b޾4ٯP/�wc���Q҆ �S�A�Z��p}C����V���wu��h+ּ�n�0xH��is-��l�(����q�,�z���O0�v:9�Cؓ�e�;����(+"�9��1���~�uｘ!@�\���O��V��@tƤ��\�Z0O�=��445�O�IJD#㎮����U��(�|j9	a�	��m[�Y-jc2v��2L�����'����,&@ 9�����]p�v�.�eS�p�9��)���r��wȦm-9�^���� �Bz}��!R��s5X�ȸ���[�~뭠4���G�;��r�Xe�gt.�6}$��:�� ;;Hy��愠���O�m��D׺G�o�"5�`$6��Wǌ%�\p�vԑ2d��o�����%�J��R�K�e�q�7oS�i�-�Ǐ������?2pp?�L�<�ԫ\g���I�:5��0�۶�J<Ѯƿ���FY�x�L�{����r�����M���Y�b��RI4�j�TF����vu*�!�V����9�����qC�G������X�vC�:$��|����=�-+˫�g�����M��a��ME�+�J�%��
Xb��Dc�-Ŏ=��2�m�a(S�~{?�^��?k��ܹL4�'���~s3̝{��������������~AP01x@��Y��ejz����������ٲ���:��n�CA~��Sİ�ZvjV���Ž]ҮA��'�Uo�ZV�R��ݹy��޽W���A���g�
|ZfA�=U�)��}h���eH{@�COE�i��7w�e�ېϚY�}����~��}��ȼc�g;ʣ�\��K/�J]���{��	Z�&��}�����[���^��J �v��~�s�~��0K�+����kx����x�`t��a�2C�އ�i��e�s�����,T�s�9[ct,�{'��<���k���d�E�,���G����jtP.ë�/NF3��?f�@��j�!eu�F�kh��b�+�i�ϯJz�IC��ea�x�0��P"E��P0�e8.�f�pR��x�Р-�쑂���J]z;�$��k�vH�PLR]!�;�̱.E���}T*��ahk�Y�L�ky����Yf��pd].�fN��1�%���|��H��_�ś� %�rs�����Z�r�Cۤ��O3��T��zY�>�C4�D&���Y�?�أj�o�����.�R��h1����	�bdϚ��r��l�@��ǚ:�<9�As����;v��1����7?��*5���c�cr�-����~�;�J��5>��~���?)cSCҳd�f��R�(0�Y�ci���ƺ����Ay��W�k^�z����L.{��d�д���4� u�����ΏC��޾��/K6�RY�t�|�3?�7]�&�W����O��ߧAD]�	�5 j2�D���33S̾��>y���V������y���XըkG$ݵ�Ak�Tc���>�S�+r�i���XhU�L�'&P�Z���u�r�J����2Z�:9{�)���a������>�E)� ��3�����._��w��e��6���+k����0�{+ɫ/�BυC����t7����JMpO{\�KCo��s�//��B9���ˢ�(�o}��o��|Q�_H"Ѡ̎����|�6�N\+('�;^^���ȱk�����
��>��O��'�HUncL����^q 4G�G%��oɱk�u��D�?�,��:�#2:V�k��7��V�A!Bx)E��{����%{���+$�z����s�=Ζ��;�T�{xD>�����Ij��ճB�3�8>����3�%�4���c�'H�7�@���0Dof�b+���
�!0�zqbl����e�.���s��5�p}��|!�����!H��o���;�h�39����|�<���� 7����|��M�}�u������^Xz_����>caв0�^(���g�d�-�JC0� z��p����_�\Q�#Y�c�Fa�PQ�* �F
�H����v�9{�H������y`S�$<
Kd���d֌�A$�BT�VM��ll%8f���<0+Nǎu��1;��-�mJ������1d&�3k�:�>^�ňa�^	o�`$K��l�M�^s�Lg��̰���2�NUul@@��,�EpdS5Kÿ�.Hp6(s��H/A�@��=c� d �/|�Er֙g�?��2�C��.��~~��y�]�QV%�N	
�<t��h��L3H��_��W��>�Yy�{��5�#�t�<��	�XGZ�bUL��c�wM۬
�}��ByR��f�$W\�f��jY����2S������爂��2g�ޫ_�Jyr����w�Sx�!����Ȼ�{�|���˻��!J�Y�:���2�byNz��7\&?��]?��p��Ne��u�Uo�}��Ρ/��,:P�vڹ�ʥ��X���o�	C�s�/{���۞P�n���Ԁ�F`�Q��f���{I�������3����L�N�=��#��l���Tgؤ�@��=�h=�$��=�k���	�
�������9��L�1lK���]/����ꨛ��/� =x�|冯�I�#m1ubU���f�`|K�ҙB�o|���]���[~'�_{����_x1�	���sE=���Y���#Q���3��y'�U��B�>�d�e�O~�s��x�����%z�)-��Р4���i��]s����?��
##Cr�'�5�|��Z�،|�;_�����X.���Р �L>�`���k3��xԴ�|�_�;�zd4P}Z>���˛�~���~	��zFqu�uj�t$���Z�`��LH��e��/|R����z�c�w�E�{����TƆ�8��x�
�.�LH�UG��#�`�UXu+gK��N�1mN<F� 6\36�x|M��:d�Yj4ս�W.���'��w��s2� ���u�%e#?jؕ���� ��g�,W�q���B���/ۣF�k��6������=�Ѻ�g����-��oe�[���}/+3u���&��sT��e;*@y& �H5(p�6�n�F�߇�H8�4�����#��o�_�G����P�Z߶�.$�F�c���:���!u��0����F=�zON����
R�U��&��į�¯8���q����dY���ׅ A �FY���XF�����w�Ú��M����!/RFY�@R"�1��6Y�<��$Si��O�W(0��}���K�{8��C��GӖh*��,�k�BPp|>O:�6Ԯ��w�S/�B�a�Ȃ��5�Q���vu��$7��U�n�:3�U�Z�u�l�*���cc8�E C!�������n���my��K����G�N����$�:H�smm���l��͕p<$�xT����,���l��3N���ۡ��I�u�����[���&�6�i�����2M$eŪ��tYD�y�eϾ�jD��s.|��tu��I��P�Ҭ�T���}rpD5���_g�w��~.��앓6=O.~�k�:JШי���a��D��K^�b��7$_����7�7�q�|��_������oO�mA#k�k�(�P?z H�@H�O>!7���{�5�˯�T�xӥr��>+7��^���i��a^�^� �"���}�d��ٔ86.?O�9�l'�uc�-�XE��|�$A(��DY��}�a��������K�3+A��D����!u�Q�g�fY�b����D9�쳨�p�i�j:!�rA��	�Kx���B1�o3S\�2�+k�+���d]�ڪ5ꉰ�WV��D��!S?f�:�� �IO�th����s��[�([~PN޴�}j�� X��6�O�3� H"w���s�fYw�J�t�2Y�|���%/c����4��Y=�:L��0�X,V�M�3*`3�r�o���#�7n��.��=v���T�����8$�qIϾ��7櫱�'Y�Q��f�`������
!�M��-H����@���zn�{oy�{o�ˋ6NὟ�X;��9�P�²h�ay�L�����-'�J�kt^�h,��L=yw^��d�~��
%Pf��&ǅ��f�ft�^f�9W8^��A\36Bt�c��~d�#�j.��0gYj��y�wA��5�L���O'N�@��?�C	sdʌ�'�'X��� 4Q�1#�i oAF�$�����+�1�&7�@��c�1 ����&2+A�Y+]�l�\��a)�B�I����CA����fzԩ�l�J��d,��a�P����&�����h(��X0t5<U)/z�ºN�~ͩ�A�鵁��3��e
kj0A����g�]'&���G���&�Olod�7�Q�=O�"�]�c2�����'�KP��?��!��ՊQ���Lhm�6rD��r5��D���(K~(w�@����3�)T,C����1�l�]<�F�o{"�T]��a	ֵ	�`H�*D=��i��M?�����o0�N�YÚ�����`zM�N/h����d��M����5�:�ǟ��;�I{W?���u?��>�F��m�!Vr��r��Tc�{�l�t��Ǐ-��G�Ε��_���n�_޵U�z�j4��z��W��%1��◉&���R�r����#i������Vg@���S����a��_���7~C����y���˞#�I�w��^2�(����J��%K�J{O���n���æS�'q=<��K�!}v�NǞ䉽�tIa������e�_I��˖ˎ]ٳ�����v������?�Ϩg@*��tw�Psd@��_m���b�h;�*��)�y��Wݑ&Z",�j�{�w�}�r��_��W���N����e�<OS'�g߰2S�Vu���������<�W�w�_k@�H.y���#Ǭ�������R6o�&��)R肘�X��l��R��d��7!���
9m�:y�;�$�y�t-t�J"�=�L��W�!�Հ&I���!y��'e��������e�[�Δ��|���O��Ndp�"'��Q�mR���̄��g T���c��N�$�?��f��˲E�r�K.�+��Y�o˘���\�J���-��:�]�*t���F7��ζ��ʵ��,����;C.{�%���n���;��=�����yҳ��@�_�u����d6g롽�,�ғE��4 0�Pw��4��	]� ����tC�j��w��c��K�Z�i9��X�\��B�F��2�g��ZYZ+�m	��q$sq��R\B�����HY8��W�������6�P��*���[Yd�ɶ@
��!j#뫃�ĝ�9���XLiU�k����m�A6y��g��~�jb�W�w@5D�~�� g]�� #n!��([��g���=04��=}�R��(���f4=�k��F</��J�Q�Ԝ�P�\:���w��M�l>fي\ �01d?�����Ĳё�sf�r�ө�1��ב�g!uh� u��y=V
�5%qh�7kޣ�Lߘ�!�k�B ����}]D���4��	��ͩZ��Ox�.�%e)��A%��L��K߂ʊ�~���p�ʡ�S�g5�JCȯ�"G1�vL���SSb���C"��VD�s2ҙ���i� x-���}�k �� �m���p�r讽 ��k��c@ ��o_�A����-[)U��뺀��.�P �`�7�\��Z��^���5/�0��k^�*��O�A_@���������ȃ�wH$������V�l���8˹�m�O~��R!s��U+�7�z?p�X�B6'A `u=���8pH��K?U�A�+ң�nJ�1k������gd Ѯ`S�[����hWH*�<��S������k�3���:��b��ړ�/�Owj�Pa�Կ�b��p-�*��-[��y�|�_�b.�{�*���I�{Xn�կI������8P�p_$VRüb�J�����={�����<��6f�0�tK�]}��L�YAkP�^��Q�5��5I�k�LFz�3SSQ�<h�'��i�� �e�Zٷ�����H\mƙ�#���J��?\Gs�����><�~�GU���ȸ��IIh xx�3���Hn��6��|��W���y�,_}�|��?����2�Q�V�LƣiIh�Z�3[����7��?"����̳N�^�����%�zϻ���:�'4�J�Y�%��K6gD��]��9|x�|�[ߓ�����q�)�~�:9�s�s_��<�mP>�o_��xFi�>�3�x$��^�d���F9/������[o��k��+_�J��=W�k.�J�y����и�Gs^a7��g0Q����3�%�H���<�����[�cW��'�,W��r9����){�~���mVDqMV�c���#@a'�@R�6Az��g[��i>��+����@��f~�����?X���z.z@X������.!�z ���V���6j;;Rj<��֞�n5�292�Pd~�[8t��͟�[�g.��V���
�[1��.g��2��UIЭzx?�:2���UzG����]�|�mT��Ba.�at�M�.�h�K�Q���p�����G���V��B�ОV���(m�6�K�%����Y�|�P���z������/{힗��nv�����Lw�~����;��ۭ�W#��@0��V)��(B��e�N���1Nf�.���Hc)��~�M��]3U=����ဖ���KUF�Fi��yZ��XA�9���Sf2����fƾD���-P.�X��4�f�w���kQ�K
s��c���:���d)83�rh���R4��A�Ro��� �Uil1�8�\p��iF�J���~��2��)[Mob�s�M���d��R*r�tu�F�-���\F���fR%I�c��\� +��"���;���*���FCz=����˙ua��,���lP���]�HRy�LՉD�횅���PNt�����/
ֿ�|�oIR���'�~���ч�d�Nt�	r��-�{ծ0���x{ǀL�L�m��!���f�ǣF�S���|�c��w[%ܩ�-��j��l�]������Uk�I5�W��mrꆓ�=�!?�����m�ID?��>���9����L5tm�\�z��5=��	��~^^�ru^+��R�����������C˖�h|��:�8�w}�Bi։��|�7�o7o��-\g�MN04Ț%��Jp�>�v N�`�mO��cC ��^k{w;{ݹ�q����z�Y+����E���Lh �(�r��w���S��t�.�`9���� ���#eu4PL�͌KGO���vȜ:�ى��}�LIiv=��VjJ��i�1��LNO�#	�e�x����5 ��|�ߕ/�Fy�^&�_q�:�~^��lrF��J��e��6���A/��,.��7�l���s�Ҭ���_.�W��{�f*2�)H]�˒�%��۷KVϣ��J�ջ���9�y۝r�ͷȆMgȺSNeF��N�U�wB�ܩ���	sm���jc�D��Q��}�ɝ�'Vs�o���H6�'�.Ce� �)��Yk85�ٞm�`J۴>�W�?���T�Z���V�}�׿���������\8�`���)��o�^G�P�h�B�V^k9*����GOO�kfff����5r���a��'�����
 ^ߚB�����[�*12���q�e�Ey�z�a�lkArd�l���s�_�.�q�k��G[Zf�����׵������8f�=�7|�������SB�P�)s]���'4ˏ��Ԭ�$��h$����ؿhq�O��}����s���7�@��_<ԋN?>��_����|��w<�����]��kn֮F��(6�#���Is
�5�n�![�z*1�6�P��S5�/ȊeKdjlL�GG䜳6�ʵ��S��~9�K�IaV"~G����p�{��-8�	���5�A����R�Ԁ�����ב��$9�MP�"�<�y�ȹ瞫k;'O<��d��԰��E�De ��H�B������<�4���<Aщ�=;�U��Gnf�=�p�-��(�ց���e%��x?ѳ����O��folw�G��4f����LN� ȋ�lA�
�&�@Z�#�*j�5�������z	�q���)h�L0Y�J�(?���}���}��e@g�:������"C�0��i1iVj��ެ��Yq�L����5NOM��}��n���ưPa�\?�G na|=�n��5��%�mٺu++���z6��(����߃J���C�WCR���mFqQ~��[d�c���!H�VD��]R�3�ٞ�|��ɉZ���J���pǧ�9Eejr�6+��8�Ȱ��1�-Z*�bU�VW�� ����-I�����T��.kLhd�'���m�~ݫ[6�̀�Mp� ���v�;�:�I,�_.��f��4p	���*�ɨ��KU2��B^�B:Ej�|#+=KW��TF�NH2���= � 4�1ud�HX�mLϙ�\V�{:�L��F\a��m�r�t�/6�Q��ҩ�C^��S�O�:�F�B�X:"�D��{����η������?�F�����T���~�9�Hi���\�ṫ�����ڭ��*yL)Db�=<����CO ���㣲l�"�鍏��i���I*�Ԟ��������Ͳ��=Pw�h�!��ZB�?F�P��9E�%�)FU���}�Y{|�����o�}��ع����>��h R�J�_�v��`���_.��"b[#�Y}hO�ڭ�1�1~s�2�z�Өnx�q��,���W�>/>��e�f@@0�k$7Mn�c�N�&�R[p�V����큮Z_G���lW�1q@�G�c�h��y�z^��p�#���0�AGC��\3�7"�O�B}���in�cZD3(~����=�Nr횵��C�ý���^��w|��W_:�?y�o���	��~�����o���G����狕v��P���p����fU�g{���09�$�2�YGT��qǮ���	��K2�+�}��:Q5Bp�w�~�:��^sj�؁L��W,O�ð��12����A�W�D'#��Lu��=к���j���򖷼�@�A5씡�IY�j������N ��wi���G%��c�k� ԉ ��aHhd�~;h��Lu�5XFJ��'��3ڞ� �5@m��u ��ef	T��� G�o��������G�� �o����-� Z�p����Y�t�^�/��k��'��Ma�r�.�x�Y+Z(N�$��6�t��w�Yl�8��~�٧�����;�l�hR�B�f�"�]M3�D4('�=I�8u#��s��2�T[���>,w?�����$���:���U�5���3r���{-鿫aT'cH�r,�-Z.���/�Su���*%i�<�T��wȚ5'H,`�c��!���j�����L�3��96�V�Ҟ4��Q5�ͪ_��p���B�%�ީ�N,�v��Kr�@�4��)����6��ȺC��K��!T�4X���\Vci�~A�v<K�2��D	P���1��.ӳ��n}o̊C�`btJN<~��u��
zjGl)d3�[�r�>�}��ݩ�.}_�R��=թ�<
+�/���,G��ռ�i �}<33$I�j�6ɔ�	��1��MJA<��A�����[Ȍ���������qR �t�23b����h������)f������0�סvU�R/e�#�J�.3���u�L���&��ߧg<;1&�T�D�qR��Cz���ptO��}�j��\ӽ�T�_l�L�S��
�wN�S��B�c���3e.[\.�U����J���
w�xZ,��v��S��w�����e�8���s��	��W�h���j������x}!��h� �' H������\�
F왃&�Q�� *�+������v=�a�M;�r`���@��#Jۭl�ԥ�S��\�1��=%81���Q#u�w����QD��'h��o�ڀP���1^-��x%k�mF¦&��g���R��4� ����H5X��V��GЌ ����Ittw����L,|�}�]�?v��ƍK�޻}Ǿ�n�H��hG{[���Y�EK �"�x;�r��������l�K5��+W�3����fx�r�ϓS7n�=;w���c�x�4�5f�L�q��)���N4m�R}j�-�O�t4E�nx3��v�
�9������7���ttvʹ/�@6�z�|��ҀhX6�v��.5 ~���}hPӬ<`�,h@xh)D4���7�=�QU�OY^��=j3�l�K�"�Gv(bH&�YnoMz8h�W�U���y5��� '�����+9�8�s�R`�H��dD���o�5~�:H�;�72*�,Fu��i�~�/�����k�,�CIS�z�(���Q��o?$mm>R�"ϩ�@���G�v���Ȉ~��iW����:�h�����Mj��m���\I�3�֬grZ�4��$N�'��n��5�Kk S:;7������7.7h� ��x~�/?0 �k�#oJ�r�7~!���m�RxDs]7K6�t�\�޿RG��A&�fG�aU3I0����?��ȁ}��9j�0)pʶ��Wɫ^y�P�����x�vfs"�n~H��߿Js97+��mb�~�(f��rl#��z�ઋ�:i���,�n�W�JW����sp�f��ට�d��a����[�u�IY��k6����#���g4 ��Q���XW�����=�����ጓ�A�	�<�s����6ѣ$�l���ޮ�;������ȹ�%O<��,_�/'�p��ݪt�w�	;���H3�q��;��sRӽ�H�ٺ������W��Ç��K�~	��$��w��q�=26>e�.A�(���l����sx&��2���Jcf.'����>9�������*���P;���)����t�
���+t���p��/Y��M��iӵ��#�?%?��{)H�j����9x�G�>�H�B�UL� �j�Y��L9t�q�����������zN�_u���s�UC�,���j��W3Yy�d�M�B��j�]�UC���-O�d
���F,���?Iu�ݔ���VL�vϝai�g��EtLÛ��PX�I8�d:E�����F�A��1f՚C�#��p�(�pf|Ao{LZ��<�p5���P:$ 	U����z�u�ޯc@���s��Y���8��2����X��K)�@D�����k@~l�n�II&�@�5�����\t�_������|�y'g�|�M�~�?}�:ցH$v\�<x��՚P5�����YL`���twvHv�*+�-��N���/��|	.�����{el�0g��D�Z�\7����l8d����%�r7,��^[ khF���V*s24��U���=ݙ�w��]239�k�8��'�������5� z ������ه�Gﻢ��^�%S�i�N:���+��C��x� "�x���Q�cuK�3*AȌ[���6�G�9"����i])��[)c�����c�>�=���׭YT6������o�WfY����6	8&Geﮧ��c�r�AiP�ux����-ۦ�iE�5�NQ����eyu���<%�''l$4���=���A��ֿh	����9�Am-�NLiM��2z횁����He�� :5f4ܝf�:�9�d�d�^b�g\�'��IqvJ
SU���ɩ�g��XA+�mF	J���k�ǯ೛��\�������p��: Q�e��%t��j���]�e1�{	d+z~5 �=�X�e&>�8i _�T�<8��!�)�4��slODY��Sܹ�1ڿ_b᤾wNv?������yJv��E��Z\3ђ�8G+$��*�Kp����$�̂w���Q�}��M��R�ը���E����]��#��kvD6o�/;v< 1P��=�J�YR�sTF����
eV��������I�B2W�˗���	 K�"��-�k��`_�jS��ǥ���z���9i]b%o��&y�: �����Xi�֔��/#��Q[���eU����k����\}΁PK&K�HC;15-�W,�v�fL	����޻��J�36M�+d0T��9�Qx��S��N�A0��ɶ%�s�v��3`����^��+/X?�����¡Wl;���-�0�n�&4���q|��D�\5��:O�\�4m۪�W��t��5��\n����/���]����̽fph򲮞EI<��V9�F��ȴS&G��"��8�	�����nLd���V�Z�
�0��B� ��F�P��{Y ��Ȫ��' Ã�V t�!㇙T��}`�W���<K�5�����1�����e�����~V�"�'�x��Y�j�� �[�w�o`\߳Z�2pX�j�^�IT�ڼ�
T�u�f3��U+���w��W>�G?�_y��oy�O�<�팙�ɞX�����B�#gpxx(��b����0��,8�����[�~�>([�W3���K3
<���q�����F����}�Op^�^����Q�\`EL&0�v:�>@`��޳g�L��pA�F�b�$W��r�=j(מ�����%���,�����8�Z!;'��0��tϠ��j;Z>0���q����QDbt�h݈��{��Q�z|�0���[' `���<)N�H�R�i�@!�+��`h��l)�2*@m]D�>�3宻7���H��g�^=[���ɇ?�y��ߥ��I*_y:��>f�q�;�-n��R�%���9aI�u�/~�9��iyۛ���9 ����������E��Ï�/n��c��|0�&�����?~\^�ȚK�:@A�=�͏1�A5�۶?�Ye���~� 5�;�=$7~���ҋ/�!���PĈ���x4�@tFm���e���9͐��c+�1������'�����{﹋������A���?��ϥ�QT�0�,�#hp�G�e�&H�s�R��z�C�%݆`@m�ڑ��t/7e�޳�Z���:���6=G��<��ݞ����!(hV��^�/�w"i65��`	x��ܔ ���ig�����4��d�3���R�@��a��w�i� n�����?�Zm]���f�P�t�$;W�tT��@�k@�ogV��8"���X�"��e�8*��u�Q1������ʌ���i�^����{d����9��/�g�_n��f
1��g�aO'��܌��.9��>�U���>#���<��b�U��L���M�Г#Piz�E����eqt�ҩ6��=U(�H#<
�5}�|%�cQW������3����CWc��v�m����4���^�c[�f�ϻ`�ٴ�����O=����Z.~ı�C��矟=�E/�ӭt�G?��=�F�陊��"25>"v�>���rhh����-3��M�Q p�O������s����`�
��'��i4�#QC��erE= � �7����M�ddrz�\�@���`�_��W�r=�F�Ոv�� F�s�1Df���jF�������h�Zf���;n��3�5�>9.%������� �+}����T(Đ�g�p80}�yg�j���S����d��-��-�X9�-D|~C��������z��*l3DX>eS�է"+"@AÁ����>���wo�g��"(�5��4�@S=͔�1�~������_z4�������$,�)D ю�Cc�g�yu�j,���ܷe+���ӧ��U�>�f犎D�!V!�ecd��w�<�����0�@ R+f��ҽ��>DP�K�����{�U����C���G�n-.�R�8��:c1���OV�Z˟?|��4�^��:ŧ�,ZL�$@�U���쾎�}�9�V�">x�f�z]�HZ�	"�)�m��Ի4{��/|�s��]J�<p�p}�l<����;�0�����,$2�P�0ރ���η���7d������p�&3�G�j�3TS�p��~-w� U���FxT�L~V=�4�w�sN��rwW�:���{@>��/ K�	�Em�1U�|�8�~��06���ej�/��W4�s]�D�<����&Q<!�j_�+�I����q~�4��"@�49���4�Rm/GMsN1ɡ���,��M�OnF�>�����D�Hŉ��uG��v��ٲ��Mi������>�+���{�M����]�xG�-Cfd�@��1��A�=א�M ��˨C��{g����Ms��;>5Ɋ"�`��[�L�%$7��v�aa*���\�
9/ٲ�V��7��"�c���k	����J��O��!(mԁkH�yZ�5�w8��w����U��'"����F! �`HQ]�Y�+��\����hj@Pid���S���Cff�����3	M�YY���o�A�9���N%6�m���L��-�D�����������w��9�r���A	�;������ޭ�Gr�^��ԧ����O4F&2�oxN�ƌ>���N���S7+�fb��/�Z3�׌����p�O��'����r���s#�5�D��[-ӳ�<���(���D����x�܀y=,Ȝ �I��P�*�}l�R�x�i�p�Z5�yRY���fr���i�[�%"9�nho�[��C �-��%R$�l��Y~V��pJ��"�~Mn��f�Zń�n�B�,�h�����'oX��������VN.Z<045�Ӡ��-21a}���3,l�JѲ�åc׃�U?�8�lْ��L�Nr�#���;:�\��֡��b2�G��g�+�#�f��TI�9�.^���W�^�:ͪ���8˄�
zjc�*�� @/+���7\�����U������CY#�F��V��&���s^U�8�����^��J^�!0+�qk6h�2#d�#�%$$�� ���>�ѡ}�pN�d[:IU�٩:Ƕ�~���[�� y%�G�`S���1c�&h"���3�D�Z3E�G�5�dh�R�������q�Ų�q�݂^{2Р H�]��@@B��l����t����iF�-����Z�������{�^r�bf0��`�2*#�77��5�#*�d��U�U"+Ya�jXS����5K<,���v֔�]#��W-[L;r���' WНׅ��8�, �C���2�5��o�>u��� "@ݿQ�� g�Qf��2�έQՀI�`��'���F6[aI�!@�T��z��\�Hv?�Cz�5H���3�Q�SF�鷼�[��f��)��P�jp`F�0p#b+� �D9z������K���-�����5�9��:�G��525v���lU4{_�|1�~�9�03�<��cW0������y@�2�QO}�(l��� ��R�3v�[�RE�%ݓc#��j�2�l�F�`XP�E�(��MCM�h�c©\��d��Z � ���-<ô~&���S"d&�L��.��t��>GRЗ�Ź�]�J�^?�����=�H8���_�j�����7K3���������4�?��ωC�C����C�p4Y%�-��͙Ќ�*���k"�p$Ѷ?�$�}Ao{t��s�(Jo�6�Z�{3�%KԀ�����235�Q� �=p�>͎M��Dx��Ű���F�gmׄ:��J������ɍ������4f��xf�a٧�@,
��J��:���ذ������ݲs�^�	w�������+�C�TչP#]��(I3t�zm�D*:����+�'|��|y��o���ᑇ^�j
�?y��w8n���f[t��R��Խ}��t$V���h���"���m�S6�|��o[���O�hd^�� �X�l0��8oI��R	J3�D\ʠ�uM��Enu�5(�#3i���[ڻ����X�T�r%u�]2�ې�&=}�hT�պ��G`�`,����a�Wᰇ���U��0}Aq����|N��fh��1�W���8 8xd�LP�����C�L{��3�,�y`�
��2d�~d��Q#�fz��>s�/ƁA������5sI�C=��YuE<�(��j�qMM2��T�n��zo��Z��53L��N���l�3F �
dr�hf2n"X�eW�EL���&��.���b!�A�NTw��5�hNY>�k��2�<�|�,�Oؠ�{��I��z�E��g�V��?�#Ȁf�-�B����p���i���#Q'g��g\�u\/���N�jf�S ��!���?�lnI�%[!ص*K�]��%vm��:~ 12آ:nq3�͍J ��l���m���q���)�ϢB��N��|� :�� �\͙*��L��P�X�њ5+d��ܛ;{��(���Ӡ�Z�%}��Y)��S�8a�瀟���i�-����ol�5�M�	�����3���5x��P�y�q�u/OIo{T�bR�kG���z�
�G��Q[�����	��3�̳#�G���)PݡZS�= �/���ݖ�qHl��G�aIj���w�}��׬ߑD[Lf����aY�jEC�����ж��,��e�}���\r���R���C�c_�������V�a��"VeD��c���趿Iz.d���Mo7�,C��$f�+���v��}X���/_��Y#fAqZ*�x�ºP��j��e�YpM����� t�a# O���epdJ>��$oz��ҥYÖ{�aFE2�E~�df��^)���=��F���-[��=*�ӳ���%�D��:��Uu�Q�*� ��?��a9��k�B�?:�:����=��bŝ|1�Ӯwx<jӀMc�M��4Kܹ�i9��Mt��EX�-� L;'�.��|&D  "|2���NL��p4� ����-���a\�b˽(��w�;X��e����p>%yV|6��k�ʕ2N�%��R��f�ad�(�7 ����ei1`{U��� ����m!��Iww�������p�83�^ՠ���$hYձf=�	\_�_���kWk�=�ٸe�Y4��gg�� p�{v?���

�o��V�
��gw�h#��O��~v��$���-��<36Z�rŰ'R�R�{:��z���m���76�ۄg$���*��$��\2Y=SadVP���ءH�@V3m�h�ķ�pĸ�|\O�'��|6�Vf?�J%��2����f���Uk�Œ��q��'G8��rԺh1�N�'���8�`p�G�%��s�~�#E�����>���4�jr���d�J��FG�$��XNY�ˢ�@�~5| �M�q3�h�:�;U�Q�j�8P�@`��c��z=$Du�f1֩�+˖V���FI�]2�B`�nB��f�~h�g&�l7�"���>�S ��C�F��E0]���h�?z(m#q�&�Ys��*xNj�ʅ��kT�Ùf����@���v�;�|�	��чGN~�\��4�^ `�8�K�(�j���
������L����|�2o�*�sj;��rĳ�g�:k��d�$0��d[�ڼ��fF3z�O����e/��w���3�[�g�Ёx�����{�p�����!3
d���N��l�� M��l��m_�4�� �Hw�GZ3�s#j�}�(�90�6!ܻc8]��1��lSJu��){�t��r#�O���q�r�ò��{�(�"�������=� h`Q,���E����286+�v��{eي�z�U�L>��
=�Y^��T�H�REY�r��ϊD,����pE���(CE��"J����E�@� �[k����4Ȼ�쑍''6�"�<x�|`2���{���Z���E<C�8O���=_����՛5�8��mr�O:�961��:ʉ�����,�\���S6n�g��5Ǭ�� ��|�2��P�i�"�IХ��6ԝ��!� k[��*����+ 2���L�(i�w�jvaP���k1$/��C���[Kn��8�
Ȅ���ۦ�������K��Pe{�T20_\�+�GA<�<ᕒ:ހ���edpAz`/����pݒ����mUCZ:�!�Ly``@��R�e��ic�g�%5K�����me�SC����.���Ү�S��*�m�`@�jޔ@m�M�S	��MtU�T�k��@P�A�B �c�c �M�p�z���{�e�Գ��#�<��8J��Q���sM0��n�������O��;"����ظ��[B�,�� U�u�/��O����>V?�ѿ'����@*��$��=�_��<�HP�� ��jU0c -�P��cFF����3M�j�2�?[̐�ε�V���M�Yrk�á�NaRE�D�Tg|��F6%���Q��#� ɯ�qߕ9)dƨw��7*V�8��r�s����s�(�{�D��ޣz�p�z����|پ}�<��A� ���3plpʦ&�R�^��w<ժieU-�QQw7{�>��i�T�BS=�=�sss���Z>7��w�p=�B^b��#͊���b>�oT���؇?p�����9s���:rY��+�('� �.S�s�&�mv�̆�jٲ��:������T���iJ�\�+��@F���P�0>�@a�n���4�FI
�Τ7�fѝgx���v}�ޅ����xr7��,_��i�7nxlu�0����Ⱦ#�}�nu�����	�<	�*Ah@�Tא(�=�d�i@J��ڶkܣ���/��z�Ơ7<E7���9���zY,��+�n�6��q`�����u���Er���h���3kf�8`-yЖ�j�lG��Q��ǚ�h_�U�<�?LG<�䓬`䧣�KV�Y)/|�E�R���
��
`�����[&���d~���Q�"�m�Y������>�Egg� B���UA�!�12��()��f�/�#�Tu�$3�b~Όm�W��X$x���w��] �A�d��C\��HF35��6�P�rs{C߷Q ����1.�R��߇"9 l��I��98IЭ�r�R;� <�����G��X��V���Y<�GC������333�iqbZ�����:��m�������iNOMG�h�I����Wj'ׄ�_բ��3zz�dx�tu��x8(�#�����}f+���V�=[^s���d ��Bx�Q�=|������Y�T��^�j9��U�˗�8�{�&�,Oת��/�k�5H�Y���zY������.�!��gC����0�c��*����7
A�A=;hS�t:t�I�O&:uπ��	��(}wv�o�"�v ��`������`��f�!�Y�����沙y�E���W�kp�5i0�������-E�a�������UǌjŶ���sf�2uj9�����ho�����l[�{��j}P�V�>;o306�$a�G[��$��H�4)LI� =��^p��p�����r�U�ں��9�6"����SK�8k��ϐ�@���̈́�7�Z�a�<��F�Py(2�Q i��0�]ҍ
[��㩰n��LLN�r̶�`�A�L��òH�A�Sgi�Ԑ�(� adb�����&�f)�5���G�\@���iZejz��dR3_�:�I:+��]ʒ�l�����r��=�S>�����5�z�0��]� �,G�9SJ���/�#O5���>?zu���w��Y�T֬\F���]����$��0\���V&�^�M[� R;�)�7��ke[��)�F�c�z-�N8�`�2�c֬�%���sNZ
�,�Ho_��zU#�h�b90:3���L�F�*u#�rf��¶1�t�>�w�����ׂ�s�S��C	��V�c*R��8�lY�����q �� ֭��
�P�؇p���dB���� ��������@���,�`�ld,�k�W���-���*�4��!/�u�uO�>Cv�c�?*(y9U���h���F��" (�&S⟙5׈��1AsP���K�����$�g�*�~���cC�� ")�`�X�Vu���a�C�>�\'��6Y5q�T���j��M�����0���������A���D	Lz^ Fd����/'��G�i�� �M܏:{�ޗr��sD��L���g�Y�3��1X�_�Zn�<�� ��H:���cT��Q��πO1�Ӧk��U@`�R8�u*B��pzlF:�| �A(��;��2tx�k4����-�S�Rտ�Y�(�J��o�v��}-��4P,�1}�Oݻ�R��pȨ�e.�JJ�%�vJ�[�m3��V�Z-��w>��3�ʓ��V}�| �Ǽx��~�SѶþ��jfx���=]����&G���6{.+j�֢����_���_|�s����r�%��a���1�kt�^%��A�\UL	���>7�PP~ئ?mf$9�A��2��?�,�Y�n�ٹ��^m	�}���"��2c���d�2��z#�e�~θf
��@)W`�����	��v�F����B�
���X��j���=�gȦN1�
ʌ�S&�Aӓ(m�T�1��j�����?�3��<�6>1�F\�a�畽M����I��9�L�B��=*���A���q�}[e�ꕲ���8i��\ۛo�� z��;����lt��62�JX~��*N���F��A���j_-�?\oWW���՗���w�~f�����Փ���uvuI��
�!C�C-�:�0��(��U� ��z�➄�6 >0���k�
R`/�v�|1�*�M�����j��8
d||��#dD��p�k���EeLv�i�,�Y�&D:X`D@#l�M;(o<C���r��	�J�b����|K���3JS��f�$��AO�XY�(�/����O�<.�ep+dڪН$���3�S7�{�E�]� ;����3g�gkη�id���˲M�={�+PvE��{\�K��H�r�	F�NӫL� ��0z����N�c�'����f`F�I�z�uP޳k�\}�r����vC�JM� �3�X1�U˖�7hODҟ���h�7jM26�y�>��B�����2�F�0���`�O���8�g�@o
���W�T̕�v��?⡑ab`rz%;@R"���"h�W*��灙q�'���|��B��M 3P�qM�S/�&��蔯[�^�ٻW�S�?����p܎��&���O`SM���z<����9<k�;����w�d�����a3��K�ϒ�Ez�r�Sz%W!P�]����#\�c�ퟕC�3�HLG�U=�aI��>�,D�O�"v,��!ؿ?�Ǿ�L�T =˞��"d�ao3�{��L�X7nؔ��� �L�kG��FfThèG� ��piI,�5�M������q`��0@��Kv�xJ��(S"��J�����&	�CoԵ̨F��1n�p(n�k����ڲirr�q���g�oס������v*:�-���cpG�d�A�>��,��
���;)Q��F��HB�'f�[7�@6m�(����r=�}4 E��%Rj�%�t��$S!����!�+�k尲Q�}0:6�4 Z3M�f�c����SO>���&��g�%h��tjP6=9#%͆#�)�'&u�Pb������P.H'��Ѭ�-!�7/��J�e
?���t�f`� �Lk�Gl� O���[$��� q�L��I<�4�����3����O�u@P��|@c�cr�guf�&��'p�9���#�^�ا��W|���h�pL� �4�|�`K�˒Lǌ���CF�U�{�p���NQOC�p2�O�7�K��c��1�x�,3����~��=5侮�x�-�4UQ����6���i� ;��h�m`Yp�1��V2��`l�{���:��0�Ha:m��빍�wH"q����O����&���Y7�Xh{�/)�;��0�'DR�y���p�9�����V[���E�	Ѵ_]v�_]/�Ϡ{���JeĴ��`��>�� 57�QP��[g`� A9�&y��/de�<��8F��j��r�/"�6J@�4 �@jр�U�,p#?����R�g�����Y�T������Ԍ&)�GKv%d�0%ղ���zF�͞����v�:���ú����v Vh��$W�+���3�3	���q=�#ȗ$�N=�vkj2���&���ko��:^��.��<t����J�X%]<a��,���Vm��O	x�2��V?Հ[}�g9/�pKԔ�4���0��t�ht2��r�"�C6f�%~dZ���1�k���-Q�@�23>1�,�=�4���l�t��^w�Z��u�p���n���2P!ZmSӳnݼy����?�Y<⺁�~�3kʵf�f��p�O"K�|�[=bl��D[�{F'�Yn	�=j�J=��e�3�YR��	f �Y(�t_�����?�l����p�s5�t���!���]�"U��q)8��<y�g3���T��^}����F���7��E`���E�F��V#95;!�]��Y�ȷ�@��J�0�C/H �Ys056A�MiQo�,@�� ��Y���;���X|���(��^�bk���dG��^deh5��`�[d5���{j�`��4�!1`O�*-��h8���u��/|3mbF3]� �������n��@�GJ�$�����%U+��Z
�G��uM�6��ڂ#��ǽq� �	��3Z�a*IM��ϴF`'v�������E���D�ۦ�B�!o�����4��<H	�:&(w�#�<�ѤFき�ƽ>�� �Dm*��"�a�zr��ip�*�)�7=��$�*b5�r�;�UpO"�
�:��@;K���6��o8uTxLo��}?޳����OEL�c�6�{��������1Y�h�<��J�jۀQ�1�g��#�7����hx��4���7�˞�hz{���i���<R>������]f�'�ĉ蘪��[<�U�Vi���@k������T⾠��@�������?C���9�82�@啄�l�+P'�\�5�EF�>��JgM�e&�-{�<�&+FϨ�r�	����P�>n_ ��^��ay��#�m3U��M�yalh��F�M������i	�v�+F��`���c4�{�ɴ�,kȃ�o
���D��b�ƲS�禟���]�&�w��k�%^O����m�R���Z��O����ie�VaY�ϵ�F9{�.˯���� �`���"e-S1�D���F)�����k��hc�ǄɁ��4�c�?[Sҕ�#A+DF�c������6H"�i ��ACԿl/����^�b$:c�ijd�b�:]V��G_����\�b�#P���fpM5_D��9�]��::Q��@��OO��<�U�˘ٻ�b1���k4�BA0�ՉՈFS��QfN]ρ~���������y~�����B��G�� �f ��"�ֆz	�0��%�j���f=����; ��)7d�2?��0x-6?S�=��������\���'ۢ^�w�';̊�w=��_x~-2���ۼ�2�{�h���8hF���8�{؉��wo9��W���`��4�ES��5
�&���d-oT��Z��}b�9��r�����y������
8o�0��F�+0_�ka7Z#-Nj�L���2.�L�@�M>����YJs��W��;����Q�=ͅj���f�D76&!�k�T+�`>k<>������s� �_�䌑���2�^`b�7�xd,�	-q]#څ�f����16J��gK9�V��+�Sh�R󜸧���b^]=�Ʒ��џ�C?E��{>?2�Q,J��ɠ��X�o";�B�s��5����w���N6�Hzs��|�����R���g\���7���;��Q�o���"?CXo62���1� g<����mo�ú j	�3z�b���::I�0=5McM�%�d���1�@+C�+*M4�=���y?�喇w��?vRoo��,n���o}�篝�ɞ$�D���IG2-��[!C��p���q[��`�7F��;��-gi��f%0�A��`$o� ��`���2�L��}�G��G��Y:/�G&��;��y����`%S���l&7,��q�1����N}��Ġȁq��?�jn\wa���Yb��
�7 �4�y  �a�0����P��aR��`�1�-۪�3T�,z�3#����I�
�A��=dZqސC�L}j���f��N��t�|鈽^y�7hX���Ϋ��8�"�_s�Qۦ��5��fm3��2�x��{bμ��;�֫�P�~ƿOͱu}����2��ubWZcKGz�G��/�F �i"�~Akm�#BC���=�z��	
Iy��R�C����m��چ�i.��7�@A�l�q��	dI�������� � B�˫�w��eq�G,�'i�Yj�䴪%f$�9_Yl=�VF��2��-�����u�d;p��n�;��簆ã�\O�t�Y73���wQ���AA+0�{�L��O��h�����y㐭g���jd���GkOL�3����//�����I��{�������t�{����e�)#�!	q "	�l� ȋ Yd�mVFVYd ��_p IȰ��%�4dZ����{���U����7��νU= �V�YS�U��>��;��w.��@+�Z�9�!��z��}��?yQ�s���F�4�D L�Gy�(t�\��I[�37�j}1W��^�a�5�B���Wt��z�m�����eg5�����|C$R��=]��u�q{ȱ��0���ذ@$�� ���/�fy����176Ӎ뢟�O-J����j�m��ͦn����5����G����_~y��g~W������~��|���k��V<�J���D�4)請���8f����Nc,�5����{b]�����PsF�Ň���>BȽS���;����S���k�Ũgf#(�*U,��#T�c'!�2=�~2�ڤ�$��P�V���*�?��Z��!�[��K/<mB�j�?���\}G6��^�:�7�AO�~F;B@����Gf �/�#��΂>��!l]l$��������el.����HJk |����h��'���~�����4׋я>��P�] �
7J9�]�j��w�n%~~!��V�x����m�Q~�иe����Wb9��D;����^xT6�=�?�%�N!ǋ�@�'��1����)ok)-�|x��:����W~��At�ҥ+�be��N{-y~���3��N(��ܢ�����ӽ��;�
��-����G�k�	�r)�~A��1C������Ç����6��h�;�s{�ɼX�I!�1�� �Sx��є�2S�GKcH��ȯ�ޠ$Б]�dݢ���� �b���[<�����9�an�0��@pc�1S�AA�e�
��hL%�����J�R��t���!���=E ��O!��k�� H�jzU�a������T�<�9�)M6VV�[���?y�a����2/�x� �z���;��F���4��͕6�lz::��,K��y��1gf4��CK�S�ױ���GP�f5�F	���|4��3Ft�M�<,ʳ���Ăa;���O��"8�K�.��O��N%S�1���_<�K�?"�F�,��7���V.�������?X���џ����������������>������o�u�?����Ooݹ����~!���pcSm�L0�(B��\�\(&"����.k�Q
��<��M�ya���ϯ���U�KA�	�,�"�f54�_Q�̨M�2"�:�b�Vd<���K� �6m���(�[���J�r8��0Έq�76��pm��F<u_���
��`DT]c"�e������V���`AIS-s�~ﹼ����o�3H7�� (36-��>ڰjHR)X��2ͭ��,ЃY�@�g��	s�@ǣT�$�Ȕ3�ʥ�T�Ƥ�q��![
\��S�%�2��%-jX�s}w�?�a���HG��i͝ks���S�a�<Ϟ��/"f)�!`S�9]��޸�R��Q�S��t^70&��}�	��r�	h{�-p
�+C�3�5.y��GT�0Z�/G�䤡�D�������ηJ�L�4G����}�ôr�0�Б,~�s�e�y��x�@�7X��H�
���Tʚf���R*E���5�-R\�ݼi^}�؇�Y,�M�cF,x�Xw)J�q�>���'���RONN�	���9A*�M�c��I�Rx�>��=m�(�i�pzm�������Y2���aSY�l$�fKs}��,�,w��٬3���L)t�������(f3�@N�2��e1[���1��n@3�u���������38�&c]��Yb��F�lEa���,Z��=��p�B甇�x�#� `���2GŎR��瞰iY:K��}2=��1�<�+�N޼T�̝]���-J�Ξ1�jl�������^9�N�?��ᵓ���߼�������֍���魭I�e͠,��~[�T��o޾����/���k�w^�y~�{;@�)+��2�q-��0Z
F��(��!Xc�H{ã%&�h�Bׂ�'��V��>�S�πT�^ ��/0�a�{ay�^uk��hO�C㽠�s=z���-����g.���l�`�u��G4��xU�s��X�a��$T˂��W���ޡ�X�pvTV �a�s0z���z����u�X�+�Q�W/_��@l�h�	���O��Rh�:�P��aO�"0P�A
OB�굑�{�6�{p�b�m��u��� �=2��`�(�{��������T�Cr|��
�L)������A5 ���05(���Gg�)���bp+cg��خ2c���'O��a����E����@�4��;��q���@v|tBs��u��~,�&6k������Q��؟�ۤ���~��) ��Q׌�w2����R`'��b)�:=S!�&���q?>�gv|p����~��:�|(��ۯ���W�w����|�p�@�ޥw��V�M�5c~JY�趇�$[.��@j%��_D�'"#"�~N��?z��T�o���_�q���H����?:Z�UH�,��Tr!#2M+Pf�� :F��LӢ�H����F�2����>�ː~+:�,�r1V8F"�P���s�51.0��H({�� ���X�Oc>��R�8z��2�0�T7�F�XY���b|W��\� �s];�GDrb���0F�Z��3�~�d;6���.hT�4M��.� OY~8���#�ki�0��n�N����,R�����D��o����:[)H)� ����#�� P�R���J�Ճ�ն6�7N操���l���w޻u��[w�VW�綨rq�'�v�d:�vpx��l6�6�UD	.lf�gX��R��̼��ǅ�1cP�Az!���Y������D�1K�����wt�V�Xk��㸑sz�H=(P� cWΨK����J��5pJا�JV?I\2��ަ�:jh�{"����DWMGl�H�,�m>��C�By�����|�W�+/?g��#S�?2�G���\cM-�?��!�@�g�������k75��F��0gyW�`�j�ԭMY�t����+��A�̎;`)���޽O���ի��3ϳ�(���ԵsfJ��[�,��T`�Lw���{$��`	�z�4
��b/�tԓ �P��]?:rŗTV��3k�e�r���7+�y%��m_o�s�
 �����G��H�qO�;7��[���_��ٰ����6���AX.h�����C	Dz�2�z9�<֮��K*̜�t6��X���׎El�鍖Ϊo��e57�������7�nU��Dp5�3�0���*�@�O]}�e��UP��h�`��@�ٝ�����%dؔ�o;��Y�?��jdH�
��D��uK��a��������y�o��v�k"���a���@Jf���	{v��9,�+Ox[gϛ���_׽*r��;w�o��Dh�Xy�� ���vP c��H#��k�x0f�Ps�J!�ZĐ0�#w�_��ԋ��� Ym.�ucuC�:D����n���!�Oy|���^zq���m�/ԇ�`��l�������G��
��Z^x�=�V<?�^gAa�L�)�<��(Hx,�;N*JO���c�f�M>�L���� �.~&�u��np�ˮ�����s�EE�����=@jM�@�{t��ؼ��{�;�3��evEo�L�ۀ��f=�v]�s}R|Ɇ��^�!+d�����u�/[��gu;i��J�=��<=n��x�s-1`QZ�u��K�q�@n�3�2�9��2��f�r.��/�WaH�K��5O���4���_�8��;-�,Q����f1��^����!��s�[@�B@ �E��m({U*"Xv̠74� =1��,durL��≐%k� �&j���ͽ��'"h6.�CY�"�̹�W�_�B5g���Vb	�����	qШdg�\Y[eר��y��3qUh5P��j�#���Kf�W^}V��C2x}����xy���g X;��Jc ��V��3��f+(��q�&�xe0��2ocD �e[O��}�Øc�tEOA�D��9��@e�j���#ݗX��R�xag�:�7%b�e�@�8�0Gc5���k�BG�t�P�d���J�%X"�5t;a�����h��"C�������i���nP�.�概Y�'��Ne����|�K����u*!T�t�|{��.[�UD
0H� %�W����_���Ǐ?6��C�GT�T".^�j�����&�(O���8�tD-pb��Ν_g�eH��W��	87BX�b=`��D�U40���ߥ�x�)�֢�Hg��*���M�p�cͧj! ����ɺ�:w�l�='sv��h�!kֱ�.����`�eo>z���w*���d�贩̙�-Yk��U1�/��d>������-RPon�3�8Kc1\/?u�T��<�~D*c�U �=�	y}1.IX$�� ��G=b�6y��_0o��[4� ��w��
Hݽb%�TE���)��g�7���o���Wo����>hm����D��.�!�b��	`fl� r�e�!'�ō�yf�Sð8�z�	)���3��5�r3��}��fi�ŰB�
�3$�>��Q�(��C�Í�	rgm|,k��EHc1I���v��2�{֧�_ϐn�!Z�
 Iu����zz��x�Q�痵���gOb�]�"�4$�l�9���њT�|:
�R��Q�R��F���%�z}��4�N����@.�e�JdRW�FhJ\]^��g$�V�L��1���|C���Z<���J/ê�����ks*�;>���jϔ~?:5��j����3ċ�:e����ɑYo�yr�ɃL�V^���ѫ��\og�H�،�L+&D���LP_l{2>E�3��#�:�+�|~�z�����d��� Gxfz�P����`a�=�����S
P����>=¡F^Ę1)}˒D#����^+�ˢ� \#GAD�ó�Y�9��l���/P���S.�N"2as&����# �H���p��sd|���)_�/�tZ�����(�]�Φ�h���J ��;NSvVyP0����ɨc����2��&��W�j0�*��/�O�:��_bm<�tG )�_�F�O��f�v�'�
B��#�&
z(78787��d��#��/���j��9t�D��\�:>8�*
^����@����g9ǵ3s����Y���8<s�g�]4�/\fEɵ�o�jֈA�F֭�1*���,M!�{(�����c����sb %`R�l�S�n�k��d́����e� �˯�b�,�m��g���T����)��������{�������Fv�ˢV�va�C5[JI��B����*X�����(�9Ȭ�U]xU`cg2��}B7��H�4�ZE=<�[j�b"c��S�����1���?�3��#�z���P��A���3܉�9�l_�C>��"R8�����T�@O�1� z��M�#GH��D�9��m�8�����b)�b�q`�?�:��=�6M�"�5"�`)R�����b�ī�z:���,U:x�hQ �Vh��B�}\�p���ජ���*Rp��_�pb
z\���pa6�����`�<��-]��#��"�SΉ�c ��p�a��h��_j� ^����x�)��ը�[�^� OD#�Y/�l^f�NU�Ε?g�d�}ԁ�� cG"�0�5�C�l�$��xU�,º˩D"+���v�����4�gh�9Mo�\������8S)CM�L��]�Β, ��q����А_x
a�+W�q�c	��+[��0�N�0 +գC�#W��.`�i9pC�@������w��="����E��o�������@�SN��O5�ʆ�%��c([�q���QE=	��H��,�����n�1i�˲l�]��S9n�C	-�@�g�r�yI@�L�qC�@AeS�'�����Mt<� K�y"�(<�3{���|&LΟ��\t,��a���#���|������,�խ�4 �k�fgw�e��(f4���|m��q��`����ڤ������)���}���Y��@\��Uo��<=M���{���|��������)t_��������ћo�����U�7d�lT~��Bl�5&^Hȕ���:���FVT-�r�*�Q#�m�;��S������m��܎�3lg�l� +������% E�A���V�3��@Q�z%�qrǢ�z2"B;�Ŝ\^���_�9y2��6�YR�[܄����� %�]��f��*9l�ޠ/��XZ�`��)ߐMl[�	�[$x��ޤ  	@IDAT�kĨ��;D-�.���F�6���w�^ФE����p&� ؘ�P;@�A!b��[/�wD탋����~5�����|�Em���s �z��hƹ�]���̻ 
\�rM�2.Wnu4���Z���S2�2�NlA����GͼGj9�Br��d�����)#"����$�:&]�&��z���d̻�7*��.l�(ā�n�+<���&��X��>��=3�j�o��"WL�"�	\�v[dD���
}��~a����}P9�s��(�`�������:��<hi��[�JbO�u1�b ��cyB��Z:|ޫa>�J���t0&��W�Nl�5�P�����ıo��^�ڼܫ`����[׶�&GhG,r(�A����������/2��(���^*A��"�[z�aQ��"�i���=�Q��	V�:������K.��zGOF���G/]?k��\oQ����(Ѣ]�GN�Yb���~��a��>4nauiDN�"v�m�� �U|��t���5�S�kȽ�t�j^��\�|b�O<>v(d�:eΪE7F�7ZI������ǻZe�{�q�l�A{t�9��+RG���i? ��=*ox�0*h̰��.��΁���qɀ����U3}��>z���?~���?������+�����g�����^x��Y=>WM&��|�Y�\��V�d" f]�9�E-���,Tsm����BCcWtxm��E��6�
Y4���'�8�����}-���%�����a��E&"ʉ����񆑀���):�u5"�-)�Tt7��d� ��
�{�)���l,%�[�*��Z.�+6N��],~�d׈�e��d�����k�/E?�z��܀�~���+㉛��`'�ߠ�E�3�ᚎH����@�����uy�&�Q���v��=�(P��)�Wx@�6�u
h�]�Z�u4h��v袁�?Kِ0�>��a��n�;`��
N;��d��<:��i�؄�,�Z;hڮ�[�9*'����s4=�������@e��ڰ4u3+&�G�,rQ$a6i��"o��=�M.B��ۼ��MS�\��!P�"w��$�cG�dM3�ɂ�I�^k� ��,"�"!��/+���]jP?��^�"�s1.���V��;y޲����3yz)M�,�K|���(�:�qA� �Qs��.�j���]�.�r�FYqp��e�<���7��!�u�O'�mi�K���k��M�@��o���>/]S�e'Ƹ���!vŚx�Ӣ�6?<�ӓI)K�'
|JtVM{uUm�����uSȸ���a���G�F��\�'`���u�� ��^�P��xu�(]�Zy^�{��@�7��}��͉�rB���� �Uv�5��iЈ9+6�@[���-���D�Dޅݶ05�%@�ṧ�P �BRa�4֑:��eU!ZD/$� %B�!Z�̶���v�<������=5xRt�]�8R��
�-JR#�ȑ g� ���h]���J�\�jRd��rB�R<^`���@�4$��+�R -$�l��H�@������?��Ё-���XW��`K&������nQ���_��o�濹m~N�gV���uk1����������]�.���K;��;�	��s�U��9S�����{"��}�؝��p�-��4P��K�����p.�	�~�]�r03�3Sd��4_2tG?'b���'ڜ{t�������1%�����e{�=�U/�e�>�x��fw�Y�����Q�r6ݳۃ��0��ɇ�Y���U78س���G߬W�������L�Y�=q����=~��ѡ�x�t���~{{`�?�����࠴x�������μp�WX?�!l�^�*�f�n�B�V�A��L�F�U'k��u�1�a�N����,7�w3g��ySTkE�r ���t�+�Z����d����I~47G���$�vu��V�<Ԧ*��>X*31�ꐣ�Y)�e6�d�'������7�h�3��e�O��GS�c�������'py�s���Y��1b�&+:Q�aj���ć�S��5ѸM�f��du	}�ս��mC{U���]9�ۺ�Qq�L^
<�x��s9�Z�t#�5����Cl����Q�Y�.��@��(be8ۿb�1�2�c��m'�nK�F#�滁B��a�E	
�{_�Q'#$> �O�z���Yy>��-� ��8H�5����p�H! M0>9�����Mf��r�=0n0xD�0�I.��\F������x<�r���K�ݹ[���JN'Pృ�U3F-�idjq���pKK>�G�w�_�_y�W���7�Z���� �Dʄ��    IEND�B`�PK   W�X4K��  �M     jsons/user_defined.json�[mo��+�>������|������	,;9�\�$B�+�6� ����%���5)�
l �����yf(~���.�����*,�!��O��7ay5o��pE�/W�u�ѫ�~[�8�_�g�v &?_\�UӬ�L�}�	gW�s���'��`~r�h���t��9k-�������!��E�(ƣ�4vڡ�}�Z^��`Õ[�/W#�����k��V�	d�ǈS0o��e��ZZ�cu���]�G��L�|�.��ί./��As��RZ���c��N���=Sqf�y���������0�ő���s0>l?�\�ہ�/Z�ؘ�HeԞ�2��`~��p_�%<��ꅭC��?����^�>�/9Nۏ���	����^ : (�����pl� �~��C ��,�� 1@T��fg�go��?�麟f�Η��ß��eX���l9���Ng��B�y����6Ԩ����c��|���z�,�b�a�p������������wgݗp?�?�]N��X���2 r��Y�6r��q�"2�J�U^����/`����!�j� ���4�\d��Z��3ZiI�I1��
VҐr�mpE��r�	��IŇ�~t��N4���a������L�d"�"�Q�@�N5�.CA�H���0te�K���%ҋ��􉗄�B�뺃���I�����E�c�1ϲ��['	2cHvk�4o���d�d�����C\fʼ���L&��W�� ��/�P��6� o	�'X���,q^ �P��|�!�ru9�� ��3貘�n)���xM�o�]�_�!��߆n�Pf���e1�j�2���
��&d� �_n��G�ئ��43���%fK�<�����no��@�ZН�;Н#Y�AD�z��Лɪ����l.'���b��}�,�`_�eV�ͼ�#�H�mA�a��Q�j�qr�tw�a�������P	�k��T1�h�Gm�k�0�����s���5��0c�����C���DW�S-R���J�K~A*%83{�ޛ�jX�8:����M��߀�>�����_
D�ƾT��Q��'?��g?Oޝ��??��%��;`�RI���]�{�vRe�G{7���W���O>\.C�}�� ���؄�e5�H��\�1�>�� 7�{c�E�&q�9��q�b�]t��2
r(�	�:�z{�^!;�b�d\�=���R�gzoCN��<���zo�|�/���;�/)�����		�����q銣6��7\��� d����V"x��}�������d�9[?�t`��xI�����E39��S����1\�D@�`�$#�:��>�^���LpE��Y��KD�odǠ�U�!X�Q/Q�-H���*�>�VDjg��{_�^��4h��zi��&F� _x����	���c���7�UI�rB�0~��R������sI~ā�/�Y�zz��=�r�q�FbYHG�N���D�p���|9�ogo�����q*�U�_�%��f@� t^"l*��P�*�]��{E�ݶ1��As��/)� ���{I�Ѕ���I�y	%}����I�yIY��~a��]R^l��4;�/i_RQ�!~��Z����S�L� B��x�!G%�L�!��Bv��Ih9�P�H�2I��/� ��6��$L�b�~�%ڙ�����9h�XB/�}4��e9��HdgU�Kz�J�R U��%F�R���Dۗb�K�D�Ae���/��A{"E�r�~.�D��;0� ��w�2޵˶���
��,'O��҆�$�rb8rVz��MD�	A��P:���;���E^G��SP�Fj��"�ߧ#>P���"e|׍W��R�����A�Փ�
�9�Pq��x�!>��ni��O���� ���j�'3�?V�Ͳ�'���D�B4q���H�背�6J�7{2c_y�+�}屯���W�����>�����8/~yfjk �0AI��(��#�P�zI���i_�!<��3�v�b��JӺMł&������E�� �J��i]q	���<=9>8/��>�P�%A:�랈���d5I�D�\V�~�dE��uW��HT����W<�t�W�����>���J6A6��2}��,�>�8��S`1��3� �i{��0j������xF6���gd��xF6���gd��xF�L����3��l<#���Ggd���B�x!|�>^/��������B�3����'C���PK
   W�X�Ή�0  Jt                  cirkitFile.jsonPK
   V��W�vh� `� /             �0  images/360150f7-d3d3-484d-baeb-b64063d02086.pngPK
   "��W��L�h� �� /             - images/40f7d2e4-4064-4959-8822-d1932a7058e9.pngPK
   "��W��L�h� �� /             � images/505d58e4-7e58-4ce3-be43-3c0c0a024e39.pngPK
   Ŧ�X�i�R�I �I /             p�	 images/5472dc22-a170-4182-a291-403007edeea8.pngPK
   ��6X\�
�@ 6 /             �, images/56cf4bf5-9c71-4f2a-9d5e-98f1de214099.pngPK
   ���W|�߮�  ��  /             ;G images/61b75eda-77d0-43e1-8746-2b678f56ccab.pngPK
   ��6X\�
�@ 6 /             6� images/846d17e9-ef90-4979-be28-74fde6feb977.pngPK
   ��W������ �� /             � images/8db8bc11-a89c-44df-83ef-15ccf3dbf879.pngPK
   繆X�=z� C� /             �� images/9595c21f-5942-45df-b2b2-1a139a6dc1aa.pngPK
   ���W|�߮�  ��  /             �A images/9c4d998a-0b1e-4d84-acc4-3fb4cfcfde1c.pngPK
   V��W�vh� `� /             {� images/d74878c5-97d0-42cc-abc5-9bd8c586a2df.pngPK
   ��W������ �� /             ��" images/dabb1173-90ac-46dc-83f0-6b94d38ee5f8.pngPK
   繆X.h�G� � /             �v' images/f072ed7c-bdca-4b42-938b-e27227333132.pngPK
   Ŧ�X_��.
 �	 /             . images/f557da7c-7f17-4077-a29c-07168c914697.pngPK
   W�X4K��  �M               �%3 jsons/user_defined.jsonPK      �  �.3   